magic
tech sky130A
magscale 1 2
timestamp 1685731389
<< obsli1 >>
rect 1104 2159 104144 105009
<< obsm1 >>
rect 14 1844 105050 105040
<< metal2 >>
rect 3882 106594 3938 107394
rect 7746 106594 7802 107394
rect 11610 106594 11666 107394
rect 15474 106594 15530 107394
rect 19338 106594 19394 107394
rect 23202 106594 23258 107394
rect 27066 106594 27122 107394
rect 30930 106594 30986 107394
rect 34794 106594 34850 107394
rect 38658 106594 38714 107394
rect 42522 106594 42578 107394
rect 46386 106594 46442 107394
rect 50250 106594 50306 107394
rect 54758 106594 54814 107394
rect 58622 106594 58678 107394
rect 62486 106594 62542 107394
rect 66350 106594 66406 107394
rect 70214 106594 70270 107394
rect 74078 106594 74134 107394
rect 77942 106594 77998 107394
rect 81806 106594 81862 107394
rect 85670 106594 85726 107394
rect 89534 106594 89590 107394
rect 93398 106594 93454 107394
rect 97262 106594 97318 107394
rect 101126 106594 101182 107394
rect 104990 106594 105046 107394
rect 18 0 74 800
rect 3882 0 3938 800
rect 7746 0 7802 800
rect 11610 0 11666 800
rect 15474 0 15530 800
rect 19338 0 19394 800
rect 23202 0 23258 800
rect 27066 0 27122 800
rect 30930 0 30986 800
rect 34794 0 34850 800
rect 38658 0 38714 800
rect 42522 0 42578 800
rect 46386 0 46442 800
rect 50250 0 50306 800
rect 54758 0 54814 800
rect 58622 0 58678 800
rect 62486 0 62542 800
rect 66350 0 66406 800
rect 70214 0 70270 800
rect 74078 0 74134 800
rect 77942 0 77998 800
rect 81806 0 81862 800
rect 85670 0 85726 800
rect 89534 0 89590 800
rect 93398 0 93454 800
rect 97262 0 97318 800
rect 101126 0 101182 800
<< obsm2 >>
rect 20 106538 3826 106865
rect 3994 106538 7690 106865
rect 7858 106538 11554 106865
rect 11722 106538 15418 106865
rect 15586 106538 19282 106865
rect 19450 106538 23146 106865
rect 23314 106538 27010 106865
rect 27178 106538 30874 106865
rect 31042 106538 34738 106865
rect 34906 106538 38602 106865
rect 38770 106538 42466 106865
rect 42634 106538 46330 106865
rect 46498 106538 50194 106865
rect 50362 106538 54702 106865
rect 54870 106538 58566 106865
rect 58734 106538 62430 106865
rect 62598 106538 66294 106865
rect 66462 106538 70158 106865
rect 70326 106538 74022 106865
rect 74190 106538 77886 106865
rect 78054 106538 81750 106865
rect 81918 106538 85614 106865
rect 85782 106538 89478 106865
rect 89646 106538 93342 106865
rect 93510 106538 97206 106865
rect 97374 106538 101070 106865
rect 101238 106538 104934 106865
rect 20 856 105044 106538
rect 130 31 3826 856
rect 3994 31 7690 856
rect 7858 31 11554 856
rect 11722 31 15418 856
rect 15586 31 19282 856
rect 19450 31 23146 856
rect 23314 31 27010 856
rect 27178 31 30874 856
rect 31042 31 34738 856
rect 34906 31 38602 856
rect 38770 31 42466 856
rect 42634 31 46330 856
rect 46498 31 50194 856
rect 50362 31 54702 856
rect 54870 31 58566 856
rect 58734 31 62430 856
rect 62598 31 66294 856
rect 66462 31 70158 856
rect 70326 31 74022 856
rect 74190 31 77886 856
rect 78054 31 81750 856
rect 81918 31 85614 856
rect 85782 31 89478 856
rect 89646 31 93342 856
rect 93510 31 97206 856
rect 97374 31 101070 856
rect 101238 31 105044 856
<< metal3 >>
rect 0 106768 800 106888
rect 0 102688 800 102808
rect 104450 102688 105250 102808
rect 0 98608 800 98728
rect 104450 98608 105250 98728
rect 0 94528 800 94648
rect 104450 94528 105250 94648
rect 0 90448 800 90568
rect 104450 90448 105250 90568
rect 0 86368 800 86488
rect 104450 86368 105250 86488
rect 0 82288 800 82408
rect 104450 82288 105250 82408
rect 0 78208 800 78328
rect 104450 78208 105250 78328
rect 0 74128 800 74248
rect 104450 74128 105250 74248
rect 0 70048 800 70168
rect 104450 70048 105250 70168
rect 0 65968 800 66088
rect 104450 65968 105250 66088
rect 0 61888 800 62008
rect 104450 61888 105250 62008
rect 0 57808 800 57928
rect 104450 57808 105250 57928
rect 104450 53728 105250 53848
rect 0 53048 800 53168
rect 0 48968 800 49088
rect 104450 48968 105250 49088
rect 0 44888 800 45008
rect 104450 44888 105250 45008
rect 0 40808 800 40928
rect 104450 40808 105250 40928
rect 0 36728 800 36848
rect 104450 36728 105250 36848
rect 0 32648 800 32768
rect 104450 32648 105250 32768
rect 0 28568 800 28688
rect 104450 28568 105250 28688
rect 0 24488 800 24608
rect 104450 24488 105250 24608
rect 0 20408 800 20528
rect 104450 20408 105250 20528
rect 0 16328 800 16448
rect 104450 16328 105250 16448
rect 0 12248 800 12368
rect 104450 12248 105250 12368
rect 0 8168 800 8288
rect 104450 8168 105250 8288
rect 0 4088 800 4208
rect 104450 4088 105250 4208
rect 104450 8 105250 128
<< obsm3 >>
rect 880 106688 104450 106861
rect 800 102888 104450 106688
rect 880 102608 104370 102888
rect 800 98808 104450 102608
rect 880 98528 104370 98808
rect 800 94728 104450 98528
rect 880 94448 104370 94728
rect 800 90648 104450 94448
rect 880 90368 104370 90648
rect 800 86568 104450 90368
rect 880 86288 104370 86568
rect 800 82488 104450 86288
rect 880 82208 104370 82488
rect 800 78408 104450 82208
rect 880 78128 104370 78408
rect 800 74328 104450 78128
rect 880 74048 104370 74328
rect 800 70248 104450 74048
rect 880 69968 104370 70248
rect 800 66168 104450 69968
rect 880 65888 104370 66168
rect 800 62088 104450 65888
rect 880 61808 104370 62088
rect 800 58008 104450 61808
rect 880 57728 104370 58008
rect 800 53928 104450 57728
rect 800 53648 104370 53928
rect 800 53248 104450 53648
rect 880 52968 104450 53248
rect 800 49168 104450 52968
rect 880 48888 104370 49168
rect 800 45088 104450 48888
rect 880 44808 104370 45088
rect 800 41008 104450 44808
rect 880 40728 104370 41008
rect 800 36928 104450 40728
rect 880 36648 104370 36928
rect 800 32848 104450 36648
rect 880 32568 104370 32848
rect 800 28768 104450 32568
rect 880 28488 104370 28768
rect 800 24688 104450 28488
rect 880 24408 104370 24688
rect 800 20608 104450 24408
rect 880 20328 104370 20608
rect 800 16528 104450 20328
rect 880 16248 104370 16528
rect 800 12448 104450 16248
rect 880 12168 104370 12448
rect 800 8368 104450 12168
rect 880 8088 104370 8368
rect 800 4288 104450 8088
rect 880 4008 104370 4288
rect 800 208 104450 4008
rect 800 35 104370 208
<< metal4 >>
rect 4208 2128 4528 105040
rect 19568 2128 19888 105040
rect 34928 2128 35248 105040
rect 50288 2128 50608 105040
rect 65648 2128 65968 105040
rect 81008 2128 81328 105040
rect 96368 2128 96688 105040
<< obsm4 >>
rect 3923 2048 4128 104685
rect 4608 2048 19488 104685
rect 19968 2048 34848 104685
rect 35328 2048 50208 104685
rect 50688 2048 65568 104685
rect 66048 2048 80928 104685
rect 81408 2048 96288 104685
rect 96768 2048 100405 104685
rect 3923 1667 100405 2048
<< labels >>
rlabel metal2 s 11610 106594 11666 107394 6 clk
port 1 nsew signal input
rlabel metal2 s 93398 0 93454 800 6 ext_address[0]
port 2 nsew signal output
rlabel metal3 s 104450 86368 105250 86488 6 ext_address[10]
port 3 nsew signal output
rlabel metal3 s 0 61888 800 62008 6 ext_address[11]
port 4 nsew signal output
rlabel metal3 s 0 70048 800 70168 6 ext_address[12]
port 5 nsew signal output
rlabel metal2 s 66350 106594 66406 107394 6 ext_address[13]
port 6 nsew signal output
rlabel metal2 s 77942 106594 77998 107394 6 ext_address[14]
port 7 nsew signal output
rlabel metal3 s 0 8168 800 8288 6 ext_address[15]
port 8 nsew signal output
rlabel metal3 s 0 48968 800 49088 6 ext_address[16]
port 9 nsew signal output
rlabel metal3 s 104450 74128 105250 74248 6 ext_address[17]
port 10 nsew signal output
rlabel metal3 s 104450 57808 105250 57928 6 ext_address[18]
port 11 nsew signal output
rlabel metal3 s 104450 4088 105250 4208 6 ext_address[19]
port 12 nsew signal output
rlabel metal3 s 0 82288 800 82408 6 ext_address[1]
port 13 nsew signal output
rlabel metal2 s 66350 0 66406 800 6 ext_address[20]
port 14 nsew signal output
rlabel metal2 s 89534 0 89590 800 6 ext_address[21]
port 15 nsew signal output
rlabel metal3 s 104450 24488 105250 24608 6 ext_address[22]
port 16 nsew signal output
rlabel metal2 s 54758 106594 54814 107394 6 ext_address[23]
port 17 nsew signal output
rlabel metal3 s 0 90448 800 90568 6 ext_address[24]
port 18 nsew signal output
rlabel metal2 s 30930 106594 30986 107394 6 ext_address[25]
port 19 nsew signal output
rlabel metal3 s 104450 98608 105250 98728 6 ext_address[26]
port 20 nsew signal output
rlabel metal2 s 62486 106594 62542 107394 6 ext_address[27]
port 21 nsew signal output
rlabel metal3 s 104450 20408 105250 20528 6 ext_address[28]
port 22 nsew signal output
rlabel metal3 s 0 57808 800 57928 6 ext_address[29]
port 23 nsew signal output
rlabel metal2 s 42522 0 42578 800 6 ext_address[2]
port 24 nsew signal output
rlabel metal3 s 0 36728 800 36848 6 ext_address[30]
port 25 nsew signal output
rlabel metal3 s 104450 16328 105250 16448 6 ext_address[31]
port 26 nsew signal output
rlabel metal2 s 74078 106594 74134 107394 6 ext_address[3]
port 27 nsew signal output
rlabel metal3 s 0 74128 800 74248 6 ext_address[4]
port 28 nsew signal output
rlabel metal2 s 23202 0 23258 800 6 ext_address[5]
port 29 nsew signal output
rlabel metal3 s 0 4088 800 4208 6 ext_address[6]
port 30 nsew signal output
rlabel metal2 s 97262 106594 97318 107394 6 ext_address[7]
port 31 nsew signal output
rlabel metal2 s 11610 0 11666 800 6 ext_address[8]
port 32 nsew signal output
rlabel metal3 s 0 20408 800 20528 6 ext_address[9]
port 33 nsew signal output
rlabel metal2 s 104990 106594 105046 107394 6 ext_instruction
port 34 nsew signal output
rlabel metal2 s 85670 106594 85726 107394 6 ext_read_data[0]
port 35 nsew signal input
rlabel metal3 s 104450 90448 105250 90568 6 ext_read_data[10]
port 36 nsew signal input
rlabel metal3 s 104450 102688 105250 102808 6 ext_read_data[11]
port 37 nsew signal input
rlabel metal3 s 104450 44888 105250 45008 6 ext_read_data[12]
port 38 nsew signal input
rlabel metal3 s 104450 36728 105250 36848 6 ext_read_data[13]
port 39 nsew signal input
rlabel metal2 s 34794 106594 34850 107394 6 ext_read_data[14]
port 40 nsew signal input
rlabel metal2 s 38658 106594 38714 107394 6 ext_read_data[15]
port 41 nsew signal input
rlabel metal3 s 104450 82288 105250 82408 6 ext_read_data[16]
port 42 nsew signal input
rlabel metal2 s 50250 106594 50306 107394 6 ext_read_data[17]
port 43 nsew signal input
rlabel metal2 s 27066 0 27122 800 6 ext_read_data[18]
port 44 nsew signal input
rlabel metal2 s 42522 106594 42578 107394 6 ext_read_data[19]
port 45 nsew signal input
rlabel metal3 s 104450 8 105250 128 6 ext_read_data[1]
port 46 nsew signal input
rlabel metal2 s 58622 106594 58678 107394 6 ext_read_data[20]
port 47 nsew signal input
rlabel metal3 s 0 78208 800 78328 6 ext_read_data[21]
port 48 nsew signal input
rlabel metal2 s 27066 106594 27122 107394 6 ext_read_data[22]
port 49 nsew signal input
rlabel metal3 s 104450 8168 105250 8288 6 ext_read_data[23]
port 50 nsew signal input
rlabel metal3 s 104450 94528 105250 94648 6 ext_read_data[24]
port 51 nsew signal input
rlabel metal2 s 89534 106594 89590 107394 6 ext_read_data[25]
port 52 nsew signal input
rlabel metal2 s 77942 0 77998 800 6 ext_read_data[26]
port 53 nsew signal input
rlabel metal2 s 38658 0 38714 800 6 ext_read_data[27]
port 54 nsew signal input
rlabel metal3 s 104450 28568 105250 28688 6 ext_read_data[28]
port 55 nsew signal input
rlabel metal3 s 0 40808 800 40928 6 ext_read_data[29]
port 56 nsew signal input
rlabel metal3 s 0 53048 800 53168 6 ext_read_data[2]
port 57 nsew signal input
rlabel metal2 s 101126 0 101182 800 6 ext_read_data[30]
port 58 nsew signal input
rlabel metal2 s 19338 106594 19394 107394 6 ext_read_data[31]
port 59 nsew signal input
rlabel metal2 s 81806 0 81862 800 6 ext_read_data[3]
port 60 nsew signal input
rlabel metal3 s 0 98608 800 98728 6 ext_read_data[4]
port 61 nsew signal input
rlabel metal3 s 0 16328 800 16448 6 ext_read_data[5]
port 62 nsew signal input
rlabel metal2 s 7746 0 7802 800 6 ext_read_data[6]
port 63 nsew signal input
rlabel metal2 s 30930 0 30986 800 6 ext_read_data[7]
port 64 nsew signal input
rlabel metal2 s 97262 0 97318 800 6 ext_read_data[8]
port 65 nsew signal input
rlabel metal3 s 104450 53728 105250 53848 6 ext_read_data[9]
port 66 nsew signal input
rlabel metal3 s 104450 32648 105250 32768 6 ext_ready
port 67 nsew signal input
rlabel metal2 s 74078 0 74134 800 6 ext_valid
port 68 nsew signal output
rlabel metal3 s 0 86368 800 86488 6 ext_write_data[0]
port 69 nsew signal output
rlabel metal3 s 0 65968 800 66088 6 ext_write_data[10]
port 70 nsew signal output
rlabel metal3 s 0 24488 800 24608 6 ext_write_data[11]
port 71 nsew signal output
rlabel metal3 s 104450 40808 105250 40928 6 ext_write_data[12]
port 72 nsew signal output
rlabel metal3 s 104450 70048 105250 70168 6 ext_write_data[13]
port 73 nsew signal output
rlabel metal2 s 85670 0 85726 800 6 ext_write_data[14]
port 74 nsew signal output
rlabel metal3 s 104450 78208 105250 78328 6 ext_write_data[15]
port 75 nsew signal output
rlabel metal2 s 50250 0 50306 800 6 ext_write_data[16]
port 76 nsew signal output
rlabel metal3 s 0 106768 800 106888 6 ext_write_data[17]
port 77 nsew signal output
rlabel metal3 s 0 44888 800 45008 6 ext_write_data[18]
port 78 nsew signal output
rlabel metal2 s 18 0 74 800 6 ext_write_data[19]
port 79 nsew signal output
rlabel metal2 s 62486 0 62542 800 6 ext_write_data[1]
port 80 nsew signal output
rlabel metal2 s 15474 106594 15530 107394 6 ext_write_data[20]
port 81 nsew signal output
rlabel metal2 s 46386 106594 46442 107394 6 ext_write_data[21]
port 82 nsew signal output
rlabel metal3 s 0 12248 800 12368 6 ext_write_data[22]
port 83 nsew signal output
rlabel metal3 s 0 102688 800 102808 6 ext_write_data[23]
port 84 nsew signal output
rlabel metal2 s 15474 0 15530 800 6 ext_write_data[24]
port 85 nsew signal output
rlabel metal2 s 3882 0 3938 800 6 ext_write_data[25]
port 86 nsew signal output
rlabel metal2 s 93398 106594 93454 107394 6 ext_write_data[26]
port 87 nsew signal output
rlabel metal2 s 70214 106594 70270 107394 6 ext_write_data[27]
port 88 nsew signal output
rlabel metal2 s 46386 0 46442 800 6 ext_write_data[28]
port 89 nsew signal output
rlabel metal2 s 101126 106594 101182 107394 6 ext_write_data[29]
port 90 nsew signal output
rlabel metal3 s 104450 12248 105250 12368 6 ext_write_data[2]
port 91 nsew signal output
rlabel metal2 s 3882 106594 3938 107394 6 ext_write_data[30]
port 92 nsew signal output
rlabel metal3 s 104450 61888 105250 62008 6 ext_write_data[31]
port 93 nsew signal output
rlabel metal2 s 19338 0 19394 800 6 ext_write_data[3]
port 94 nsew signal output
rlabel metal2 s 34794 0 34850 800 6 ext_write_data[4]
port 95 nsew signal output
rlabel metal2 s 54758 0 54814 800 6 ext_write_data[5]
port 96 nsew signal output
rlabel metal3 s 104450 65968 105250 66088 6 ext_write_data[6]
port 97 nsew signal output
rlabel metal2 s 58622 0 58678 800 6 ext_write_data[7]
port 98 nsew signal output
rlabel metal3 s 0 28568 800 28688 6 ext_write_data[8]
port 99 nsew signal output
rlabel metal2 s 81806 106594 81862 107394 6 ext_write_data[9]
port 100 nsew signal output
rlabel metal2 s 7746 106594 7802 107394 6 ext_write_strobe[0]
port 101 nsew signal output
rlabel metal2 s 23202 106594 23258 107394 6 ext_write_strobe[1]
port 102 nsew signal output
rlabel metal2 s 70214 0 70270 800 6 ext_write_strobe[2]
port 103 nsew signal output
rlabel metal3 s 0 32648 800 32768 6 ext_write_strobe[3]
port 104 nsew signal output
rlabel metal3 s 0 94528 800 94648 6 meip
port 105 nsew signal input
rlabel metal3 s 104450 48968 105250 49088 6 reset
port 106 nsew signal input
rlabel metal4 s 4208 2128 4528 105040 6 vccd1
port 107 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 105040 6 vccd1
port 107 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 105040 6 vccd1
port 107 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 105040 6 vccd1
port 107 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 105040 6 vssd1
port 108 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 105040 6 vssd1
port 108 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 105040 6 vssd1
port 108 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 105250 107394
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 33314604
string GDS_FILE /data/yinguohua/Cyberrio/openlane/user_proj_example/runs/23_06_02_18_23/results/signoff/core.magic.gds
string GDS_START 1318596
<< end >>

