* NGSPICE file created from core.ext - technology: sky130A

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_8 abstract view
.subckt sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_2 abstract view
.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_8 abstract view
.subckt sky130_fd_sc_hd__mux2_8 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_4 abstract view
.subckt sky130_fd_sc_hd__and4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_4 abstract view
.subckt sky130_fd_sc_hd__a22o_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_2 abstract view
.subckt sky130_fd_sc_hd__and4b_2 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_2 abstract view
.subckt sky130_fd_sc_hd__mux4_2 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_4 abstract view
.subckt sky130_fd_sc_hd__o31a_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_2 abstract view
.subckt sky130_fd_sc_hd__o22ai_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_4 abstract view
.subckt sky130_fd_sc_hd__o22a_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_2 abstract view
.subckt sky130_fd_sc_hd__a21bo_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_4 abstract view
.subckt sky130_fd_sc_hd__nand2b_4 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_4 abstract view
.subckt sky130_fd_sc_hd__and3b_4 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_2 abstract view
.subckt sky130_fd_sc_hd__a32o_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_4 abstract view
.subckt sky130_fd_sc_hd__o32a_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_4 abstract view
.subckt sky130_fd_sc_hd__a2111o_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_4 abstract view
.subckt sky130_fd_sc_hd__and4b_4 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_4 abstract view
.subckt sky130_fd_sc_hd__and4bb_4 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_4 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_6 abstract view
.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_1 abstract view
.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_4 abstract view
.subckt sky130_fd_sc_hd__a21boi_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_2 abstract view
.subckt sky130_fd_sc_hd__nand3b_2 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_2 abstract view
.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_2 abstract view
.subckt sky130_fd_sc_hd__o32a_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_4 abstract view
.subckt sky130_fd_sc_hd__a31o_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_4 abstract view
.subckt sky130_fd_sc_hd__nor4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_2 abstract view
.subckt sky130_fd_sc_hd__o221ai_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_4 abstract view
.subckt sky130_fd_sc_hd__a221o_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_4 abstract view
.subckt sky130_fd_sc_hd__o2111a_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_4 abstract view
.subckt sky130_fd_sc_hd__o22ai_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_2 abstract view
.subckt sky130_fd_sc_hd__or4bb_2 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_4 abstract view
.subckt sky130_fd_sc_hd__a221oi_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_4 abstract view
.subckt sky130_fd_sc_hd__and2b_4 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_1 abstract view
.subckt sky130_fd_sc_hd__a2111oi_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_4 abstract view
.subckt sky130_fd_sc_hd__a41o_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__bufbuf_16 abstract view
.subckt sky130_fd_sc_hd__bufbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_8 abstract view
.subckt sky130_fd_sc_hd__inv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_4 abstract view
.subckt sky130_fd_sc_hd__nor3b_4 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_4 abstract view
.subckt sky130_fd_sc_hd__or4bb_4 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_2 abstract view
.subckt sky130_fd_sc_hd__a2111o_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_8 abstract view
.subckt sky130_fd_sc_hd__clkinv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_4 abstract view
.subckt sky130_fd_sc_hd__nand3b_4 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_4 abstract view
.subckt sky130_fd_sc_hd__nand4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_4 abstract view
.subckt sky130_fd_sc_hd__o221ai_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

.subckt core clk ext_address[0] ext_address[10] ext_address[11] ext_address[12] ext_address[13]
+ ext_address[14] ext_address[15] ext_address[16] ext_address[17] ext_address[18]
+ ext_address[19] ext_address[1] ext_address[20] ext_address[21] ext_address[22] ext_address[23]
+ ext_address[24] ext_address[25] ext_address[26] ext_address[27] ext_address[28]
+ ext_address[29] ext_address[2] ext_address[30] ext_address[31] ext_address[3] ext_address[4]
+ ext_address[5] ext_address[6] ext_address[7] ext_address[8] ext_address[9] ext_instruction
+ ext_read_data[0] ext_read_data[10] ext_read_data[11] ext_read_data[12] ext_read_data[13]
+ ext_read_data[14] ext_read_data[15] ext_read_data[16] ext_read_data[17] ext_read_data[18]
+ ext_read_data[19] ext_read_data[1] ext_read_data[20] ext_read_data[21] ext_read_data[22]
+ ext_read_data[23] ext_read_data[24] ext_read_data[25] ext_read_data[26] ext_read_data[27]
+ ext_read_data[28] ext_read_data[29] ext_read_data[2] ext_read_data[30] ext_read_data[31]
+ ext_read_data[3] ext_read_data[4] ext_read_data[5] ext_read_data[6] ext_read_data[7]
+ ext_read_data[8] ext_read_data[9] ext_ready ext_valid ext_write_data[0] ext_write_data[10]
+ ext_write_data[11] ext_write_data[12] ext_write_data[13] ext_write_data[14] ext_write_data[15]
+ ext_write_data[16] ext_write_data[17] ext_write_data[18] ext_write_data[19] ext_write_data[1]
+ ext_write_data[20] ext_write_data[21] ext_write_data[22] ext_write_data[23] ext_write_data[24]
+ ext_write_data[25] ext_write_data[26] ext_write_data[27] ext_write_data[28] ext_write_data[29]
+ ext_write_data[2] ext_write_data[30] ext_write_data[31] ext_write_data[3] ext_write_data[4]
+ ext_write_data[5] ext_write_data[6] ext_write_data[7] ext_write_data[8] ext_write_data[9]
+ ext_write_strobe[0] ext_write_strobe[1] ext_write_strobe[2] ext_write_strobe[3]
+ meip reset vccd1 vssd1
XFILLER_79_380 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_127 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09671_ _14042_/Q _13326_/A0 _09690_/S vssd1 vssd1 vccd1 vccd1 _14042_/D sky130_fd_sc_hd__mux2_1
X_06883_ _15399_/Q _06688_/Y _15398_/Q _06691_/Y vssd1 vssd1 vccd1 vccd1 _06883_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_39_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08622_ _13463_/Q _08684_/A2 _08691_/A2 _13598_/Q _08621_/X vssd1 vssd1 vccd1 vccd1
+ _08622_/X sky130_fd_sc_hd__a221o_1
XFILLER_82_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08553_ _13777_/Q _08573_/S _08552_/X vssd1 vssd1 vccd1 vccd1 _13777_/D sky130_fd_sc_hd__o21a_1
XFILLER_82_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07504_ _07783_/A _07504_/B _07504_/C vssd1 vssd1 vccd1 vccd1 _08025_/C sky130_fd_sc_hd__or3_1
X_08484_ _14592_/Q _08465_/B _08487_/B _09435_/A vssd1 vssd1 vccd1 vccd1 _08484_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_51_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07435_ _13664_/Q _07483_/A2 _07483_/B1 _14692_/Q _07434_/X vssd1 vssd1 vccd1 vccd1
+ _07435_/X sky130_fd_sc_hd__a221o_1
XFILLER_168_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07366_ _14716_/Q _08817_/B vssd1 vssd1 vccd1 vccd1 _13318_/C sky130_fd_sc_hd__nand2_8
XFILLER_148_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09105_ _13949_/Q _13691_/Q _09425_/S vssd1 vssd1 vccd1 vccd1 _09105_/X sky130_fd_sc_hd__mux2_1
XFILLER_149_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07297_ _07297_/A vssd1 vssd1 vccd1 vccd1 _07297_/Y sky130_fd_sc_hd__inv_2
XFILLER_164_845 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09036_ _13913_/Q _13139_/S _09035_/X vssd1 vssd1 vccd1 vccd1 _13913_/D sky130_fd_sc_hd__a21o_1
XFILLER_164_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09938_ _11858_/A1 _14298_/Q _09958_/S vssd1 vssd1 vccd1 vccd1 _14298_/D sky130_fd_sc_hd__mux2_1
XFILLER_89_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09869_ _11680_/A0 _14231_/Q _09892_/S vssd1 vssd1 vccd1 vccd1 _14231_/D sky130_fd_sc_hd__mux2_1
XFILLER_92_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11900_ _12268_/A _11900_/B vssd1 vssd1 vccd1 vccd1 _11900_/X sky130_fd_sc_hd__and2_1
XTAP_3235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12880_ _15408_/Q _15593_/Q _12918_/S vssd1 vssd1 vccd1 vccd1 _15408_/D sky130_fd_sc_hd__mux2_1
XFILLER_45_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_172_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11831_ _15253_/Q _13331_/A0 _11849_/S vssd1 vssd1 vccd1 vccd1 _15253_/D sky130_fd_sc_hd__mux2_1
XTAP_2534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14550_ _15209_/CLK _14550_/D vssd1 vssd1 vccd1 vccd1 _14550_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_228 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11762_ _11870_/A1 _15190_/Q _11775_/S vssd1 vssd1 vccd1 vccd1 _15190_/D sky130_fd_sc_hd__mux2_1
XFILLER_26_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13501_ _13565_/CLK _13501_/D vssd1 vssd1 vccd1 vccd1 _13501_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_14_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10713_ _15038_/Q _10652_/B _10712_/X vssd1 vssd1 vccd1 vccd1 _10713_/X sky130_fd_sc_hd__a21o_1
XTAP_1877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14481_ _15300_/CLK _14481_/D vssd1 vssd1 vccd1 vccd1 _14481_/Q sky130_fd_sc_hd__dfxtp_1
X_11693_ _13335_/A0 _15124_/Q _11703_/S vssd1 vssd1 vccd1 vccd1 _15124_/D sky130_fd_sc_hd__mux2_1
XTAP_1899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13432_ _15389_/CLK _13432_/D vssd1 vssd1 vccd1 vccd1 _13432_/Q sky130_fd_sc_hd__dfxtp_2
X_10644_ _15056_/Q _10714_/A2 _10641_/X _10643_/X vssd1 vssd1 vccd1 vccd1 _10644_/X
+ sky130_fd_sc_hd__o22a_2
XFILLER_127_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13363_ _14466_/Q vssd1 vssd1 vccd1 vccd1 _14466_/D sky130_fd_sc_hd__clkbuf_2
X_10575_ _14929_/Q _10581_/B _14927_/Q vssd1 vssd1 vccd1 vccd1 _10575_/X sky130_fd_sc_hd__and3_2
X_15102_ _15675_/CLK _15102_/D vssd1 vssd1 vccd1 vccd1 _15102_/Q sky130_fd_sc_hd__dfxtp_1
X_12314_ _12383_/A _12314_/B vssd1 vssd1 vccd1 vccd1 _12314_/X sky130_fd_sc_hd__and2_1
XFILLER_127_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13294_ _12681_/Y _15626_/Q _13300_/S vssd1 vssd1 vccd1 vccd1 _15626_/D sky130_fd_sc_hd__mux2_1
XFILLER_138_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15033_ _15041_/CLK _15033_/D vssd1 vssd1 vccd1 vccd1 _15033_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_154_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12245_ _12452_/A _12245_/B vssd1 vssd1 vccd1 vccd1 _12245_/X sky130_fd_sc_hd__and2_1
XFILLER_107_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12176_ _12452_/A _12176_/B vssd1 vssd1 vccd1 vccd1 _12176_/X sky130_fd_sc_hd__and2_1
XFILLER_174_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11127_ _11414_/A _11185_/B _11126_/X _11202_/A vssd1 vssd1 vccd1 vccd1 _11127_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_68_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_593 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11058_ _11058_/A vssd1 vssd1 vccd1 vccd1 _11058_/Y sky130_fd_sc_hd__inv_2
XFILLER_95_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10009_ _13330_/A0 _14367_/Q _10028_/S vssd1 vssd1 vccd1 vccd1 _14367_/D sky130_fd_sc_hd__mux2_1
XFILLER_49_586 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14817_ _15643_/CLK _14817_/D vssd1 vssd1 vccd1 vccd1 _14817_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14748_ _15569_/CLK _14748_/D vssd1 vssd1 vccd1 vccd1 _14748_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_33_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14679_ _15619_/CLK _14679_/D vssd1 vssd1 vccd1 vccd1 _14679_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07220_ _15330_/Q _15486_/Q _07340_/S vssd1 vssd1 vccd1 vccd1 _07221_/A sky130_fd_sc_hd__mux2_8
XFILLER_177_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_108 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07151_ _07163_/A _07151_/B vssd1 vssd1 vccd1 vccd1 _07151_/X sky130_fd_sc_hd__and2_4
XFILLER_145_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07082_ _07081_/X _13606_/Q _12662_/S vssd1 vssd1 vccd1 vccd1 _07082_/X sky130_fd_sc_hd__mux2_1
XFILLER_172_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout105 _12621_/Y vssd1 vssd1 vccd1 vccd1 _12743_/A sky130_fd_sc_hd__buf_12
XFILLER_141_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout116 _12946_/Y vssd1 vssd1 vccd1 vccd1 _13116_/C sky130_fd_sc_hd__buf_8
XFILLER_99_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout127 fanout138/X vssd1 vssd1 vccd1 vccd1 _13140_/S sky130_fd_sc_hd__buf_6
Xfanout138 _06782_/Y vssd1 vssd1 vccd1 vccd1 fanout138/X sky130_fd_sc_hd__buf_12
XFILLER_102_948 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout149 _12885_/S vssd1 vssd1 vccd1 vccd1 _12906_/S sky130_fd_sc_hd__buf_12
X_07984_ _13562_/Q _13561_/Q _13560_/Q _07984_/D vssd1 vssd1 vccd1 vccd1 _07995_/D
+ sky130_fd_sc_hd__and4_2
XFILLER_68_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09723_ _13104_/B2 _14093_/Q _09723_/S vssd1 vssd1 vccd1 vccd1 _14093_/D sky130_fd_sc_hd__mux2_1
X_06935_ _14501_/Q _06936_/B _14500_/Q _06724_/Y vssd1 vssd1 vccd1 vccd1 _06941_/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_74_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09654_ _14027_/Q _11876_/A1 _09660_/S vssd1 vssd1 vccd1 vccd1 _14027_/D sky130_fd_sc_hd__mux2_1
XFILLER_27_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06866_ _06873_/B _14514_/Q _13506_/Q _06692_/Y vssd1 vssd1 vccd1 vccd1 _06882_/A
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_103_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08605_ _08722_/A _08605_/B _08605_/C vssd1 vssd1 vccd1 vccd1 _08605_/X sky130_fd_sc_hd__or3_1
XFILLER_103_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09585_ _13961_/Q _13341_/A0 _09589_/S vssd1 vssd1 vccd1 vccd1 _13961_/D sky130_fd_sc_hd__mux2_1
X_06797_ _06797_/A vssd1 vssd1 vccd1 vccd1 _06797_/Y sky130_fd_sc_hd__inv_2
XFILLER_103_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08536_ _08536_/A _08536_/B _08536_/C vssd1 vssd1 vccd1 vccd1 _08538_/B sky130_fd_sc_hd__or3_4
XFILLER_179_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08467_ hold5/A _09829_/B _06988_/A _08490_/A1 _08466_/X vssd1 vssd1 vccd1 vccd1
+ _08467_/X sky130_fd_sc_hd__a221o_2
XFILLER_23_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07418_ _14656_/Q _07474_/B _07482_/C vssd1 vssd1 vccd1 vccd1 _07418_/X sky130_fd_sc_hd__and3_1
X_08398_ _13732_/Q _13140_/S _08394_/X _14591_/Q vssd1 vssd1 vccd1 vccd1 _13732_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_183_428 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07349_ _07306_/Y _07307_/X _07278_/X vssd1 vssd1 vccd1 vccd1 _07350_/D sky130_fd_sc_hd__a21oi_1
XFILLER_109_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10360_ _10360_/A _10360_/B vssd1 vssd1 vccd1 vccd1 _10360_/X sky130_fd_sc_hd__and2_2
XFILLER_12_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09019_ _08507_/A _09018_/X _09017_/X _09524_/A vssd1 vssd1 vccd1 vccd1 _09019_/X
+ sky130_fd_sc_hd__o211a_1
X_10291_ _14676_/Q _14829_/Q _10735_/S vssd1 vssd1 vccd1 vccd1 _14676_/D sky130_fd_sc_hd__mux2_1
XFILLER_128_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12030_ _12582_/A _12030_/B vssd1 vssd1 vccd1 vccd1 _12030_/X sky130_fd_sc_hd__or2_1
XFILLER_2_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13981_ _15133_/CLK _13981_/D vssd1 vssd1 vccd1 vccd1 _13981_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_77_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12932_ _15460_/Q _15646_/Q _12932_/S vssd1 vssd1 vccd1 vccd1 _15460_/D sky130_fd_sc_hd__mux2_1
XTAP_3021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15651_ _15651_/CLK _15651_/D vssd1 vssd1 vccd1 vccd1 _15651_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12863_ _14757_/Q _15391_/Q _12866_/S vssd1 vssd1 vccd1 vccd1 _15391_/D sky130_fd_sc_hd__mux2_1
XTAP_3065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14602_ _14892_/CLK _14602_/D vssd1 vssd1 vccd1 vccd1 _14602_/Q sky130_fd_sc_hd__dfxtp_1
X_11814_ _15237_/Q _11847_/A1 _11817_/S vssd1 vssd1 vccd1 vccd1 _15237_/D sky130_fd_sc_hd__mux2_1
XTAP_2364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15582_ _15582_/CLK _15582_/D vssd1 vssd1 vccd1 vccd1 _15582_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12794_ _06861_/Y _12791_/Y _12792_/X _12793_/X vssd1 vssd1 vccd1 vccd1 _12794_/X
+ sky130_fd_sc_hd__a31o_1
XTAP_1641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_712 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14533_ _15315_/CLK _14533_/D vssd1 vssd1 vccd1 vccd1 _14533_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11745_ _11853_/A1 _15173_/Q _11775_/S vssd1 vssd1 vccd1 vccd1 _15173_/D sky130_fd_sc_hd__mux2_1
XFILLER_18_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_795 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14464_ _15556_/CLK _14464_/D vssd1 vssd1 vccd1 vccd1 _14464_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_174_406 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11676_ _14714_/Q _14715_/Q _13318_/C _11851_/A vssd1 vssd1 vccd1 vccd1 _11676_/X
+ sky130_fd_sc_hd__or4_4
XFILLER_144_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13415_ _13803_/CLK _13415_/D vssd1 vssd1 vccd1 vccd1 _13415_/Q sky130_fd_sc_hd__dfxtp_1
X_10627_ _15004_/Q _10717_/A2 _10652_/B _13723_/Q _10717_/C1 vssd1 vssd1 vccd1 vccd1
+ _10627_/X sky130_fd_sc_hd__a221o_1
XFILLER_139_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14395_ _15081_/CLK _14395_/D vssd1 vssd1 vccd1 vccd1 _14395_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_973 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13346_ _13346_/A0 _15676_/Q _13350_/S vssd1 vssd1 vccd1 vccd1 _15676_/D sky130_fd_sc_hd__mux2_1
XFILLER_127_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10558_ _10558_/A _10558_/B _10558_/C vssd1 vssd1 vccd1 vccd1 _11240_/A sky130_fd_sc_hd__nor3_2
XFILLER_183_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13277_ _15361_/Q _15608_/Q _13300_/S vssd1 vssd1 vccd1 vccd1 _15608_/D sky130_fd_sc_hd__mux2_1
XFILLER_170_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10489_ _11561_/A _11563_/A vssd1 vssd1 vccd1 vccd1 _10491_/A sky130_fd_sc_hd__or2_1
X_15016_ _15017_/CLK _15016_/D vssd1 vssd1 vccd1 vccd1 _15016_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_170_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12228_ _12504_/A _12228_/B _12228_/C vssd1 vssd1 vccd1 vccd1 _12228_/X sky130_fd_sc_hd__and3_1
XFILLER_123_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_572 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12159_ _12596_/A _12159_/B _12159_/C vssd1 vssd1 vccd1 vccd1 _12159_/X sky130_fd_sc_hd__and3_1
XFILLER_123_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_1027 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06720_ _14502_/Q vssd1 vssd1 vccd1 vccd1 _06720_/Y sky130_fd_sc_hd__inv_2
XFILLER_80_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_206 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09370_ _14379_/Q _15195_/Q _13834_/Q _14573_/Q _09535_/S _08494_/B vssd1 vssd1 vccd1
+ vccd1 _09371_/B sky130_fd_sc_hd__mux4_1
XFILLER_178_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08321_ _11283_/A _08319_/X _08320_/Y _10403_/A vssd1 vssd1 vccd1 vccd1 _08321_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_71_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_1039 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08252_ _11351_/C1 _10895_/B _11437_/A _08224_/X vssd1 vssd1 vccd1 vccd1 _13713_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_32_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07203_ _15334_/Q _15490_/Q _07335_/S vssd1 vssd1 vccd1 vccd1 _07204_/A sky130_fd_sc_hd__mux2_8
X_08183_ _08150_/S input24/X _08185_/A vssd1 vssd1 vccd1 vccd1 _08183_/X sky130_fd_sc_hd__and3b_1
XFILLER_146_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_4_12_0_clk clkbuf_3_6_0_clk/X vssd1 vssd1 vccd1 vccd1 clkbuf_5_25_0_clk/A
+ sky130_fd_sc_hd__clkbuf_8
X_07134_ _14847_/Q _14839_/Q _07146_/S vssd1 vssd1 vccd1 vccd1 _07134_/X sky130_fd_sc_hd__mux2_1
XFILLER_119_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07065_ _07064_/X _14754_/Q _07077_/S vssd1 vssd1 vccd1 vccd1 _13600_/D sky130_fd_sc_hd__mux2_1
XFILLER_160_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07967_ _13557_/Q _07973_/D vssd1 vssd1 vccd1 vccd1 _07967_/X sky130_fd_sc_hd__or2_1
X_09706_ _13328_/A0 _14076_/Q _09723_/S vssd1 vssd1 vccd1 vccd1 _14076_/D sky130_fd_sc_hd__mux2_1
X_06918_ _06918_/A _13468_/Q vssd1 vssd1 vccd1 vccd1 _06918_/X sky130_fd_sc_hd__or2_1
X_07898_ _07903_/A _07898_/B vssd1 vssd1 vccd1 vccd1 _07898_/Y sky130_fd_sc_hd__nand2_1
X_09637_ _14010_/Q _13326_/A0 _09660_/S vssd1 vssd1 vccd1 vccd1 _14010_/D sky130_fd_sc_hd__mux2_1
XFILLER_83_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06849_ _14906_/Q _06848_/X _06682_/Y _14923_/Q _06847_/X vssd1 vssd1 vccd1 vccd1
+ _06849_/X sky130_fd_sc_hd__o2111a_1
XFILLER_28_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_183 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09568_ _13944_/Q _11649_/A0 _09594_/S vssd1 vssd1 vccd1 vccd1 _13944_/D sky130_fd_sc_hd__mux2_1
X_08519_ _08519_/A _08519_/B vssd1 vssd1 vccd1 vccd1 _08519_/X sky130_fd_sc_hd__and2_4
X_09499_ _14257_/Q _14289_/Q _14321_/Q _14353_/Q _09535_/S _08494_/B vssd1 vssd1 vccd1
+ vccd1 _09499_/X sky130_fd_sc_hd__mux4_1
XFILLER_168_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11530_ _13215_/B _11532_/B vssd1 vssd1 vccd1 vccd1 _11530_/X sky130_fd_sc_hd__and2_1
XFILLER_168_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11461_ _11440_/A _11440_/B _11450_/B vssd1 vssd1 vccd1 vccd1 _11461_/X sky130_fd_sc_hd__a21bo_1
XFILLER_168_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13200_ _13217_/A _13199_/B _11496_/A vssd1 vssd1 vccd1 vccd1 _13200_/Y sky130_fd_sc_hd__a21oi_1
X_10412_ _11414_/C _11399_/A _10395_/A vssd1 vssd1 vccd1 vccd1 _10412_/X sky130_fd_sc_hd__or3b_1
X_14180_ _14225_/CLK _14180_/D vssd1 vssd1 vccd1 vccd1 _14180_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_104_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11392_ _11401_/B _11401_/C vssd1 vssd1 vccd1 vccd1 _11394_/A sky130_fd_sc_hd__nand2_1
XFILLER_136_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_600 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13131_ _13131_/A _14610_/Q _13131_/C vssd1 vssd1 vccd1 vccd1 _13131_/Y sky130_fd_sc_hd__nor3_1
XFILLER_136_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10343_ _14728_/Q _14921_/Q _10343_/S vssd1 vssd1 vccd1 vccd1 _14728_/D sky130_fd_sc_hd__mux2_1
XFILLER_152_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10274_ _14659_/Q _14812_/Q _10630_/S vssd1 vssd1 vccd1 vccd1 _14659_/D sky130_fd_sc_hd__mux2_1
XFILLER_174_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13062_ _12960_/X _13118_/A2 _13114_/B1 _13324_/A0 vssd1 vssd1 vccd1 vccd1 _13062_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_105_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12013_ _12592_/A1 _12012_/X _12594_/S vssd1 vssd1 vccd1 vccd1 _12013_/X sky130_fd_sc_hd__a21o_1
XFILLER_3_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_opt_2_0_clk clkbuf_5_12_0_clk/X vssd1 vssd1 vccd1 vccd1 clkbuf_opt_2_0_clk/X
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_19_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout480 _12548_/S vssd1 vssd1 vccd1 vccd1 _12559_/A sky130_fd_sc_hd__buf_8
XFILLER_48_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout491 _07104_/C vssd1 vssd1 vccd1 vccd1 _08093_/B sky130_fd_sc_hd__buf_4
X_13964_ _14405_/CLK _13964_/D vssd1 vssd1 vccd1 vccd1 _13964_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12915_ _15443_/Q _15629_/Q _12918_/S vssd1 vssd1 vccd1 vccd1 _15443_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13895_ _15293_/CLK _13895_/D vssd1 vssd1 vccd1 vccd1 _13895_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_111_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15634_ _15634_/CLK _15634_/D vssd1 vssd1 vccd1 vccd1 _15634_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_46_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12846_ _14740_/Q _15374_/Q _12871_/S vssd1 vssd1 vccd1 vccd1 _15374_/D sky130_fd_sc_hd__mux2_1
XFILLER_181_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_520 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15565_ _15569_/CLK _15565_/D vssd1 vssd1 vccd1 vccd1 _15565_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12777_ _12789_/C _12777_/B vssd1 vssd1 vccd1 vccd1 _12778_/B sky130_fd_sc_hd__and2b_1
XFILLER_14_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14516_ _14517_/CLK _14516_/D vssd1 vssd1 vccd1 vccd1 _14516_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11728_ _15157_/Q _13336_/A0 _11742_/S vssd1 vssd1 vccd1 vccd1 _15157_/D sky130_fd_sc_hd__mux2_1
X_15496_ _15523_/CLK _15496_/D vssd1 vssd1 vccd1 vccd1 _15496_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_175_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14447_ _15662_/CLK _14447_/D vssd1 vssd1 vccd1 vccd1 _14447_/Q sky130_fd_sc_hd__dfxtp_1
X_11659_ _13082_/B2 _15091_/Q _11670_/S vssd1 vssd1 vccd1 vccd1 _15091_/D sky130_fd_sc_hd__mux2_1
XFILLER_7_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14378_ _15295_/CLK _14378_/D vssd1 vssd1 vccd1 vccd1 _14378_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_183_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_686 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_994 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13329_ _13329_/A0 _15659_/Q _13345_/S vssd1 vssd1 vccd1 vccd1 _15659_/D sky130_fd_sc_hd__mux2_1
XFILLER_50_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_3_1_0_clk clkbuf_3_1_0_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_3_0_clk/A sky130_fd_sc_hd__clkbuf_8
XFILLER_131_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08870_ _13891_/Q _11868_/A1 _08880_/S vssd1 vssd1 vccd1 vccd1 _13891_/D sky130_fd_sc_hd__mux2_1
XFILLER_96_220 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07821_ _13519_/Q _13518_/Q _07825_/D vssd1 vssd1 vccd1 vccd1 _07821_/X sky130_fd_sc_hd__and3_1
XFILLER_69_467 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07752_ _13501_/Q _07757_/D _13502_/Q vssd1 vssd1 vccd1 vccd1 _07752_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_56_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06703_ _13502_/Q vssd1 vssd1 vccd1 vccd1 _06703_/Y sky130_fd_sc_hd__inv_2
XFILLER_65_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07683_ _13483_/Q _07687_/C vssd1 vssd1 vccd1 vccd1 _07686_/B sky130_fd_sc_hd__and2_1
XFILLER_92_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09422_ _14028_/Q _13996_/Q _09425_/S vssd1 vssd1 vccd1 vccd1 _09422_/X sky130_fd_sc_hd__mux2_1
XFILLER_64_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09353_ _13865_/Q _14218_/Q _09521_/S vssd1 vssd1 vccd1 vccd1 _09353_/X sky130_fd_sc_hd__mux2_1
XFILLER_12_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08304_ _11349_/B _13178_/B vssd1 vssd1 vccd1 vccd1 _11045_/A sky130_fd_sc_hd__nor2_1
X_09284_ _09543_/A _09284_/B vssd1 vssd1 vccd1 vccd1 _09284_/X sky130_fd_sc_hd__or2_1
XFILLER_127_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08235_ _07337_/A _10457_/A2 _08234_/X vssd1 vssd1 vccd1 vccd1 _08235_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_165_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_247 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08166_ _13670_/Q _10695_/S _08155_/X _08165_/X vssd1 vssd1 vccd1 vccd1 _13670_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_118_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07117_ _07131_/A _07117_/B vssd1 vssd1 vccd1 vccd1 _07117_/X sky130_fd_sc_hd__and2_2
XFILLER_134_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08097_ _08093_/Y _08095_/X _08096_/X _10344_/S _13649_/Q vssd1 vssd1 vccd1 vccd1
+ _13649_/D sky130_fd_sc_hd__a32o_1
XFILLER_134_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07048_ _14628_/Q _14660_/Q _07078_/S vssd1 vssd1 vccd1 vccd1 _07048_/X sky130_fd_sc_hd__mux2_1
XFILLER_161_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_1000 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_231 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08999_ _14427_/Q _08540_/B _08520_/B _08998_/X vssd1 vssd1 vccd1 vccd1 _08999_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_134_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10961_ _11023_/A _11626_/A vssd1 vssd1 vccd1 vccd1 _10963_/A sky130_fd_sc_hd__or2_2
XFILLER_44_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12700_ _15348_/Q _12765_/B _12699_/X _12809_/C1 vssd1 vssd1 vccd1 vccd1 _15348_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_71_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13680_ _14892_/CLK _13680_/D vssd1 vssd1 vccd1 vccd1 _13680_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10892_ _13807_/Q _10892_/B _10891_/X vssd1 vssd1 vccd1 vccd1 _10892_/X sky130_fd_sc_hd__or3b_1
X_12631_ _13583_/Q _12630_/X _12785_/B vssd1 vssd1 vccd1 vccd1 _12631_/X sky130_fd_sc_hd__mux2_1
XFILLER_34_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_1083 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15350_ _15630_/CLK _15350_/D vssd1 vssd1 vccd1 vccd1 _15350_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_70_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12562_ _13968_/Q _13710_/Q _12568_/S vssd1 vssd1 vccd1 vccd1 _12563_/B sky130_fd_sc_hd__mux2_1
XFILLER_141_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14301_ _15181_/CLK _14301_/D vssd1 vssd1 vccd1 vccd1 _14301_/Q sky130_fd_sc_hd__dfxtp_1
X_11513_ _11546_/A _11508_/B _11501_/A vssd1 vssd1 vccd1 vccd1 _11516_/A sky130_fd_sc_hd__a21bo_1
XFILLER_156_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_202 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15281_ _15281_/CLK _15281_/D vssd1 vssd1 vccd1 vccd1 _15281_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_156_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12493_ _13965_/Q _13707_/Q _12499_/S vssd1 vssd1 vccd1 vccd1 _12494_/B sky130_fd_sc_hd__mux2_1
X_14232_ _15273_/CLK _14232_/D vssd1 vssd1 vccd1 vccd1 _14232_/Q sky130_fd_sc_hd__dfxtp_1
X_11444_ _11430_/X _11440_/Y _11441_/X _11474_/S vssd1 vssd1 vccd1 vccd1 _11444_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_138_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14163_ _15172_/CLK _14163_/D vssd1 vssd1 vccd1 vccd1 _14163_/Q sky130_fd_sc_hd__dfxtp_1
X_11375_ _13165_/B _11375_/B _11375_/C vssd1 vssd1 vccd1 vccd1 _11377_/B sky130_fd_sc_hd__and3b_1
XFILLER_4_964 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13114_ _13038_/X _13118_/A2 _13114_/B1 _07500_/X vssd1 vssd1 vccd1 vccd1 _13114_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_152_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10326_ _07498_/B _14904_/Q _10730_/S vssd1 vssd1 vccd1 vccd1 _14711_/D sky130_fd_sc_hd__mux2_1
XFILLER_98_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14094_ _15676_/CLK _14094_/D vssd1 vssd1 vccd1 vccd1 _14094_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13045_ _09382_/A _11743_/C _08817_/Y _09466_/A vssd1 vssd1 vccd1 vccd1 _13045_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_140_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10257_ _14642_/Q hold6/X _10610_/S vssd1 vssd1 vccd1 vccd1 _14642_/D sky130_fd_sc_hd__mux2_1
XFILLER_79_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10188_ _11874_/A1 _14572_/Q _10197_/S vssd1 vssd1 vccd1 vccd1 _14572_/D sky130_fd_sc_hd__mux2_1
XFILLER_121_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14996_ _15558_/CLK _14996_/D vssd1 vssd1 vccd1 vccd1 _14996_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_971 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13947_ _15657_/CLK _13947_/D vssd1 vssd1 vccd1 vccd1 _13947_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13878_ _15202_/CLK _13878_/D vssd1 vssd1 vccd1 vccd1 _13878_/Q sky130_fd_sc_hd__dfxtp_1
X_15617_ _15617_/CLK _15617_/D vssd1 vssd1 vccd1 vccd1 _15617_/Q sky130_fd_sc_hd__dfxtp_1
X_12829_ _15073_/Q _12834_/B vssd1 vssd1 vccd1 vccd1 _12829_/X sky130_fd_sc_hd__or2_1
XFILLER_22_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_570 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15548_ _15548_/CLK _15548_/D vssd1 vssd1 vccd1 vccd1 _15548_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_187_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15479_ _15525_/CLK _15479_/D vssd1 vssd1 vccd1 vccd1 _15479_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_150_clk clkbuf_5_25_0_clk/X vssd1 vssd1 vccd1 vccd1 _15618_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_129_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08020_ _08022_/B _08018_/Y _08019_/Y input35/X vssd1 vssd1 vccd1 vccd1 _13571_/D
+ sky130_fd_sc_hd__a211oi_1
XFILLER_163_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_987 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09971_ _11858_/A1 _14330_/Q _09991_/S vssd1 vssd1 vccd1 vccd1 _14330_/D sky130_fd_sc_hd__mux2_1
XFILLER_131_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_272 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08922_ _15650_/Q _13384_/Q _09557_/S vssd1 vssd1 vccd1 vccd1 _08922_/X sky130_fd_sc_hd__mux2_1
XFILLER_130_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08853_ _10032_/A _11851_/A vssd1 vssd1 vccd1 vccd1 _08853_/Y sky130_fd_sc_hd__nor2_8
XFILLER_84_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07804_ _07813_/D _07803_/Y _07816_/A vssd1 vssd1 vccd1 vccd1 _07804_/Y sky130_fd_sc_hd__o21ai_1
XTAP_3609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08784_ _14714_/Q _14716_/Q _11743_/C _13318_/D vssd1 vssd1 vccd1 vccd1 _08784_/X
+ sky130_fd_sc_hd__or4_4
X_07735_ _13497_/Q _07739_/C vssd1 vssd1 vccd1 vccd1 _07736_/B sky130_fd_sc_hd__xnor2_1
XFILLER_26_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07666_ _07664_/Y _07672_/C _07777_/A vssd1 vssd1 vccd1 vccd1 _07666_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_164_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09405_ _09405_/A _09405_/B _09405_/C vssd1 vssd1 vccd1 vccd1 _09405_/X sky130_fd_sc_hd__and3_1
XFILLER_81_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_996 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_164 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07597_ _07594_/Y _07599_/B _07607_/A vssd1 vssd1 vccd1 vccd1 _07597_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_164_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09336_ _13144_/A0 _09334_/X _09335_/X vssd1 vssd1 vccd1 vccd1 _09340_/B sky130_fd_sc_hd__a21o_1
XFILLER_179_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09267_ _14472_/Q _09558_/A2 _09266_/X _13049_/A1 vssd1 vssd1 vccd1 vccd1 _09267_/X
+ sky130_fd_sc_hd__a211o_1
Xclkbuf_leaf_141_clk clkbuf_5_28_0_clk/X vssd1 vssd1 vccd1 vccd1 _15548_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_138_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08218_ _13709_/Q _11847_/A1 _08221_/S vssd1 vssd1 vccd1 vccd1 _13709_/D sky130_fd_sc_hd__mux2_1
XFILLER_166_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09198_ _13921_/Q _09197_/X _12481_/A vssd1 vssd1 vccd1 vccd1 _13921_/D sky130_fd_sc_hd__mux2_1
XFILLER_14_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08149_ _08150_/S input25/X vssd1 vssd1 vccd1 vccd1 _08185_/B sky130_fd_sc_hd__and2b_1
XFILLER_162_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11160_ _11129_/A _11113_/X _11129_/Y vssd1 vssd1 vccd1 vccd1 _11199_/B sky130_fd_sc_hd__a21oi_2
XFILLER_136_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10111_ _14497_/Q _14745_/Q _10131_/S vssd1 vssd1 vccd1 vccd1 _14497_/D sky130_fd_sc_hd__mux2_1
XFILLER_161_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11091_ _11380_/A _11177_/B _10984_/Y vssd1 vssd1 vccd1 vccd1 _11091_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10042_ _14399_/Q _13328_/A0 _10059_/S vssd1 vssd1 vccd1 vccd1 _14399_/D sky130_fd_sc_hd__mux2_1
XFILLER_1_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14850_ _15500_/CLK _14850_/D vssd1 vssd1 vccd1 vccd1 _14850_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_76_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_64 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13801_ _15646_/CLK _13801_/D vssd1 vssd1 vccd1 vccd1 _13801_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_35_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14781_ _15599_/CLK _14781_/D vssd1 vssd1 vccd1 vccd1 _14781_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11993_ _14071_/Q _14039_/Q _11993_/S vssd1 vssd1 vccd1 vccd1 _11993_/X sky130_fd_sc_hd__mux2_1
XFILLER_91_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13732_ _15530_/CLK _13732_/D vssd1 vssd1 vccd1 vccd1 _13732_/Q sky130_fd_sc_hd__dfxtp_2
X_10944_ wire360/X _10944_/B vssd1 vssd1 vccd1 vccd1 _10944_/Y sky130_fd_sc_hd__nand2_1
XFILLER_91_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13663_ _14774_/CLK _13663_/D vssd1 vssd1 vccd1 vccd1 _13663_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10875_ _13731_/Q _14907_/Q _13129_/A vssd1 vssd1 vccd1 vccd1 _14907_/D sky130_fd_sc_hd__mux2_1
XFILLER_31_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15402_ _15587_/CLK _15402_/D vssd1 vssd1 vccd1 vccd1 _15402_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_176_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12614_ _14098_/Q _14066_/Q _12614_/S vssd1 vssd1 vccd1 vccd1 _12614_/X sky130_fd_sc_hd__mux2_1
XFILLER_188_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13594_ _15630_/CLK _13594_/D vssd1 vssd1 vccd1 vccd1 _13594_/Q sky130_fd_sc_hd__dfxtp_2
XPHY_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15333_ _15670_/CLK _15333_/D vssd1 vssd1 vccd1 vccd1 _15333_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_157_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12545_ _14095_/Q _14063_/Q _12545_/S vssd1 vssd1 vccd1 vccd1 _12545_/X sky130_fd_sc_hd__mux2_1
XFILLER_129_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_132_clk clkbuf_5_28_0_clk/X vssd1 vssd1 vccd1 vccd1 _15397_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_129_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15264_ _15336_/CLK _15264_/D vssd1 vssd1 vccd1 vccd1 _15264_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12476_ _14092_/Q _14060_/Q _12476_/S vssd1 vssd1 vccd1 vccd1 _12476_/X sky130_fd_sc_hd__mux2_1
XFILLER_138_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14215_ _15275_/CLK _14215_/D vssd1 vssd1 vccd1 vccd1 _14215_/Q sky130_fd_sc_hd__dfxtp_1
X_11427_ _11437_/A _11436_/A _11437_/B _13229_/A vssd1 vssd1 vccd1 vccd1 _11428_/B
+ sky130_fd_sc_hd__a31o_1
XANTENNA_5 _08744_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15195_ _15336_/CLK _15195_/D vssd1 vssd1 vccd1 vccd1 _15195_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_126_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14146_ _15664_/CLK _14146_/D vssd1 vssd1 vccd1 vccd1 _14146_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_152_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11358_ _11357_/B _11357_/C _13159_/B vssd1 vssd1 vccd1 vccd1 _11359_/B sky130_fd_sc_hd__a21oi_1
XFILLER_180_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10309_ _14694_/Q _14879_/Q _10665_/S vssd1 vssd1 vccd1 vccd1 _14694_/D sky130_fd_sc_hd__mux2_1
X_14077_ _15133_/CLK _14077_/D vssd1 vssd1 vccd1 vccd1 _14077_/Q sky130_fd_sc_hd__dfxtp_1
X_11289_ _11259_/X _11288_/X _11297_/S vssd1 vssd1 vccd1 vccd1 _11289_/X sky130_fd_sc_hd__mux2_1
XFILLER_3_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13028_ _15489_/Q _10892_/B _13116_/C _13027_/X vssd1 vssd1 vccd1 vccd1 _15489_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_100_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_199_clk clkbuf_5_17_0_clk/X vssd1 vssd1 vccd1 vccd1 _15211_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_39_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14979_ _14988_/CLK _14979_/D vssd1 vssd1 vccd1 vccd1 _14979_/Q sky130_fd_sc_hd__dfxtp_1
X_07520_ _14750_/Q _13429_/Q _07529_/S vssd1 vssd1 vccd1 vccd1 _13429_/D sky130_fd_sc_hd__mux2_1
XFILLER_81_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07451_ _13668_/Q _07483_/A2 _07483_/B1 _14696_/Q _07450_/X vssd1 vssd1 vccd1 vccd1
+ _07451_/X sky130_fd_sc_hd__a221o_1
XFILLER_34_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_179_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07382_ _14647_/Q _07498_/B _07498_/C vssd1 vssd1 vccd1 vccd1 _07382_/X sky130_fd_sc_hd__and3_1
XFILLER_176_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_1081 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09121_ _14465_/Q _14433_/Q _13854_/Q _14207_/Q _09190_/S _09429_/S1 vssd1 vssd1
+ vccd1 vccd1 _09121_/X sky130_fd_sc_hd__mux4_1
XFILLER_31_882 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_123_clk clkbuf_5_31_0_clk/X vssd1 vssd1 vccd1 vccd1 _15385_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_148_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09052_ _09419_/A2 _09050_/X _09051_/X _09421_/A1 vssd1 vssd1 vccd1 vccd1 _09052_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_136_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08003_ _13567_/Q _08003_/B vssd1 vssd1 vccd1 vccd1 _08003_/X sky130_fd_sc_hd__xor2_1
XFILLER_163_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09954_ _11874_/A1 _14314_/Q _09963_/S vssd1 vssd1 vccd1 vccd1 _14314_/D sky130_fd_sc_hd__mux2_1
X_08905_ _14357_/Q _15173_/Q _13812_/Q _14551_/Q _09469_/S _09546_/S1 vssd1 vssd1
+ vccd1 vccd1 _08906_/B sky130_fd_sc_hd__mux4_1
XFILLER_103_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09885_ _13338_/A0 _14247_/Q _09897_/S vssd1 vssd1 vccd1 vccd1 _14247_/D sky130_fd_sc_hd__mux2_1
XFILLER_140_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08836_ _13859_/Q _11868_/A1 _08846_/S vssd1 vssd1 vccd1 vccd1 _13859_/D sky130_fd_sc_hd__mux2_1
XFILLER_58_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08767_ _13125_/B _08769_/B vssd1 vssd1 vccd1 vccd1 _08767_/Y sky130_fd_sc_hd__nor2_1
XTAP_2705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07718_ _07715_/Y _07724_/C _07713_/A vssd1 vssd1 vccd1 vccd1 _07718_/Y sky130_fd_sc_hd__o21ai_1
XTAP_2738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08698_ _13452_/Q _08746_/A2 _08750_/A2 _13516_/Q _08696_/X vssd1 vssd1 vccd1 vccd1
+ _08698_/X sky130_fd_sc_hd__a221o_1
XFILLER_82_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07649_ _14763_/Q _07644_/A _07648_/Y _08016_/C1 vssd1 vssd1 vccd1 vccd1 _13474_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_53_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10660_ _14750_/Q _10659_/X _10710_/S vssd1 vssd1 vccd1 vccd1 _14750_/D sky130_fd_sc_hd__mux2_1
XFILLER_40_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09319_ _15096_/Q _08519_/B _09519_/B1 _08501_/A vssd1 vssd1 vccd1 vccd1 _09319_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_22_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_114_clk _15447_/CLK vssd1 vssd1 vccd1 vccd1 _15379_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_166_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10591_ _14997_/Q _10569_/B _10733_/B1 _14933_/Q _10732_/C1 vssd1 vssd1 vccd1 vccd1
+ _10591_/X sky130_fd_sc_hd__a221o_1
X_12330_ _12615_/B1 _12327_/X _12616_/C1 vssd1 vssd1 vccd1 vccd1 _12330_/X sky130_fd_sc_hd__o21a_1
XFILLER_182_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12261_ _12500_/B1 _12258_/X _12501_/C1 vssd1 vssd1 vccd1 vccd1 _12261_/X sky130_fd_sc_hd__o21a_1
XFILLER_5_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14000_ _15130_/CLK _14000_/D vssd1 vssd1 vccd1 vccd1 _14000_/Q sky130_fd_sc_hd__dfxtp_1
X_11212_ _10399_/A _15001_/Q _11237_/S vssd1 vssd1 vccd1 vccd1 _15001_/D sky130_fd_sc_hd__mux2_1
XFILLER_134_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12192_ _12500_/B1 _12189_/X _12501_/C1 vssd1 vssd1 vccd1 vccd1 _12192_/X sky130_fd_sc_hd__o21a_1
XFILLER_150_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput42 _07178_/X vssd1 vssd1 vccd1 vccd1 ext_address[16] sky130_fd_sc_hd__clkbuf_2
Xoutput53 _07189_/X vssd1 vssd1 vccd1 vccd1 ext_address[27] sky130_fd_sc_hd__clkbuf_2
X_11143_ _08233_/B _11142_/X _10984_/Y vssd1 vssd1 vccd1 vccd1 _11143_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_150_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput64 _07170_/X vssd1 vssd1 vccd1 vccd1 ext_address[8] sky130_fd_sc_hd__clkbuf_2
XFILLER_96_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput75 _07135_/X vssd1 vssd1 vccd1 vccd1 ext_write_data[17] sky130_fd_sc_hd__clkbuf_2
Xoutput86 _07155_/X vssd1 vssd1 vccd1 vccd1 ext_write_data[27] sky130_fd_sc_hd__clkbuf_2
XFILLER_49_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput97 _07117_/X vssd1 vssd1 vccd1 vccd1 ext_write_data[8] sky130_fd_sc_hd__clkbuf_2
XFILLER_95_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11074_ _11017_/X _11027_/X _11330_/A vssd1 vssd1 vccd1 vccd1 _11074_/X sky130_fd_sc_hd__mux2_1
X_14902_ _15540_/CLK _14902_/D vssd1 vssd1 vccd1 vccd1 _14902_/Q sky130_fd_sc_hd__dfxtp_1
X_10025_ _11879_/A1 _14383_/Q _10029_/S vssd1 vssd1 vccd1 vccd1 _14383_/D sky130_fd_sc_hd__mux2_1
XFILLER_48_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14833_ _15497_/CLK _14833_/D vssd1 vssd1 vccd1 vccd1 _14833_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_48_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14764_ _14892_/CLK _14764_/D vssd1 vssd1 vccd1 vccd1 _14764_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_3984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11976_ _15309_/Q _13081_/A2 _11975_/X vssd1 vssd1 vccd1 vccd1 _15309_/D sky130_fd_sc_hd__a21o_1
XFILLER_60_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13715_ _14468_/CLK _13715_/D vssd1 vssd1 vccd1 vccd1 _13715_/Q sky130_fd_sc_hd__dfxtp_1
X_10927_ _11536_/A _10929_/B vssd1 vssd1 vccd1 vccd1 _10927_/Y sky130_fd_sc_hd__nand2_1
XFILLER_60_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14695_ _15452_/CLK _14695_/D vssd1 vssd1 vccd1 vccd1 _14695_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13646_ _15372_/CLK _13646_/D vssd1 vssd1 vccd1 vccd1 _13646_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_158_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10858_ _14890_/Q _13778_/Q _12933_/S vssd1 vssd1 vccd1 vccd1 _14890_/D sky130_fd_sc_hd__mux2_1
XFILLER_13_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_176_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_105_clk clkbuf_5_26_0_clk/X vssd1 vssd1 vccd1 vccd1 _15641_/CLK sky130_fd_sc_hd__clkbuf_16
X_13577_ _15372_/CLK _13577_/D vssd1 vssd1 vccd1 vccd1 _13577_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_169_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10789_ _14821_/Q _15453_/Q _12929_/S vssd1 vssd1 vccd1 vccd1 _14821_/D sky130_fd_sc_hd__mux2_1
XPHY_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15316_ _15664_/CLK _15316_/D vssd1 vssd1 vccd1 vccd1 _15316_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_185_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12528_ _15333_/Q _13154_/S _12527_/X vssd1 vssd1 vccd1 vccd1 _15333_/D sky130_fd_sc_hd__a21o_1
XFILLER_9_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15247_ _15279_/CLK _15247_/D vssd1 vssd1 vccd1 vccd1 _15247_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12459_ _15330_/Q _13119_/S _12458_/X vssd1 vssd1 vccd1 vccd1 _15330_/D sky130_fd_sc_hd__a21o_1
X_15178_ _15178_/CLK _15178_/D vssd1 vssd1 vccd1 vccd1 _15178_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_153_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14129_ _15672_/CLK _14129_/D vssd1 vssd1 vccd1 vccd1 _14129_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout309 _07452_/X vssd1 vssd1 vccd1 vccd1 _13338_/A0 sky130_fd_sc_hd__buf_6
XFILLER_67_1088 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06951_ _14488_/Q _06751_/Y _14487_/Q _06754_/Y _06960_/A vssd1 vssd1 vccd1 vccd1
+ _06951_/X sky130_fd_sc_hd__a221o_1
XFILLER_39_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09670_ _14041_/Q _13325_/A0 _09690_/S vssd1 vssd1 vccd1 vccd1 _14041_/D sky130_fd_sc_hd__mux2_1
X_06882_ _06882_/A _06882_/B _06882_/C _06882_/D vssd1 vssd1 vccd1 vccd1 _06882_/Y
+ sky130_fd_sc_hd__nor4_1
XFILLER_55_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08621_ _13527_/Q _08683_/A2 _08693_/B1 _13630_/Q vssd1 vssd1 vccd1 vccd1 _08621_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_94_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08552_ _08722_/A _08552_/B _08552_/C vssd1 vssd1 vccd1 vccd1 _08552_/X sky130_fd_sc_hd__or3_1
XFILLER_130_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07503_ _14720_/Q _14719_/Q vssd1 vssd1 vccd1 vccd1 _08037_/C sky130_fd_sc_hd__nand2b_2
XFILLER_35_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08483_ _13771_/Q _08482_/X _12906_/S vssd1 vssd1 vccd1 vccd1 _13771_/D sky130_fd_sc_hd__mux2_1
XFILLER_74_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07434_ _14660_/Q _07474_/B _07482_/C vssd1 vssd1 vccd1 vccd1 _07434_/X sky130_fd_sc_hd__and3_1
XFILLER_161_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07365_ _07365_/A _07365_/B vssd1 vssd1 vccd1 vccd1 _14925_/D sky130_fd_sc_hd__xnor2_1
XFILLER_148_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09104_ _09449_/A1 _09102_/X _09103_/X _09449_/B2 _09101_/X vssd1 vssd1 vccd1 vccd1
+ _09104_/X sky130_fd_sc_hd__a221o_2
XFILLER_182_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07296_ _13918_/Q _15505_/Q _07339_/S vssd1 vssd1 vccd1 vccd1 _07297_/A sky130_fd_sc_hd__mux2_8
XFILLER_148_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09035_ _09033_/X _09034_/X _12596_/A _09024_/X vssd1 vssd1 vccd1 vccd1 _09035_/X
+ sky130_fd_sc_hd__o211a_2
XFILLER_184_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09937_ _11857_/A1 _14297_/Q _09963_/S vssd1 vssd1 vccd1 vccd1 _14297_/D sky130_fd_sc_hd__mux2_1
XFILLER_58_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09868_ _13321_/A0 _14230_/Q _09897_/S vssd1 vssd1 vccd1 vccd1 _14230_/D sky130_fd_sc_hd__mux2_1
XTAP_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08819_ _13318_/D _10065_/A vssd1 vssd1 vccd1 vccd1 _08819_/Y sky130_fd_sc_hd__nor2_8
XTAP_3225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09799_ _14165_/Q _13321_/A0 _09828_/S vssd1 vssd1 vccd1 vccd1 _14165_/D sky130_fd_sc_hd__mux2_1
XTAP_3247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11830_ _15252_/Q _13330_/A0 _11849_/S vssd1 vssd1 vccd1 vccd1 _15252_/D sky130_fd_sc_hd__mux2_1
XTAP_2524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11761_ _11761_/A0 _15189_/Q _11775_/S vssd1 vssd1 vccd1 vccd1 _15189_/D sky130_fd_sc_hd__mux2_1
XTAP_1834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13500_ _13565_/CLK _13500_/D vssd1 vssd1 vccd1 vccd1 _13500_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10712_ _15580_/Q _10706_/B _10733_/B1 _14957_/Q vssd1 vssd1 vccd1 vccd1 _10712_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_1867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14480_ _15558_/CLK _14480_/D vssd1 vssd1 vccd1 vccd1 _14480_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11692_ _13082_/B2 _15123_/Q _11703_/S vssd1 vssd1 vccd1 vccd1 _15123_/D sky130_fd_sc_hd__mux2_1
XFILLER_42_999 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13431_ _15383_/CLK _13431_/D vssd1 vssd1 vccd1 vccd1 _13431_/Q sky130_fd_sc_hd__dfxtp_2
X_10643_ _14975_/Q _10718_/A2 _10722_/B1 _14943_/Q _10642_/X vssd1 vssd1 vccd1 vccd1
+ _10643_/X sky130_fd_sc_hd__a221o_1
XFILLER_9_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_52 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13362_ _14465_/Q vssd1 vssd1 vccd1 vccd1 _14465_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_42_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10574_ _14929_/Q _14994_/Q _10569_/B _10731_/B _15553_/Q vssd1 vssd1 vccd1 vccd1
+ _10574_/X sky130_fd_sc_hd__a32o_1
X_15101_ _15133_/CLK _15101_/D vssd1 vssd1 vccd1 vccd1 _15101_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_158_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12313_ _14021_/Q _13989_/Q _12614_/S vssd1 vssd1 vccd1 vccd1 _12314_/B sky130_fd_sc_hd__mux2_1
XFILLER_166_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13293_ _12673_/X _15625_/Q _13300_/S vssd1 vssd1 vccd1 vccd1 _15625_/D sky130_fd_sc_hd__mux2_1
XFILLER_182_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15032_ _15042_/CLK _15032_/D vssd1 vssd1 vccd1 vccd1 _15032_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_182_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12244_ _14018_/Q _13986_/Q _12246_/S vssd1 vssd1 vccd1 vccd1 _12245_/B sky130_fd_sc_hd__mux2_1
XFILLER_182_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12175_ _14015_/Q _13983_/Q _12246_/S vssd1 vssd1 vccd1 vccd1 _12176_/B sky130_fd_sc_hd__mux2_1
XFILLER_122_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11126_ _11371_/A _11124_/X _11125_/X vssd1 vssd1 vccd1 vccd1 _11126_/X sky130_fd_sc_hd__a21o_1
XFILLER_110_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_275 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11057_ _11053_/X _11056_/X _11252_/A vssd1 vssd1 vccd1 vccd1 _11058_/A sky130_fd_sc_hd__mux2_2
XFILLER_49_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_82 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_716 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10008_ _13072_/B2 _14366_/Q _10028_/S vssd1 vssd1 vccd1 vccd1 _14366_/D sky130_fd_sc_hd__mux2_1
XFILLER_76_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_598 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14816_ _15634_/CLK _14816_/D vssd1 vssd1 vccd1 vccd1 _14816_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_184_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14747_ _15569_/CLK _14747_/D vssd1 vssd1 vccd1 vccd1 _14747_/Q sky130_fd_sc_hd__dfxtp_4
X_11959_ _14359_/Q _15175_/Q _13814_/Q _14553_/Q _12269_/S _12268_/A vssd1 vssd1 vccd1
+ vccd1 _11959_/X sky130_fd_sc_hd__mux4_1
XFILLER_44_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14678_ _15616_/CLK _14678_/D vssd1 vssd1 vccd1 vccd1 _14678_/Q sky130_fd_sc_hd__dfxtp_1
X_13629_ _15386_/CLK _13629_/D vssd1 vssd1 vccd1 vccd1 _13629_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07150_ _14855_/Q _14847_/Q _14839_/Q _14831_/Q _07146_/S _07104_/C vssd1 vssd1 vccd1
+ vccd1 _07151_/B sky130_fd_sc_hd__mux4_1
XFILLER_146_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07081_ _14639_/Q _14671_/Q _07096_/S vssd1 vssd1 vccd1 vccd1 _07081_/X sky130_fd_sc_hd__mux2_1
XFILLER_161_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout106 _12621_/Y vssd1 vssd1 vccd1 vccd1 _12737_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_141_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout117 _12944_/Y vssd1 vssd1 vccd1 vccd1 _13024_/A2 sky130_fd_sc_hd__clkbuf_16
XFILLER_141_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout128 _10759_/S vssd1 vssd1 vccd1 vccd1 _10764_/S sky130_fd_sc_hd__buf_12
X_07983_ _14754_/Q _07971_/A _07982_/Y vssd1 vssd1 vccd1 vccd1 _13561_/D sky130_fd_sc_hd__o21a_1
Xfanout139 _12320_/A vssd1 vssd1 vccd1 vccd1 _12481_/A sky130_fd_sc_hd__buf_12
XFILLER_86_126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09722_ _13344_/A0 _14092_/Q _09723_/S vssd1 vssd1 vccd1 vccd1 _14092_/D sky130_fd_sc_hd__mux2_1
X_06934_ _06730_/Y _13488_/Q _14496_/Q _06732_/Y vssd1 vssd1 vccd1 vccd1 _06934_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_55_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09653_ _14026_/Q _13342_/A0 _09661_/S vssd1 vssd1 vccd1 vccd1 _14026_/D sky130_fd_sc_hd__mux2_1
X_06865_ input33/X _06865_/B _13316_/S _06997_/B vssd1 vssd1 vccd1 vccd1 _15615_/D
+ sky130_fd_sc_hd__and4_2
XFILLER_28_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08604_ _14507_/Q _08748_/B1 _08602_/X _08603_/X vssd1 vssd1 vccd1 vccd1 _08605_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_43_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09584_ _13960_/Q _11873_/A1 _09594_/S vssd1 vssd1 vccd1 vccd1 _13960_/D sky130_fd_sc_hd__mux2_1
X_06796_ _14597_/Q _06796_/B vssd1 vssd1 vccd1 vccd1 _06797_/A sky130_fd_sc_hd__nor2_1
XFILLER_24_900 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08535_ _08910_/S _08668_/B _08724_/C _08668_/D vssd1 vssd1 vccd1 vccd1 _08535_/X
+ sky130_fd_sc_hd__and4_2
XFILLER_35_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08466_ _08421_/Y _08465_/X _14614_/Q vssd1 vssd1 vccd1 vccd1 _08466_/X sky130_fd_sc_hd__o21a_1
XFILLER_50_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07417_ _13329_/A0 _13393_/Q _07481_/S vssd1 vssd1 vccd1 vccd1 _13393_/D sky130_fd_sc_hd__mux2_1
XFILLER_149_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08397_ _13731_/Q _13140_/S _08394_/X _14592_/Q vssd1 vssd1 vccd1 vccd1 _13731_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_149_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_150 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07348_ _07348_/A _07348_/B _07287_/X vssd1 vssd1 vccd1 vccd1 _07351_/C sky130_fd_sc_hd__or3b_1
XFILLER_164_621 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07279_ _13921_/Q _15508_/Q _07339_/S vssd1 vssd1 vccd1 vccd1 _07280_/A sky130_fd_sc_hd__mux2_8
XFILLER_164_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09018_ _15279_/Q _15247_/Q _15215_/Q _15146_/Q _09073_/S _09234_/S1 vssd1 vssd1
+ vccd1 vccd1 _09018_/X sky130_fd_sc_hd__mux4_1
XFILLER_88_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_570 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10290_ _14675_/Q _14828_/Q _10610_/S vssd1 vssd1 vccd1 vccd1 _14675_/D sky130_fd_sc_hd__mux2_1
XFILLER_151_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_859 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout640 fanout647/X vssd1 vssd1 vccd1 vccd1 _07938_/C1 sky130_fd_sc_hd__buf_4
XFILLER_59_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13980_ _14415_/CLK _13980_/D vssd1 vssd1 vccd1 vccd1 _13980_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_120_768 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12931_ _15459_/Q _15645_/Q _12933_/S vssd1 vssd1 vccd1 vccd1 _15459_/D sky130_fd_sc_hd__mux2_1
XFILLER_46_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12862_ _14756_/Q _15390_/Q _12866_/S vssd1 vssd1 vccd1 vccd1 _15390_/D sky130_fd_sc_hd__mux2_1
X_15650_ _15650_/CLK _15650_/D vssd1 vssd1 vccd1 vccd1 _15650_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_74_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14601_ _15536_/CLK _14601_/D vssd1 vssd1 vccd1 vccd1 _14601_/Q sky130_fd_sc_hd__dfxtp_4
X_11813_ _15236_/Q _11879_/A1 _11817_/S vssd1 vssd1 vccd1 vccd1 _15236_/D sky130_fd_sc_hd__mux2_1
XTAP_3099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15581_ _15581_/CLK _15581_/D vssd1 vssd1 vccd1 vccd1 _15581_/Q sky130_fd_sc_hd__dfxtp_1
X_12793_ _13438_/Q _12647_/B _08030_/Y _13605_/Q _12743_/A vssd1 vssd1 vccd1 vccd1
+ _12793_/X sky130_fd_sc_hd__a221o_2
XTAP_1620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14532_ _15674_/CLK _14532_/D vssd1 vssd1 vccd1 vccd1 _14532_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11744_ _11852_/A1 _15172_/Q _11774_/S vssd1 vssd1 vccd1 vccd1 _15172_/D sky130_fd_sc_hd__mux2_1
XFILLER_57_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1076 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14463_ _15663_/CLK _14463_/D vssd1 vssd1 vccd1 vccd1 _14463_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_186_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11675_ _13350_/A0 _15107_/Q _11675_/S vssd1 vssd1 vccd1 vccd1 _15107_/D sky130_fd_sc_hd__mux2_1
XFILLER_169_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13414_ _15326_/CLK _13414_/D vssd1 vssd1 vccd1 vccd1 _13414_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10626_ _15563_/Q _10706_/B vssd1 vssd1 vccd1 vccd1 _10626_/X sky130_fd_sc_hd__and2_1
XFILLER_186_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14394_ _15108_/CLK _14394_/D vssd1 vssd1 vccd1 vccd1 _14394_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13345_ _13345_/A0 _15675_/Q _13345_/S vssd1 vssd1 vccd1 vccd1 _15675_/D sky130_fd_sc_hd__mux2_1
XFILLER_127_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10557_ _10557_/A _10557_/B _10557_/C vssd1 vssd1 vccd1 vccd1 _10558_/C sky130_fd_sc_hd__or3_1
XFILLER_6_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13276_ _15360_/Q _15607_/Q _13300_/S vssd1 vssd1 vccd1 vccd1 _15607_/D sky130_fd_sc_hd__mux2_1
XFILLER_142_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10488_ _07238_/X _10523_/A2 _10487_/X vssd1 vssd1 vccd1 vccd1 _11563_/A sky130_fd_sc_hd__a21o_4
XFILLER_29_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15015_ _15017_/CLK _15015_/D vssd1 vssd1 vccd1 vccd1 _15015_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_142_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12227_ _12273_/A1 _12226_/X _12225_/X _12503_/C1 vssd1 vssd1 vccd1 vccd1 _12228_/C
+ sky130_fd_sc_hd__a211o_2
XFILLER_64_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12158_ _12273_/A1 _12157_/X _12156_/X _12503_/C1 vssd1 vssd1 vccd1 vccd1 _12159_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_25_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_1039 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11109_ _11298_/A _11107_/X _11108_/X vssd1 vssd1 vccd1 vccd1 _11109_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_1_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12089_ _12273_/A1 _12088_/X _12087_/X _12503_/C1 vssd1 vssd1 vccd1 vccd1 _12090_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_37_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08320_ _11283_/A _11252_/A vssd1 vssd1 vccd1 vccd1 _08320_/Y sky130_fd_sc_hd__nor2_2
XFILLER_36_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_763 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08251_ _11129_/A _11115_/S _11259_/S _11023_/A vssd1 vssd1 vccd1 vccd1 _11437_/A
+ sky130_fd_sc_hd__and4_4
XFILLER_178_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07202_ _13935_/Q _15522_/Q _07334_/S vssd1 vssd1 vccd1 vccd1 _07202_/X sky130_fd_sc_hd__mux2_8
XFILLER_177_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08182_ _13678_/Q _10730_/S _08155_/X _08181_/X vssd1 vssd1 vccd1 vccd1 _13678_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_9_480 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07133_ _14830_/Q _07104_/X _07132_/X _07131_/A vssd1 vssd1 vccd1 vccd1 _07133_/X
+ sky130_fd_sc_hd__a22o_4
X_07064_ _07063_/X _13600_/Q _12764_/S vssd1 vssd1 vccd1 vccd1 _07064_/X sky130_fd_sc_hd__mux2_1
XFILLER_145_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07966_ _13557_/Q _07973_/D vssd1 vssd1 vccd1 vccd1 _07970_/B sky130_fd_sc_hd__nand2_1
X_09705_ _13327_/A0 _14075_/Q _09723_/S vssd1 vssd1 vccd1 vccd1 _14075_/D sky130_fd_sc_hd__mux2_1
XFILLER_56_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06917_ _15389_/Q _06711_/Y _06712_/Y _13465_/Q vssd1 vssd1 vccd1 vccd1 _06921_/B
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_114_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07897_ _13539_/Q _07897_/B vssd1 vssd1 vccd1 vccd1 _07898_/B sky130_fd_sc_hd__xor2_1
XFILLER_28_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_94_clk clkbuf_5_24_0_clk/X vssd1 vssd1 vccd1 vccd1 _15646_/CLK sky130_fd_sc_hd__clkbuf_16
X_09636_ _14009_/Q _13325_/A0 _09661_/S vssd1 vssd1 vccd1 vccd1 _14009_/D sky130_fd_sc_hd__mux2_1
XFILLER_71_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06848_ _14905_/Q _14908_/Q _14907_/Q _14909_/Q vssd1 vssd1 vccd1 vccd1 _06848_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_43_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09567_ _13943_/Q _11681_/A0 _09589_/S vssd1 vssd1 vccd1 vccd1 _13943_/D sky130_fd_sc_hd__mux2_1
X_06779_ _07096_/S _14730_/Q vssd1 vssd1 vccd1 vccd1 _10244_/S sky130_fd_sc_hd__nand2_8
XFILLER_70_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08518_ _13125_/A _08521_/A vssd1 vssd1 vccd1 vccd1 _08518_/Y sky130_fd_sc_hd__nor2_8
X_09498_ _06675_/Y _09497_/X _09496_/X _09524_/A vssd1 vssd1 vccd1 vccd1 _09498_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_90_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08449_ _08449_/A _08773_/B vssd1 vssd1 vccd1 vccd1 _08449_/X sky130_fd_sc_hd__and2_1
XFILLER_23_32 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11460_ _11425_/B _11460_/B _11460_/C _11460_/D vssd1 vssd1 vccd1 vccd1 _11464_/B
+ sky130_fd_sc_hd__and4b_2
XFILLER_165_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10411_ _10410_/A _10408_/Y _10556_/A vssd1 vssd1 vccd1 vccd1 _10411_/X sky130_fd_sc_hd__a21o_1
XFILLER_87_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11391_ _11390_/B _11390_/C _13171_/B vssd1 vssd1 vccd1 vccd1 _11401_/C sky130_fd_sc_hd__a21o_1
XFILLER_104_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13130_ _13123_/B _08507_/Y _13130_/B1 _13130_/C1 vssd1 vssd1 vccd1 vccd1 _13130_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_139_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10342_ _14727_/Q _14920_/Q _10343_/S vssd1 vssd1 vccd1 vccd1 _14727_/D sky130_fd_sc_hd__mux2_1
XFILLER_174_1006 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13061_ _15498_/Q _13081_/A2 _13105_/B1 _13060_/X vssd1 vssd1 vccd1 vccd1 _15498_/D
+ sky130_fd_sc_hd__a22o_1
X_10273_ _14658_/Q _14811_/Q _10650_/S vssd1 vssd1 vccd1 vccd1 _14658_/D sky130_fd_sc_hd__mux2_1
XFILLER_79_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12012_ _13880_/Q _14395_/Q _12407_/S vssd1 vssd1 vccd1 vccd1 _12012_/X sky130_fd_sc_hd__mux2_1
XFILLER_2_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1020 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout470 _12618_/A1 vssd1 vssd1 vccd1 vccd1 _12595_/A1 sky130_fd_sc_hd__buf_12
Xfanout481 _06670_/Y vssd1 vssd1 vccd1 vccd1 _12548_/S sky130_fd_sc_hd__buf_12
XFILLER_24_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_991 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout492 _15044_/Q vssd1 vssd1 vccd1 vccd1 _07104_/C sky130_fd_sc_hd__buf_12
XFILLER_150_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13963_ _15673_/CLK _13963_/D vssd1 vssd1 vccd1 vccd1 _13963_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_85_clk clkbuf_5_12_0_clk/X vssd1 vssd1 vccd1 vccd1 _14868_/CLK sky130_fd_sc_hd__clkbuf_16
X_12914_ _15442_/Q _15628_/Q _12917_/S vssd1 vssd1 vccd1 vccd1 _15442_/D sky130_fd_sc_hd__mux2_1
XFILLER_47_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13894_ _15127_/CLK _13894_/D vssd1 vssd1 vccd1 vccd1 _13894_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_46_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15633_ _15634_/CLK _15633_/D vssd1 vssd1 vccd1 vccd1 _15633_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12845_ _14739_/Q _15373_/Q _12871_/S vssd1 vssd1 vccd1 vccd1 _15373_/D sky130_fd_sc_hd__mux2_1
XTAP_2151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15564_ _15580_/CLK _15564_/D vssd1 vssd1 vccd1 vccd1 _15564_/Q sky130_fd_sc_hd__dfxtp_1
X_12776_ _15359_/Q _12776_/B vssd1 vssd1 vccd1 vccd1 _12777_/B sky130_fd_sc_hd__or2_1
XTAP_1450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11727_ _15156_/Q _11868_/A1 _11741_/S vssd1 vssd1 vccd1 vccd1 _15156_/D sky130_fd_sc_hd__mux2_1
X_14515_ _15398_/CLK _14515_/D vssd1 vssd1 vccd1 vccd1 _14515_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15495_ _15499_/CLK _15495_/D vssd1 vssd1 vccd1 vccd1 _15495_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_175_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11658_ _13333_/A0 _15090_/Q _11670_/S vssd1 vssd1 vccd1 vccd1 _15090_/D sky130_fd_sc_hd__mux2_1
X_14446_ _15518_/CLK _14446_/D vssd1 vssd1 vccd1 vccd1 _14446_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_1062 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10609_ _15049_/Q _10734_/A2 _10606_/X _10608_/X vssd1 vssd1 vccd1 vccd1 _10609_/X
+ sky130_fd_sc_hd__o22a_2
XFILLER_128_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14377_ _14485_/CLK _14377_/D vssd1 vssd1 vccd1 vccd1 _14377_/Q sky130_fd_sc_hd__dfxtp_1
X_11589_ _11582_/A _11589_/B _11589_/C vssd1 vssd1 vccd1 vccd1 _11598_/B sky130_fd_sc_hd__nand3b_1
X_13328_ _13328_/A0 _15658_/Q _13345_/S vssd1 vssd1 vccd1 vccd1 _15658_/D sky130_fd_sc_hd__mux2_1
XFILLER_155_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13259_ _15343_/Q _15590_/Q _13291_/S vssd1 vssd1 vccd1 vccd1 _15590_/D sky130_fd_sc_hd__mux2_1
XFILLER_43_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07820_ _14743_/Q _07830_/A _07819_/Y _12809_/C1 vssd1 vssd1 vccd1 vccd1 _13518_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_38_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07751_ _14758_/Q _07750_/A _07750_/Y _08002_/C1 vssd1 vssd1 vccd1 vccd1 _13501_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_38_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_76_clk clkbuf_5_15_0_clk/X vssd1 vssd1 vccd1 vccd1 _15632_/CLK sky130_fd_sc_hd__clkbuf_16
X_06702_ _15393_/Q vssd1 vssd1 vccd1 vccd1 _06702_/Y sky130_fd_sc_hd__inv_2
XFILLER_38_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07682_ _13483_/Q _07687_/C vssd1 vssd1 vccd1 vccd1 _07682_/Y sky130_fd_sc_hd__nor2_1
XFILLER_25_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09421_ _09421_/A1 _09417_/X _09420_/X _09416_/X vssd1 vssd1 vccd1 vccd1 _09421_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_52_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09352_ _14250_/Q _14282_/Q _14314_/Q _14346_/Q _09521_/S _09523_/A1 vssd1 vssd1
+ vccd1 vccd1 _09352_/X sky130_fd_sc_hd__mux4_1
XFILLER_178_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08303_ _07317_/A _10481_/B _08302_/X vssd1 vssd1 vccd1 vccd1 _13178_/B sky130_fd_sc_hd__a21oi_4
XFILLER_127_1041 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09283_ _14375_/Q _15191_/Q _13830_/Q _14569_/Q _09484_/S _08519_/A vssd1 vssd1 vccd1
+ vccd1 _09284_/B sky130_fd_sc_hd__mux4_1
XFILLER_138_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08234_ _08240_/A _13804_/Q _13772_/Q _08237_/A vssd1 vssd1 vccd1 vccd1 _08234_/X
+ sky130_fd_sc_hd__a22o_4
XFILLER_178_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08165_ _08185_/A _08165_/B vssd1 vssd1 vccd1 vccd1 _08165_/X sky130_fd_sc_hd__and2_1
XFILLER_109_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07116_ _14838_/Q _14830_/Q _07146_/S vssd1 vssd1 vccd1 vccd1 _07117_/B sky130_fd_sc_hd__mux2_1
XFILLER_180_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08096_ _10730_/S _08121_/B vssd1 vssd1 vccd1 vccd1 _08096_/X sky130_fd_sc_hd__and2_4
XFILLER_173_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07047_ _07046_/X _14748_/Q _07077_/S vssd1 vssd1 vccd1 vccd1 _13594_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_243 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08998_ _13848_/Q _14201_/Q _09005_/S vssd1 vssd1 vccd1 vccd1 _08998_/X sky130_fd_sc_hd__mux2_1
XFILLER_29_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07949_ _14745_/Q _07964_/A _07948_/Y _07949_/C1 vssd1 vssd1 vccd1 vccd1 _13552_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_75_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_67_clk clkbuf_5_11_0_clk/X vssd1 vssd1 vccd1 vccd1 _15579_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_28_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10960_ _13251_/B _11349_/C _11023_/A vssd1 vssd1 vccd1 vccd1 _10960_/X sky130_fd_sc_hd__mux2_1
XFILLER_28_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09619_ _13993_/Q _11874_/A1 _09628_/S vssd1 vssd1 vccd1 vccd1 _13993_/D sky130_fd_sc_hd__mux2_1
XFILLER_141_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10891_ _15532_/Q _06758_/Y _15533_/Q _06683_/Y vssd1 vssd1 vccd1 vccd1 _10891_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_188_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12630_ _15046_/Q _12629_/X _12834_/B vssd1 vssd1 vccd1 vccd1 _12630_/X sky130_fd_sc_hd__mux2_1
XFILLER_188_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12561_ _12618_/A1 _12556_/X _12559_/X _12560_/X _08405_/D vssd1 vssd1 vccd1 vccd1
+ _12573_/B sky130_fd_sc_hd__a221o_1
XFILLER_93_1095 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11512_ _13208_/B _11512_/B vssd1 vssd1 vccd1 vccd1 _11512_/X sky130_fd_sc_hd__and2b_1
XFILLER_157_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14300_ _15281_/CLK _14300_/D vssd1 vssd1 vccd1 vccd1 _14300_/Q sky130_fd_sc_hd__dfxtp_1
X_15280_ _15284_/CLK _15280_/D vssd1 vssd1 vccd1 vccd1 _15280_/Q sky130_fd_sc_hd__dfxtp_1
X_12492_ _12503_/A1 _12487_/X _12490_/X _12491_/X _08449_/A vssd1 vssd1 vccd1 vccd1
+ _12504_/B sky130_fd_sc_hd__a221o_1
XFILLER_156_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14231_ _15202_/CLK _14231_/D vssd1 vssd1 vccd1 vccd1 _14231_/Q sky130_fd_sc_hd__dfxtp_1
X_11443_ _11430_/X _11441_/X _11440_/Y vssd1 vssd1 vccd1 vccd1 _11443_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_109_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14162_ _15680_/CLK _14162_/D vssd1 vssd1 vccd1 vccd1 _14162_/Q sky130_fd_sc_hd__dfxtp_1
X_11374_ _11365_/B _11368_/B _11363_/X vssd1 vssd1 vccd1 vccd1 _11378_/A sky130_fd_sc_hd__a21oi_1
XFILLER_164_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13113_ _15524_/Q _13139_/S _13042_/A _13112_/X vssd1 vssd1 vccd1 vccd1 _15524_/D
+ sky130_fd_sc_hd__a22o_1
X_10325_ _07498_/C _13038_/S _10735_/S vssd1 vssd1 vccd1 vccd1 _14710_/D sky130_fd_sc_hd__mux2_1
X_14093_ _14093_/CLK _14093_/D vssd1 vssd1 vccd1 vccd1 _14093_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13044_ _06839_/X _12934_/Y _13043_/Y _06835_/X vssd1 vssd1 vccd1 vccd1 _13044_/X
+ sky130_fd_sc_hd__o211a_2
X_10256_ _14641_/Q _14794_/Q _10343_/S vssd1 vssd1 vccd1 vccd1 _14641_/D sky130_fd_sc_hd__mux2_1
XFILLER_26_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10187_ _11873_/A1 _14571_/Q _10197_/S vssd1 vssd1 vccd1 vccd1 _14571_/D sky130_fd_sc_hd__mux2_1
XFILLER_121_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_58_clk _15031_/CLK vssd1 vssd1 vccd1 vccd1 _14988_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_8_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14995_ _15556_/CLK _14995_/D vssd1 vssd1 vccd1 vccd1 _14995_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_4_11_0_clk clkbuf_3_5_0_clk/X vssd1 vssd1 vccd1 vccd1 clkbuf_5_23_0_clk/A
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_75_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13946_ _15652_/CLK _13946_/D vssd1 vssd1 vccd1 vccd1 _13946_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_71 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13877_ _15211_/CLK _13877_/D vssd1 vssd1 vccd1 vccd1 _13877_/Q sky130_fd_sc_hd__dfxtp_1
X_15616_ _15616_/CLK _15616_/D vssd1 vssd1 vccd1 vccd1 _15616_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12828_ _12828_/A _12828_/B vssd1 vssd1 vccd1 vccd1 _12828_/X sky130_fd_sc_hd__or2_1
XFILLER_188_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15547_ _15670_/CLK _15547_/D vssd1 vssd1 vccd1 vccd1 _15547_/Q sky130_fd_sc_hd__dfxtp_1
X_12759_ _15356_/Q _12759_/B vssd1 vssd1 vccd1 vccd1 _12759_/X sky130_fd_sc_hd__or2_1
XTAP_1291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15478_ _15518_/CLK _15478_/D vssd1 vssd1 vccd1 vccd1 _15478_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_147_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14429_ _15284_/CLK _14429_/D vssd1 vssd1 vccd1 vccd1 _14429_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_162_207 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09970_ _11857_/A1 _14329_/Q _09996_/S vssd1 vssd1 vccd1 vccd1 _14329_/D sky130_fd_sc_hd__mux2_1
XFILLER_171_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08921_ _14519_/Q _14132_/Q _14164_/Q _14100_/Q _08910_/S _08508_/B vssd1 vssd1 vccd1
+ vccd1 _08921_/X sky130_fd_sc_hd__mux4_1
XFILLER_170_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_115 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08852_ _09662_/B _08852_/B vssd1 vssd1 vccd1 vccd1 _11851_/A sky130_fd_sc_hd__nand2_8
XFILLER_112_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07803_ _13513_/Q _07798_/B _13514_/Q vssd1 vssd1 vccd1 vccd1 _07803_/Y sky130_fd_sc_hd__a21oi_1
X_08783_ _14712_/Q _08852_/B vssd1 vssd1 vccd1 vccd1 _13318_/D sky130_fd_sc_hd__or2_4
XFILLER_57_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_49_clk clkbuf_5_8_0_clk/X vssd1 vssd1 vccd1 vccd1 _14468_/CLK sky130_fd_sc_hd__clkbuf_16
X_07734_ _14753_/Q _07750_/A _07733_/Y _07987_/C1 vssd1 vssd1 vccd1 vccd1 _13496_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_2909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07665_ _13478_/Q _13477_/Q _07665_/C vssd1 vssd1 vccd1 vccd1 _07672_/C sky130_fd_sc_hd__and3_2
XFILLER_129_1103 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09404_ _09406_/S1 _09402_/X _09403_/X vssd1 vssd1 vccd1 vccd1 _09405_/C sky130_fd_sc_hd__a21o_1
XFILLER_80_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07596_ _07603_/C _07603_/D vssd1 vssd1 vccd1 vccd1 _07599_/B sky130_fd_sc_hd__and2_2
XFILLER_41_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09335_ _13896_/Q _13123_/B _08512_/B _14411_/Q _13123_/A vssd1 vssd1 vccd1 vccd1
+ _09335_/X sky130_fd_sc_hd__a221o_1
XFILLER_166_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09266_ _14440_/Q _08540_/B _08520_/B _09265_/X vssd1 vssd1 vccd1 vccd1 _09266_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_138_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_opt_1_0_clk clkbuf_5_7_0_clk/X vssd1 vssd1 vccd1 vccd1 clkbuf_opt_1_0_clk/X
+ sky130_fd_sc_hd__clkbuf_16
X_08217_ _13708_/Q _13346_/A0 _08221_/S vssd1 vssd1 vccd1 vccd1 _13708_/D sky130_fd_sc_hd__mux2_1
XFILLER_181_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09197_ _06676_/A _09186_/X _09195_/X _09196_/X vssd1 vssd1 vccd1 vccd1 _09197_/X
+ sky130_fd_sc_hd__o22a_2
XFILLER_181_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08148_ _13663_/Q _10285_/S _08119_/X _08147_/X vssd1 vssd1 vccd1 vccd1 _13663_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_14_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_112 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08079_ _14735_/Q _08083_/A _08078_/X _08084_/C1 vssd1 vssd1 vccd1 vccd1 _13645_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_150_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10110_ _14496_/Q _14744_/Q _10124_/S vssd1 vssd1 vccd1 vccd1 _14496_/D sky130_fd_sc_hd__mux2_1
XFILLER_171_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_947 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11090_ _11298_/A _11086_/X _11089_/X vssd1 vssd1 vccd1 vccd1 _11090_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_88_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10041_ _14398_/Q _13327_/A0 _10059_/S vssd1 vssd1 vccd1 vccd1 _14398_/D sky130_fd_sc_hd__mux2_1
XFILLER_49_917 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13800_ _14868_/CLK _13800_/D vssd1 vssd1 vccd1 vccd1 _13800_/Q sky130_fd_sc_hd__dfxtp_1
X_14780_ _15632_/CLK _14780_/D vssd1 vssd1 vccd1 vccd1 _14780_/Q sky130_fd_sc_hd__dfxtp_1
X_11992_ _11992_/A _11992_/B vssd1 vssd1 vccd1 vccd1 _11992_/X sky130_fd_sc_hd__and2_1
X_10943_ _14956_/Q _10948_/B _10942_/Y _13236_/B vssd1 vssd1 vccd1 vccd1 _14956_/D
+ sky130_fd_sc_hd__o22a_1
X_13731_ _15540_/CLK _13731_/D vssd1 vssd1 vccd1 vccd1 _13731_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_28_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_3_0_0_clk clkbuf_3_1_0_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_1_0_clk/A sky130_fd_sc_hd__clkbuf_8
X_10874_ _13732_/Q _14906_/Q _13129_/A vssd1 vssd1 vccd1 vccd1 _14906_/D sky130_fd_sc_hd__mux2_1
X_13662_ _14703_/CLK _13662_/D vssd1 vssd1 vccd1 vccd1 _13662_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_188_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15401_ _15620_/CLK _15401_/D vssd1 vssd1 vccd1 vccd1 _15401_/Q sky130_fd_sc_hd__dfxtp_2
X_12613_ _12613_/A _12613_/B vssd1 vssd1 vccd1 vccd1 _12613_/X sky130_fd_sc_hd__and2_1
X_13593_ _15630_/CLK _13593_/D vssd1 vssd1 vccd1 vccd1 _13593_/Q sky130_fd_sc_hd__dfxtp_2
XPHY_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_40 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12544_ _12544_/A _12544_/B vssd1 vssd1 vccd1 vccd1 _12544_/X sky130_fd_sc_hd__and2_1
X_15332_ _15332_/CLK _15332_/D vssd1 vssd1 vccd1 vccd1 _15332_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_177_40 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_579 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15263_ _15295_/CLK _15263_/D vssd1 vssd1 vccd1 vccd1 _15263_/Q sky130_fd_sc_hd__dfxtp_1
X_12475_ _12498_/A _12475_/B vssd1 vssd1 vccd1 vccd1 _12475_/X sky130_fd_sc_hd__and2_1
XFILLER_184_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11426_ _11425_/Y _15051_/Q _11474_/S vssd1 vssd1 vccd1 vccd1 _15051_/D sky130_fd_sc_hd__mux2_1
X_14214_ _15301_/CLK _14214_/D vssd1 vssd1 vccd1 vccd1 _14214_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_137_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15194_ _15295_/CLK _15194_/D vssd1 vssd1 vccd1 vccd1 _15194_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_6 _08744_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14145_ _15663_/CLK _14145_/D vssd1 vssd1 vccd1 vccd1 _14145_/Q sky130_fd_sc_hd__dfxtp_1
X_11357_ _13159_/B _11357_/B _11357_/C vssd1 vssd1 vccd1 vccd1 _11359_/A sky130_fd_sc_hd__and3_1
XFILLER_153_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10308_ _14693_/Q _14878_/Q _10650_/S vssd1 vssd1 vccd1 vccd1 _14693_/D sky130_fd_sc_hd__mux2_1
XFILLER_152_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14076_ _15184_/CLK _14076_/D vssd1 vssd1 vccd1 vccd1 _14076_/Q sky130_fd_sc_hd__dfxtp_1
X_11288_ _11330_/A _11272_/Y _11287_/X vssd1 vssd1 vccd1 vccd1 _11288_/X sky130_fd_sc_hd__a21o_1
X_13027_ _07484_/X _13039_/A2 _13026_/X _12944_/A vssd1 vssd1 vccd1 vccd1 _13027_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_112_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10239_ _14624_/Q _14777_/Q _10650_/S vssd1 vssd1 vccd1 vccd1 _14624_/D sky130_fd_sc_hd__mux2_1
XFILLER_121_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14978_ _15020_/CLK _14978_/D vssd1 vssd1 vccd1 vccd1 _14978_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13929_ _15678_/CLK _13929_/D vssd1 vssd1 vccd1 vccd1 _13929_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_19_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07450_ _14664_/Q _07474_/B _07482_/C vssd1 vssd1 vccd1 vccd1 _07450_/X sky130_fd_sc_hd__and3_1
XFILLER_179_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07381_ _11853_/A1 _13384_/Q _07501_/S vssd1 vssd1 vccd1 vccd1 _13384_/D sky130_fd_sc_hd__mux2_1
XFILLER_15_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09120_ _09445_/C1 _09117_/X _09119_/X _09130_/A vssd1 vssd1 vccd1 vccd1 _09120_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_187_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09051_ _14525_/Q _14138_/Q _14170_/Q _14106_/Q _09407_/S _09406_/S1 vssd1 vssd1
+ vccd1 vccd1 _09051_/X sky130_fd_sc_hd__mux4_1
XFILLER_163_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_771 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08002_ _14759_/Q _08022_/B _08001_/X _08002_/C1 vssd1 vssd1 vccd1 vccd1 _13566_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_116_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_295 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09953_ _11873_/A1 _14313_/Q _09963_/S vssd1 vssd1 vccd1 vccd1 _14313_/D sky130_fd_sc_hd__mux2_1
XFILLER_104_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08904_ _13907_/Q _08903_/X _12504_/A vssd1 vssd1 vccd1 vccd1 _13907_/D sky130_fd_sc_hd__mux2_1
XFILLER_44_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09884_ _07448_/X _14246_/Q _09897_/S vssd1 vssd1 vccd1 vccd1 _14246_/D sky130_fd_sc_hd__mux2_1
XTAP_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08835_ _13858_/Q _13334_/A0 _08846_/S vssd1 vssd1 vccd1 vccd1 _13858_/D sky130_fd_sc_hd__mux2_1
XFILLER_97_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08766_ _08758_/X _08759_/X _08764_/X _08765_/X _08763_/X vssd1 vssd1 vccd1 vccd1
+ _08766_/X sky130_fd_sc_hd__a221o_1
XFILLER_85_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07717_ _07717_/A _07717_/B _07732_/B vssd1 vssd1 vccd1 vccd1 _07724_/C sky130_fd_sc_hd__and3_2
XTAP_2728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08697_ _13573_/Q _08724_/B _08724_/C vssd1 vssd1 vccd1 vccd1 _08697_/X sky130_fd_sc_hd__and3_1
XTAP_2739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_750 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07648_ _07646_/Y _07650_/B _07651_/A vssd1 vssd1 vccd1 vccd1 _07648_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_26_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07579_ _13456_/Q _07588_/D vssd1 vssd1 vccd1 vccd1 _07579_/Y sky130_fd_sc_hd__nor2_1
X_09318_ _14538_/Q _14151_/Q _14183_/Q _14119_/Q _09481_/S _08519_/A vssd1 vssd1 vccd1
+ vccd1 _09318_/X sky130_fd_sc_hd__mux4_1
XFILLER_139_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10590_ _14736_/Q _10589_/X _10735_/S vssd1 vssd1 vccd1 vccd1 _14736_/D sky130_fd_sc_hd__mux2_1
XFILLER_139_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09249_ _14020_/Q _13988_/Q _09484_/S vssd1 vssd1 vccd1 vccd1 _09249_/X sky130_fd_sc_hd__mux2_1
XFILLER_21_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12260_ _12260_/A _12260_/B vssd1 vssd1 vccd1 vccd1 _12260_/X sky130_fd_sc_hd__or2_1
XFILLER_154_549 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11211_ _10399_/B _15000_/Q _11237_/S vssd1 vssd1 vccd1 vccd1 _15000_/D sky130_fd_sc_hd__mux2_1
X_12191_ _12490_/A _12191_/B vssd1 vssd1 vccd1 vccd1 _12191_/X sky130_fd_sc_hd__or2_1
XFILLER_108_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11142_ _11062_/X _11067_/X _11283_/A vssd1 vssd1 vccd1 vccd1 _11142_/X sky130_fd_sc_hd__mux2_1
Xoutput43 _07179_/X vssd1 vssd1 vccd1 vccd1 ext_address[17] sky130_fd_sc_hd__clkbuf_2
Xoutput54 _07190_/X vssd1 vssd1 vccd1 vccd1 ext_address[28] sky130_fd_sc_hd__clkbuf_2
Xoutput65 _07171_/X vssd1 vssd1 vccd1 vccd1 ext_address[9] sky130_fd_sc_hd__clkbuf_2
Xoutput76 _07137_/X vssd1 vssd1 vccd1 vccd1 ext_write_data[18] sky130_fd_sc_hd__clkbuf_2
Xoutput87 _07157_/X vssd1 vssd1 vccd1 vccd1 ext_write_data[28] sky130_fd_sc_hd__clkbuf_2
X_11073_ _14964_/Q _11202_/A _11064_/Y _11072_/Y vssd1 vssd1 vccd1 vccd1 _14964_/D
+ sky130_fd_sc_hd__o22a_1
Xoutput98 _07119_/X vssd1 vssd1 vccd1 vccd1 ext_write_data[9] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10024_ _13345_/A0 _14382_/Q _10028_/S vssd1 vssd1 vccd1 vccd1 _14382_/D sky130_fd_sc_hd__mux2_1
X_14901_ _15616_/CLK _14901_/D vssd1 vssd1 vccd1 vccd1 _14901_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_76_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14832_ _15536_/CLK _14832_/D vssd1 vssd1 vccd1 vccd1 _14832_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_3930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14763_ _15623_/CLK _14763_/D vssd1 vssd1 vccd1 vccd1 _14763_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_3974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11975_ _12596_/A _11975_/B _11975_/C vssd1 vssd1 vccd1 vccd1 _11975_/X sky130_fd_sc_hd__and3_2
XFILLER_56_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13714_ _14468_/CLK _13714_/D vssd1 vssd1 vccd1 vccd1 _13714_/Q sky130_fd_sc_hd__dfxtp_1
X_10926_ _11536_/B _10925_/X _10929_/B _14946_/Q vssd1 vssd1 vccd1 vccd1 _14946_/D
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_186_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14694_ _15643_/CLK _14694_/D vssd1 vssd1 vccd1 vccd1 _14694_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10857_ _14889_/Q _13779_/Q _12933_/S vssd1 vssd1 vccd1 vccd1 _14889_/D sky130_fd_sc_hd__mux2_1
X_13645_ _15372_/CLK _13645_/D vssd1 vssd1 vccd1 vccd1 _13645_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10788_ _14820_/Q _15452_/Q _12929_/S vssd1 vssd1 vccd1 vccd1 _14820_/D sky130_fd_sc_hd__mux2_1
XPHY_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13576_ _13803_/CLK _13576_/D vssd1 vssd1 vccd1 vccd1 _13576_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_173_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15315_ _15315_/CLK _15315_/D vssd1 vssd1 vccd1 vccd1 _15315_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_145_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12527_ _13134_/A _12527_/B _12527_/C vssd1 vssd1 vccd1 vccd1 _12527_/X sky130_fd_sc_hd__and3_1
XFILLER_145_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15246_ _15278_/CLK _15246_/D vssd1 vssd1 vccd1 vccd1 _15246_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_184_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12458_ _12596_/A _12458_/B _12458_/C vssd1 vssd1 vccd1 vccd1 _12458_/X sky130_fd_sc_hd__and3_1
XFILLER_160_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11409_ _13178_/B _11409_/B vssd1 vssd1 vccd1 vccd1 _11410_/B sky130_fd_sc_hd__nand2_1
X_15177_ _15278_/CLK _15177_/D vssd1 vssd1 vccd1 vccd1 _15177_/Q sky130_fd_sc_hd__dfxtp_1
X_12389_ _13134_/A _12389_/B _12389_/C vssd1 vssd1 vccd1 vccd1 _12389_/X sky130_fd_sc_hd__and3_1
XFILLER_99_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14128_ _15678_/CLK _14128_/D vssd1 vssd1 vccd1 vccd1 _14128_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_154_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06950_ _14489_/Q _06748_/Y _06750_/Y _13479_/Q vssd1 vssd1 vccd1 vccd1 _06960_/A
+ sky130_fd_sc_hd__a2bb2o_1
X_14059_ _14542_/CLK _14059_/D vssd1 vssd1 vccd1 vccd1 _14059_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06881_ _14510_/Q _06705_/Y _06878_/X _06879_/Y _06880_/X vssd1 vssd1 vccd1 vccd1
+ _06882_/D sky130_fd_sc_hd__a2111o_1
X_08620_ _13787_/Q _08626_/S _08619_/X vssd1 vssd1 vccd1 vccd1 _13787_/D sky130_fd_sc_hd__o21a_1
XFILLER_95_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08551_ _14515_/Q _08748_/B1 _08549_/X _08550_/X vssd1 vssd1 vccd1 vccd1 _08552_/C
+ sky130_fd_sc_hd__a211o_1
X_07502_ _14722_/Q _14721_/Q _14724_/Q _14723_/Q vssd1 vssd1 vccd1 vccd1 _07504_/C
+ sky130_fd_sc_hd__or4_1
XFILLER_74_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08482_ hold4/A _08465_/B _08477_/X _08451_/A _08481_/X vssd1 vssd1 vccd1 vccd1 _08482_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_50_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07433_ _13333_/A0 _13397_/Q _07481_/S vssd1 vssd1 vccd1 vccd1 _13397_/D sky130_fd_sc_hd__mux2_1
XFILLER_74_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07364_ _07355_/A _07363_/X _07359_/X _07355_/X vssd1 vssd1 vccd1 vccd1 _07365_/B
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_176_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09103_ _14238_/Q _14270_/Q _14302_/Q _14334_/Q _09444_/S _09448_/S1 vssd1 vssd1
+ vccd1 vccd1 _09103_/X sky130_fd_sc_hd__mux4_2
XFILLER_148_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07295_ _15316_/Q _15472_/Q _07340_/S vssd1 vssd1 vccd1 vccd1 _07295_/X sky130_fd_sc_hd__mux2_4
XFILLER_175_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09034_ _09524_/A _09027_/X _09030_/X _08501_/A vssd1 vssd1 vccd1 vccd1 _09034_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_164_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_172_880 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09936_ _13323_/A0 _14296_/Q _09958_/S vssd1 vssd1 vccd1 vccd1 _14296_/D sky130_fd_sc_hd__mux2_1
XFILLER_86_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09867_ _11853_/A1 _14229_/Q _09897_/S vssd1 vssd1 vccd1 vccd1 _14229_/D sky130_fd_sc_hd__mux2_1
XTAP_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08818_ _14714_/Q _14715_/Q _14716_/Q _08817_/B vssd1 vssd1 vccd1 vccd1 _10065_/A
+ sky130_fd_sc_hd__o31a_4
XTAP_3226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09798_ _14164_/Q _13320_/A0 _09828_/S vssd1 vssd1 vccd1 vccd1 _14164_/D sky130_fd_sc_hd__mux2_1
XTAP_3237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08749_ _13580_/Q _08749_/A2 _08748_/X vssd1 vssd1 vccd1 vccd1 _08749_/X sky130_fd_sc_hd__a21o_1
XTAP_2525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11760_ _11868_/A1 _15188_/Q _11774_/S vssd1 vssd1 vccd1 vccd1 _15188_/D sky130_fd_sc_hd__mux2_1
XFILLER_60_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_411 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10711_ _15021_/Q _10569_/B _10718_/A2 _14989_/Q _10732_/C1 vssd1 vssd1 vccd1 vccd1
+ _10711_/X sky130_fd_sc_hd__a221o_1
XFILLER_13_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11691_ _13333_/A0 _15122_/Q _11703_/S vssd1 vssd1 vccd1 vccd1 _15122_/D sky130_fd_sc_hd__mux2_1
XTAP_1868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13430_ _15381_/CLK _13430_/D vssd1 vssd1 vccd1 vccd1 _13430_/Q sky130_fd_sc_hd__dfxtp_2
X_10642_ _15007_/Q _10717_/A2 _10602_/B _13726_/Q _10717_/C1 vssd1 vssd1 vccd1 vccd1
+ _10642_/X sky130_fd_sc_hd__a221o_1
XFILLER_139_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13361_ _14464_/Q vssd1 vssd1 vccd1 vccd1 _14464_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_182_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10573_ _14929_/Q _14928_/Q _14927_/Q vssd1 vssd1 vccd1 vccd1 _10573_/X sky130_fd_sc_hd__and3_2
XFILLER_127_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15100_ _15673_/CLK _15100_/D vssd1 vssd1 vccd1 vccd1 _15100_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_154_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12312_ _12592_/A1 _12311_/X _12536_/A vssd1 vssd1 vccd1 vccd1 _12312_/X sky130_fd_sc_hd__a21o_1
X_13292_ _12667_/Y _15624_/Q _13309_/A vssd1 vssd1 vccd1 vccd1 _15624_/D sky130_fd_sc_hd__mux2_1
XFILLER_177_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15031_ _15031_/CLK _15031_/D vssd1 vssd1 vccd1 vccd1 _15031_/Q sky130_fd_sc_hd__dfxtp_2
X_12243_ _12477_/A1 _12242_/X _12490_/A vssd1 vssd1 vccd1 vccd1 _12243_/X sky130_fd_sc_hd__a21o_1
XFILLER_5_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_711 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12174_ _12477_/A1 _12173_/X _12502_/S vssd1 vssd1 vccd1 vccd1 _12174_/X sky130_fd_sc_hd__a21o_1
XFILLER_174_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11125_ _11047_/Y _11085_/X _11088_/X _08249_/Y _11380_/A vssd1 vssd1 vccd1 vccd1
+ _11125_/X sky130_fd_sc_hd__a221o_1
XFILLER_7_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11056_ _10960_/X _11055_/Y _11330_/A vssd1 vssd1 vccd1 vccd1 _11056_/X sky130_fd_sc_hd__mux2_1
XFILLER_3_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10007_ _11861_/A1 _14365_/Q _10028_/S vssd1 vssd1 vccd1 vccd1 _14365_/D sky130_fd_sc_hd__mux2_1
XFILLER_67_94 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14815_ _15634_/CLK _14815_/D vssd1 vssd1 vccd1 vccd1 _14815_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_97_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14746_ _15592_/CLK _14746_/D vssd1 vssd1 vccd1 vccd1 _14746_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_3793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_474 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11958_ _11954_/X _11955_/X _12582_/A vssd1 vssd1 vccd1 vccd1 _11958_/X sky130_fd_sc_hd__mux2_1
X_10909_ _14937_/Q _10908_/Y _10951_/B vssd1 vssd1 vccd1 vccd1 _14937_/D sky130_fd_sc_hd__mux2_1
X_14677_ _15462_/CLK _14677_/D vssd1 vssd1 vccd1 vccd1 _14677_/Q sky130_fd_sc_hd__dfxtp_1
X_11889_ _11885_/X _11886_/X _12260_/A vssd1 vssd1 vccd1 vccd1 _11889_/X sky130_fd_sc_hd__mux2_1
XFILLER_32_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13628_ _15381_/CLK _13628_/D vssd1 vssd1 vccd1 vccd1 _13628_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_177_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13559_ _15386_/CLK _13559_/D vssd1 vssd1 vccd1 vccd1 _13559_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_173_600 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1066 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07080_ _07079_/X _14759_/Q _07098_/S vssd1 vssd1 vccd1 vccd1 _13605_/D sky130_fd_sc_hd__mux2_1
XFILLER_146_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15229_ _15292_/CLK _15229_/D vssd1 vssd1 vccd1 vccd1 _15229_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_161_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout107 _13288_/S vssd1 vssd1 vccd1 vccd1 _13284_/S sky130_fd_sc_hd__buf_12
Xfanout118 _12944_/Y vssd1 vssd1 vccd1 vccd1 _13039_/A2 sky130_fd_sc_hd__buf_8
XFILLER_87_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07982_ _07971_/A _07981_/X input35/X vssd1 vssd1 vccd1 vccd1 _07982_/Y sky130_fd_sc_hd__a21oi_1
Xfanout129 fanout138/X vssd1 vssd1 vccd1 vccd1 _10759_/S sky130_fd_sc_hd__buf_12
XFILLER_141_596 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06933_ _06734_/Y _13486_/Q _06736_/Y _13485_/Q vssd1 vssd1 vccd1 vccd1 _06944_/A
+ sky130_fd_sc_hd__a22o_2
X_09721_ _13343_/A0 _14091_/Q _09723_/S vssd1 vssd1 vccd1 vccd1 _14091_/D sky130_fd_sc_hd__mux2_1
XFILLER_86_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09652_ _14025_/Q _13341_/A0 _09661_/S vssd1 vssd1 vccd1 vccd1 _14025_/D sky130_fd_sc_hd__mux2_1
XFILLER_27_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06864_ input35/X _12622_/A vssd1 vssd1 vccd1 vccd1 _06997_/B sky130_fd_sc_hd__nor2_4
XFILLER_28_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08603_ _13601_/Q _08691_/A2 _08685_/A2 _13562_/Q vssd1 vssd1 vccd1 vccd1 _08603_/X
+ sky130_fd_sc_hd__a22o_1
X_09583_ _13959_/Q _11872_/A1 _09594_/S vssd1 vssd1 vccd1 vccd1 _13959_/D sky130_fd_sc_hd__mux2_1
X_06795_ _14596_/Q _14595_/Q vssd1 vssd1 vccd1 vccd1 _08756_/B sky130_fd_sc_hd__or2_4
XFILLER_83_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08534_ _13572_/Q _08747_/A2 _08533_/X _08722_/A vssd1 vssd1 vccd1 vccd1 _08534_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_63_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08465_ _14589_/Q _08465_/B vssd1 vssd1 vccd1 vccd1 _08465_/X sky130_fd_sc_hd__and2b_2
XFILLER_51_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_438 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07416_ _14744_/Q _07415_/X _07480_/S vssd1 vssd1 vccd1 vccd1 _07416_/X sky130_fd_sc_hd__mux2_8
XFILLER_144_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08396_ _13730_/Q _13140_/S _08394_/X hold4/X vssd1 vssd1 vccd1 vccd1 _13730_/D sky130_fd_sc_hd__a22o_1
XFILLER_177_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07347_ _07345_/Y _07360_/D _07360_/A vssd1 vssd1 vccd1 vccd1 _07347_/X sky130_fd_sc_hd__o21ba_1
XFILLER_10_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07278_ _07278_/A _07278_/B vssd1 vssd1 vccd1 vccd1 _07278_/X sky130_fd_sc_hd__and2_1
XFILLER_128_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09017_ _09532_/A _09017_/B vssd1 vssd1 vccd1 vccd1 _09017_/X sky130_fd_sc_hd__or2_1
XFILLER_163_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_582 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_253_clk clkbuf_5_1_0_clk/X vssd1 vssd1 vccd1 vccd1 _15172_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_78_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout630 _14195_/Q vssd1 vssd1 vccd1 vccd1 _10515_/B2 sky130_fd_sc_hd__buf_12
XFILLER_137_1098 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout641 fanout647/X vssd1 vssd1 vccd1 vccd1 _08016_/C1 sky130_fd_sc_hd__buf_8
X_09919_ _13339_/A0 _14280_/Q _09930_/S vssd1 vssd1 vccd1 vccd1 _14280_/D sky130_fd_sc_hd__mux2_1
XFILLER_77_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12930_ _15458_/Q _15644_/Q _12933_/S vssd1 vssd1 vccd1 vccd1 _15458_/D sky130_fd_sc_hd__mux2_1
XTAP_3001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12861_ _14755_/Q _15389_/Q _12871_/S vssd1 vssd1 vccd1 vccd1 _15389_/D sky130_fd_sc_hd__mux2_1
XFILLER_18_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14600_ _15612_/CLK _14600_/D vssd1 vssd1 vccd1 vccd1 _14600_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_3089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11812_ _15235_/Q _13104_/B2 _11816_/S vssd1 vssd1 vccd1 vccd1 _15235_/D sky130_fd_sc_hd__mux2_1
XTAP_2344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15580_ _15580_/CLK _15580_/D vssd1 vssd1 vccd1 vccd1 _15580_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12792_ _15068_/Q _12792_/B vssd1 vssd1 vccd1 vccd1 _12792_/X sky130_fd_sc_hd__or2_1
XTAP_1621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14531_ _15659_/CLK _14531_/D vssd1 vssd1 vccd1 vccd1 _14531_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11743_ _14714_/Q _14716_/Q _11743_/C _11818_/A vssd1 vssd1 vccd1 vccd1 _11743_/X
+ sky130_fd_sc_hd__or4_4
XTAP_2399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_904 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_1088 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14462_ _14462_/CLK _14462_/D vssd1 vssd1 vccd1 vccd1 _14462_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11674_ _13349_/A0 _15106_/Q _11675_/S vssd1 vssd1 vccd1 vccd1 _15106_/D sky130_fd_sc_hd__mux2_1
XFILLER_53_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13413_ _15678_/CLK _13413_/D vssd1 vssd1 vccd1 vccd1 _13413_/Q sky130_fd_sc_hd__dfxtp_1
X_10625_ _14743_/Q _10624_/X _10710_/S vssd1 vssd1 vccd1 vccd1 _14743_/D sky130_fd_sc_hd__mux2_1
XFILLER_155_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14393_ _15202_/CLK _14393_/D vssd1 vssd1 vccd1 vccd1 _14393_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_183_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13344_ _13344_/A0 _15674_/Q _13345_/S vssd1 vssd1 vccd1 vccd1 _15674_/D sky130_fd_sc_hd__mux2_1
X_10556_ _10556_/A _10556_/B _10556_/C _10556_/D vssd1 vssd1 vccd1 vccd1 _10557_/C
+ sky130_fd_sc_hd__or4_2
XFILLER_128_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13275_ _15359_/Q _15606_/Q _13309_/A vssd1 vssd1 vccd1 vccd1 _15606_/D sky130_fd_sc_hd__mux2_1
X_10487_ _10507_/A1 _13752_/Q _15420_/Q _10515_/B2 vssd1 vssd1 vccd1 vccd1 _10487_/X
+ sky130_fd_sc_hd__a22o_1
X_15014_ _15014_/CLK _15014_/D vssd1 vssd1 vccd1 vccd1 _15014_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_170_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12226_ _12209_/X _12210_/X _12260_/A vssd1 vssd1 vccd1 vccd1 _12226_/X sky130_fd_sc_hd__mux2_1
XFILLER_135_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_244_clk clkbuf_5_4_0_clk/X vssd1 vssd1 vccd1 vccd1 _14470_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_64_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12157_ _12140_/X _12141_/X _12260_/A vssd1 vssd1 vccd1 vccd1 _12157_/X sky130_fd_sc_hd__mux2_1
XFILLER_78_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11108_ _11307_/A _11046_/X _11048_/Y _11035_/X _11414_/A vssd1 vssd1 vccd1 vccd1
+ _11108_/X sky130_fd_sc_hd__o221a_1
X_12088_ _12071_/X _12072_/X _12582_/A vssd1 vssd1 vccd1 vccd1 _12088_/X sky130_fd_sc_hd__mux2_1
X_11039_ _11036_/Y _11038_/Y _11330_/A vssd1 vssd1 vccd1 vccd1 _11039_/X sky130_fd_sc_hd__mux2_1
XFILLER_49_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14729_ _15615_/CLK _14729_/D vssd1 vssd1 vccd1 vccd1 _14729_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_33_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08250_ _11298_/A _11047_/B vssd1 vssd1 vccd1 vccd1 _11307_/A sky130_fd_sc_hd__nand2_8
XFILLER_33_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07201_ _07201_/A vssd1 vssd1 vccd1 vccd1 _07228_/B sky130_fd_sc_hd__inv_2
XFILLER_177_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08181_ _08150_/S input22/X _08185_/A vssd1 vssd1 vccd1 vccd1 _08181_/X sky130_fd_sc_hd__and3b_1
X_07132_ _14846_/Q _14838_/Q _07146_/S vssd1 vssd1 vccd1 vccd1 _07132_/X sky130_fd_sc_hd__mux2_1
XFILLER_119_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07063_ _14633_/Q _14665_/Q _07078_/S vssd1 vssd1 vccd1 vccd1 _07063_/X sky130_fd_sc_hd__mux2_1
XFILLER_146_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_235_clk clkbuf_5_5_0_clk/X vssd1 vssd1 vccd1 vccd1 _15652_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_99_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07965_ _14749_/Q _07964_/A _07964_/Y _07965_/C1 vssd1 vssd1 vccd1 vccd1 _13556_/D
+ sky130_fd_sc_hd__o211a_1
X_09704_ _13326_/A0 _14074_/Q _09723_/S vssd1 vssd1 vccd1 vccd1 _14074_/D sky130_fd_sc_hd__mux2_1
XFILLER_96_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06916_ _06712_/Y _13465_/Q _06714_/Y _13464_/Q vssd1 vssd1 vccd1 vccd1 _06916_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_114_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07896_ _14763_/Q _07903_/A _07895_/X _08012_/C1 vssd1 vssd1 vccd1 vccd1 _13538_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_74_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09635_ _14008_/Q _11857_/A1 _09661_/S vssd1 vssd1 vccd1 vccd1 _14008_/D sky130_fd_sc_hd__mux2_1
XFILLER_56_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06847_ _06806_/A _06844_/X _06846_/X _06840_/X vssd1 vssd1 vccd1 vccd1 _06847_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_82_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09566_ _13942_/Q _11680_/A0 _09589_/S vssd1 vssd1 vccd1 vccd1 _13942_/D sky130_fd_sc_hd__mux2_1
X_06778_ _07096_/S _14730_/Q vssd1 vssd1 vccd1 vccd1 _10566_/B sky130_fd_sc_hd__and2_4
X_08517_ _08517_/A _08528_/C vssd1 vssd1 vccd1 vccd1 _08521_/A sky130_fd_sc_hd__or2_4
XFILLER_24_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09497_ _15302_/Q _15270_/Q _15238_/Q _15169_/Q _09512_/S _09511_/S1 vssd1 vssd1
+ vccd1 vccd1 _09497_/X sky130_fd_sc_hd__mux4_1
XFILLER_70_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_224 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08448_ _13754_/Q _12878_/S _08426_/B _08447_/X vssd1 vssd1 vccd1 vccd1 _13754_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_139_11 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_44 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08379_ _11347_/A _08299_/B _08299_/C _08378_/Y vssd1 vssd1 vccd1 vccd1 _08379_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_149_471 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1083 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10410_ _10410_/A _10410_/B vssd1 vssd1 vccd1 vccd1 _10555_/B sky130_fd_sc_hd__nand2_1
XFILLER_165_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11390_ _13171_/B _11390_/B _11390_/C vssd1 vssd1 vccd1 vccd1 _11401_/B sky130_fd_sc_hd__nand3_2
XFILLER_165_964 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_901 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10341_ _14726_/Q _14919_/Q _10343_/S vssd1 vssd1 vccd1 vccd1 _14726_/D sky130_fd_sc_hd__mux2_1
XFILLER_164_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13060_ _12957_/X _13104_/A2 _13104_/B1 _07392_/X vssd1 vssd1 vccd1 vccd1 _13060_/X
+ sky130_fd_sc_hd__a22o_1
X_10272_ _14657_/Q _14810_/Q _10650_/S vssd1 vssd1 vccd1 vccd1 _14657_/D sky130_fd_sc_hd__mux2_1
XFILLER_180_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12011_ _12590_/A _12011_/B vssd1 vssd1 vccd1 vccd1 _12011_/X sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_226_clk clkbuf_5_7_0_clk/X vssd1 vssd1 vccd1 vccd1 _14542_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_155_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout460 _09450_/B1 vssd1 vssd1 vccd1 vccd1 _08501_/A sky130_fd_sc_hd__buf_12
Xfanout471 _06671_/Y vssd1 vssd1 vccd1 vccd1 _12618_/A1 sky130_fd_sc_hd__buf_12
XFILLER_24_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout482 _06669_/Y vssd1 vssd1 vccd1 vccd1 _12500_/A1 sky130_fd_sc_hd__buf_12
XFILLER_4_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13962_ _15328_/CLK _13962_/D vssd1 vssd1 vccd1 vccd1 _13962_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout493 _15043_/Q vssd1 vssd1 vccd1 vccd1 _07146_/S sky130_fd_sc_hd__buf_12
X_12913_ _15441_/Q _15627_/Q _12918_/S vssd1 vssd1 vccd1 vccd1 _15441_/D sky130_fd_sc_hd__mux2_1
XFILLER_171_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13893_ _15094_/CLK _13893_/D vssd1 vssd1 vccd1 vccd1 _13893_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15632_ _15632_/CLK _15632_/D vssd1 vssd1 vccd1 vccd1 _15632_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12844_ _14738_/Q _15372_/Q _12871_/S vssd1 vssd1 vccd1 vccd1 _15372_/D sky130_fd_sc_hd__mux2_1
XTAP_2141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15563_ _15570_/CLK _15563_/D vssd1 vssd1 vccd1 vccd1 _15563_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12775_ _15359_/Q _12776_/B vssd1 vssd1 vccd1 vccd1 _12789_/C sky130_fd_sc_hd__and2_1
XTAP_1451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14514_ _15398_/CLK _14514_/D vssd1 vssd1 vccd1 vccd1 _14514_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_42_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11726_ _15155_/Q _13334_/A0 _11741_/S vssd1 vssd1 vccd1 vccd1 _15155_/D sky130_fd_sc_hd__mux2_1
XTAP_1495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15494_ _15507_/CLK _15494_/D vssd1 vssd1 vccd1 vccd1 _15494_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_159_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14445_ _15517_/CLK _14445_/D vssd1 vssd1 vccd1 vccd1 _14445_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11657_ _13332_/A0 _15089_/Q _11670_/S vssd1 vssd1 vccd1 vccd1 _15089_/D sky130_fd_sc_hd__mux2_1
XFILLER_70_1074 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10608_ _14968_/Q _10733_/A2 _10733_/B1 _14936_/Q _10607_/X vssd1 vssd1 vccd1 vccd1
+ _10608_/X sky130_fd_sc_hd__a221o_2
X_14376_ _15192_/CLK _14376_/D vssd1 vssd1 vccd1 vccd1 _14376_/Q sky130_fd_sc_hd__dfxtp_1
X_11588_ _15067_/Q _11614_/S _11586_/Y _11587_/X vssd1 vssd1 vccd1 vccd1 _15067_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_7_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13327_ _13327_/A0 _15657_/Q _13345_/S vssd1 vssd1 vccd1 vccd1 _15657_/D sky130_fd_sc_hd__mux2_1
X_10539_ _11536_/A _13208_/B _10519_/B _10538_/X vssd1 vssd1 vccd1 vccd1 _10539_/Y
+ sky130_fd_sc_hd__a211oi_1
XFILLER_155_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13258_ _15342_/Q _15589_/Q _13282_/S vssd1 vssd1 vccd1 vccd1 _15589_/D sky130_fd_sc_hd__mux2_1
XFILLER_170_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_217_clk clkbuf_5_18_0_clk/X vssd1 vssd1 vccd1 vccd1 _15328_/CLK sky130_fd_sc_hd__clkbuf_16
X_12209_ _14532_/Q _14145_/Q _14177_/Q _14113_/Q _12472_/S _12465_/S1 vssd1 vssd1
+ vccd1 vccd1 _12209_/X sky130_fd_sc_hd__mux4_1
X_13189_ _13229_/A _13189_/B vssd1 vssd1 vccd1 vccd1 _13189_/Y sky130_fd_sc_hd__nor2_1
XFILLER_151_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07750_ _07750_/A _07750_/B vssd1 vssd1 vccd1 vccd1 _07750_/Y sky130_fd_sc_hd__nand2_1
XFILLER_38_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06701_ _13471_/Q vssd1 vssd1 vccd1 vccd1 _06701_/Y sky130_fd_sc_hd__inv_2
XFILLER_93_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07681_ _14739_/Q _07676_/A _07680_/Y _07938_/C1 vssd1 vssd1 vccd1 vccd1 _13482_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_64_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09420_ _14479_/Q _09536_/A2 _13130_/B1 _14447_/Q _09419_/X vssd1 vssd1 vccd1 vccd1
+ _09420_/X sky130_fd_sc_hd__a221o_1
XFILLER_18_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09351_ _08507_/A _09350_/X _09349_/X _09524_/A vssd1 vssd1 vccd1 vccd1 _09351_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_178_500 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_1080 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08302_ _10507_/A1 _13767_/Q _15405_/Q _10515_/B2 vssd1 vssd1 vccd1 vccd1 _08302_/X
+ sky130_fd_sc_hd__a22o_1
X_09282_ _13925_/Q _13149_/S _09281_/X vssd1 vssd1 vccd1 vccd1 _13925_/D sky130_fd_sc_hd__a21o_1
XFILLER_100_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08233_ _11302_/A _08233_/B vssd1 vssd1 vccd1 vccd1 _11327_/A sky130_fd_sc_hd__nand2_1
XFILLER_21_767 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08164_ _13669_/Q _10695_/S _08155_/X _08163_/X vssd1 vssd1 vccd1 vccd1 _13669_/D
+ sky130_fd_sc_hd__o22a_1
X_07115_ _14837_/Q _07115_/B _07163_/A vssd1 vssd1 vccd1 vccd1 _07115_/X sky130_fd_sc_hd__and3_4
XFILLER_106_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08095_ _08151_/S _08095_/B vssd1 vssd1 vccd1 vccd1 _08095_/X sky130_fd_sc_hd__or2_1
XFILLER_107_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07046_ _07045_/X _13594_/Q _12728_/S vssd1 vssd1 vccd1 vccd1 _07046_/X sky130_fd_sc_hd__mux2_1
XFILLER_134_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_208_clk clkbuf_5_16_0_clk/X vssd1 vssd1 vccd1 vccd1 _14420_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_88_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_1032 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08997_ _14233_/Q _14265_/Q _14297_/Q _14329_/Q _09005_/S _09523_/A1 vssd1 vssd1
+ vccd1 vccd1 _08997_/X sky130_fd_sc_hd__mux4_1
XFILLER_87_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07948_ _07961_/C _07947_/Y _07964_/A vssd1 vssd1 vccd1 vccd1 _07948_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_75_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07879_ _07881_/B _07878_/X _07874_/A vssd1 vssd1 vccd1 vccd1 _07879_/X sky130_fd_sc_hd__a21bo_1
XFILLER_28_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09618_ _13992_/Q _13340_/A0 _09628_/S vssd1 vssd1 vccd1 vccd1 _13992_/D sky130_fd_sc_hd__mux2_1
XFILLER_83_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_399 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10890_ _14922_/Q _15538_/Q _12904_/S vssd1 vssd1 vccd1 vccd1 _14922_/D sky130_fd_sc_hd__mux2_1
XFILLER_19_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09549_ _13906_/Q _08494_/Y _08512_/B _14421_/Q _13123_/A vssd1 vssd1 vccd1 vccd1
+ _09549_/X sky130_fd_sc_hd__a221o_1
XFILLER_12_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_1014 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12560_ _06670_/A _12557_/X _06671_/A vssd1 vssd1 vccd1 vccd1 _12560_/X sky130_fd_sc_hd__o21a_1
XFILLER_140_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11511_ _11536_/A _11511_/B vssd1 vssd1 vccd1 vccd1 _11512_/B sky130_fd_sc_hd__xor2_1
X_12491_ _08453_/A _12488_/X _08451_/A vssd1 vssd1 vccd1 vccd1 _12491_/X sky130_fd_sc_hd__o21a_1
XFILLER_12_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14230_ _14537_/CLK _14230_/D vssd1 vssd1 vccd1 vccd1 _14230_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11442_ _11420_/A _11430_/X _11441_/A vssd1 vssd1 vccd1 vccd1 _11442_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_137_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14161_ _15672_/CLK _14161_/D vssd1 vssd1 vccd1 vccd1 _14161_/Q sky130_fd_sc_hd__dfxtp_1
X_11373_ _11423_/A vssd1 vssd1 vccd1 vccd1 _11377_/A sky130_fd_sc_hd__inv_2
XFILLER_165_794 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13112_ _13035_/X _13118_/A2 _13114_/B1 _07496_/X vssd1 vssd1 vccd1 vccd1 _13112_/X
+ sky130_fd_sc_hd__a22o_1
X_10324_ _14896_/Q _14709_/Q _10344_/S vssd1 vssd1 vccd1 vccd1 _14709_/D sky130_fd_sc_hd__mux2_1
XFILLER_30_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14092_ _14405_/CLK _14092_/D vssd1 vssd1 vccd1 vccd1 _14092_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10255_ _14640_/Q _14793_/Q _10715_/S vssd1 vssd1 vccd1 vccd1 _14640_/D sky130_fd_sc_hd__mux2_1
XTAP_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13043_ _13125_/B _08538_/A _12934_/Y vssd1 vssd1 vccd1 vccd1 _13043_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_124_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10186_ _11872_/A1 _14570_/Q _10197_/S vssd1 vssd1 vccd1 vccd1 _14570_/D sky130_fd_sc_hd__mux2_1
XFILLER_61_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14994_ _15046_/CLK _14994_/D vssd1 vssd1 vccd1 vccd1 _14994_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout290 _07488_/X vssd1 vssd1 vccd1 vccd1 _13347_/A0 sky130_fd_sc_hd__buf_6
XFILLER_93_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13945_ _15178_/CLK _13945_/D vssd1 vssd1 vccd1 vccd1 _13945_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_163 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13876_ _15077_/CLK _13876_/D vssd1 vssd1 vccd1 vccd1 _13876_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15615_ _15615_/CLK _15615_/D vssd1 vssd1 vccd1 vccd1 _15615_/Q sky130_fd_sc_hd__dfxtp_4
X_12827_ _15366_/Q _12827_/B vssd1 vssd1 vccd1 vccd1 _12828_/B sky130_fd_sc_hd__xor2_1
XFILLER_90_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15546_ _15552_/CLK _15546_/D vssd1 vssd1 vccd1 vccd1 _15546_/Q sky130_fd_sc_hd__dfxtp_1
X_12758_ _13433_/Q _12757_/X _12764_/S vssd1 vssd1 vccd1 vccd1 _12758_/X sky130_fd_sc_hd__mux2_1
XTAP_1281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11709_ _14716_/Q _11743_/C _14714_/Q vssd1 vssd1 vccd1 vccd1 _11851_/B sky130_fd_sc_hd__or3b_4
X_15477_ _15501_/CLK _15477_/D vssd1 vssd1 vccd1 vccd1 _15477_/Q sky130_fd_sc_hd__dfxtp_1
X_12689_ _12701_/C _12689_/B vssd1 vssd1 vccd1 vccd1 _12689_/Y sky130_fd_sc_hd__nor2_1
XFILLER_30_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14428_ _14462_/CLK _14428_/D vssd1 vssd1 vccd1 vccd1 _14428_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14359_ _14525_/CLK _14359_/D vssd1 vssd1 vccd1 vccd1 _14359_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08920_ _09382_/A _08920_/B _08920_/C vssd1 vssd1 vccd1 vccd1 _08920_/X sky130_fd_sc_hd__and3_1
XFILLER_157_1079 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08851_ _13874_/Q _11883_/A1 _08851_/S vssd1 vssd1 vccd1 vccd1 _13874_/D sky130_fd_sc_hd__mux2_1
XFILLER_85_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07802_ _13512_/Q _13511_/Q _07802_/C _07802_/D vssd1 vssd1 vccd1 vccd1 _07813_/D
+ sky130_fd_sc_hd__and4_2
XFILLER_69_288 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08782_ _13810_/Q _10892_/B _08779_/X vssd1 vssd1 vccd1 vccd1 _13810_/D sky130_fd_sc_hd__a21bo_1
XFILLER_66_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07733_ _07730_/Y _07739_/C _07750_/A vssd1 vssd1 vccd1 vccd1 _07733_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_38_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07664_ _13477_/Q _07665_/C _13478_/Q vssd1 vssd1 vccd1 vccd1 _07664_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_111_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09403_ _14091_/Q _08494_/Y _09403_/B1 _14059_/Q _09391_/A vssd1 vssd1 vccd1 vccd1
+ _09403_/X sky130_fd_sc_hd__a221o_1
X_07595_ _07595_/A _07595_/B vssd1 vssd1 vccd1 vccd1 _07603_/D sky130_fd_sc_hd__nor2_1
X_09334_ _13960_/Q _13702_/Q _09342_/S vssd1 vssd1 vccd1 vccd1 _09334_/X sky130_fd_sc_hd__mux2_1
XFILLER_178_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09265_ _13861_/Q _14214_/Q _09557_/S vssd1 vssd1 vccd1 vccd1 _09265_/X sky130_fd_sc_hd__mux2_1
X_08216_ _13707_/Q _13104_/B2 _08216_/S vssd1 vssd1 vccd1 vccd1 _13707_/D sky130_fd_sc_hd__mux2_1
X_09196_ _09130_/A _09189_/X _09192_/X _09450_/B1 vssd1 vssd1 vccd1 vccd1 _09196_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_5_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_772 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_603 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08147_ _08093_/B _08145_/X _08146_/Y _08121_/X vssd1 vssd1 vccd1 vccd1 _08147_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_107_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08078_ _08078_/A _08078_/B _08083_/A vssd1 vssd1 vccd1 vccd1 _08078_/X sky130_fd_sc_hd__or3b_1
XFILLER_150_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07029_ _07028_/X _14742_/Q _07098_/S vssd1 vssd1 vccd1 vccd1 _13588_/D sky130_fd_sc_hd__mux2_1
XFILLER_96_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10040_ _14397_/Q _13326_/A0 _10059_/S vssd1 vssd1 vccd1 vccd1 _14397_/D sky130_fd_sc_hd__mux2_1
XFILLER_96_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_406 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11991_ _14007_/Q _13975_/Q _11993_/S vssd1 vssd1 vccd1 vccd1 _11992_/B sky130_fd_sc_hd__mux2_1
XFILLER_28_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13730_ _15530_/CLK _13730_/D vssd1 vssd1 vccd1 vccd1 _13730_/Q sky130_fd_sc_hd__dfxtp_2
X_10942_ _11600_/A _10948_/B vssd1 vssd1 vccd1 vccd1 _10942_/Y sky130_fd_sc_hd__nand2_1
XFILLER_43_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13661_ _14774_/CLK _13661_/D vssd1 vssd1 vccd1 vccd1 _13661_/Q sky130_fd_sc_hd__dfxtp_1
X_10873_ _13733_/Q _14905_/Q _10877_/S vssd1 vssd1 vccd1 vccd1 _14905_/D sky130_fd_sc_hd__mux2_1
XFILLER_43_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15400_ _15617_/CLK _15400_/D vssd1 vssd1 vccd1 vccd1 _15400_/Q sky130_fd_sc_hd__dfxtp_2
XPHY_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12612_ _14034_/Q _14002_/Q _12612_/S vssd1 vssd1 vccd1 vccd1 _12613_/B sky130_fd_sc_hd__mux2_1
XPHY_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13592_ _15453_/CLK _13592_/D vssd1 vssd1 vccd1 vccd1 _13592_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15331_ _15331_/CLK _15331_/D vssd1 vssd1 vccd1 vccd1 _15331_/Q sky130_fd_sc_hd__dfxtp_2
XPHY_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12543_ _14031_/Q _13999_/Q _12543_/S vssd1 vssd1 vccd1 vccd1 _12544_/B sky130_fd_sc_hd__mux2_1
XFILLER_61_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15262_ _15544_/CLK _15262_/D vssd1 vssd1 vccd1 vccd1 _15262_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_185_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12474_ _14028_/Q _13996_/Q _12476_/S vssd1 vssd1 vccd1 vccd1 _12475_/B sky130_fd_sc_hd__mux2_1
XFILLER_8_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14213_ _14373_/CLK _14213_/D vssd1 vssd1 vccd1 vccd1 _14213_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_184_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11425_ _11460_/D _11425_/B vssd1 vssd1 vccd1 vccd1 _11425_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_144_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15193_ _15304_/CLK _15193_/D vssd1 vssd1 vccd1 vccd1 _15193_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_7 _08903_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14144_ _15662_/CLK _14144_/D vssd1 vssd1 vccd1 vccd1 _14144_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11356_ _13251_/A _11356_/B _11356_/C vssd1 vssd1 vccd1 vccd1 _11357_/C sky130_fd_sc_hd__or3_1
XFILLER_125_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10307_ _14692_/Q _14877_/Q _10710_/S vssd1 vssd1 vccd1 vccd1 _14692_/D sky130_fd_sc_hd__mux2_1
XFILLER_125_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14075_ _15657_/CLK _14075_/D vssd1 vssd1 vccd1 vccd1 _14075_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_125_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11287_ _11318_/S _11305_/B _11305_/C vssd1 vssd1 vccd1 vccd1 _11287_/X sky130_fd_sc_hd__and3_1
XFILLER_112_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13026_ _10714_/X _14889_/Q _13029_/S vssd1 vssd1 vccd1 vccd1 _13026_/X sky130_fd_sc_hd__mux2_4
XFILLER_140_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10238_ _14623_/Q _14776_/Q _10630_/S vssd1 vssd1 vccd1 vccd1 _14623_/D sky130_fd_sc_hd__mux2_1
XFILLER_67_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10169_ _13322_/A0 _14553_/Q _10192_/S vssd1 vssd1 vccd1 vccd1 _14553_/D sky130_fd_sc_hd__mux2_1
XFILLER_86_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14977_ _15577_/CLK _14977_/D vssd1 vssd1 vccd1 vccd1 _14977_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_94_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13928_ _15544_/CLK _13928_/D vssd1 vssd1 vccd1 vccd1 _13928_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_179_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13859_ _15108_/CLK _13859_/D vssd1 vssd1 vccd1 vccd1 _13859_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_604 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07380_ _14735_/Q _07379_/X _07500_/S vssd1 vssd1 vccd1 vccd1 _07380_/X sky130_fd_sc_hd__mux2_8
XFILLER_15_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15529_ _15529_/CLK _15529_/D vssd1 vssd1 vccd1 vccd1 _15529_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_187_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09050_ _15115_/Q _15083_/Q _15656_/Q _13390_/Q _09407_/S _09406_/S1 vssd1 vssd1
+ vccd1 vccd1 _09050_/X sky130_fd_sc_hd__mux4_1
XFILLER_159_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08001_ _08003_/B _08000_/X _08022_/B vssd1 vssd1 vccd1 vccd1 _08001_/X sky130_fd_sc_hd__a21bo_1
XFILLER_116_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09952_ _11872_/A1 _14312_/Q _09963_/S vssd1 vssd1 vccd1 vccd1 _14312_/D sky130_fd_sc_hd__mux2_1
XFILLER_116_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08903_ _06676_/A _08892_/X _08901_/X _08902_/X vssd1 vssd1 vccd1 vccd1 _08903_/X
+ sky130_fd_sc_hd__o22a_2
XFILLER_98_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09883_ _11761_/A0 _14245_/Q _09897_/S vssd1 vssd1 vccd1 vccd1 _14245_/D sky130_fd_sc_hd__mux2_1
XFILLER_140_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08834_ _13857_/Q _13080_/B2 _08846_/S vssd1 vssd1 vccd1 vccd1 _13857_/D sky130_fd_sc_hd__mux2_1
XTAP_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08765_ _08765_/A _14595_/Q _14587_/Q _08765_/D vssd1 vssd1 vccd1 vccd1 _08765_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_73_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07716_ _13492_/Q _13491_/Q _13490_/Q _13489_/Q vssd1 vssd1 vccd1 vccd1 _07732_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_54_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08696_ _13548_/Q _08747_/A2 _08747_/B1 _13484_/Q vssd1 vssd1 vccd1 vccd1 _08696_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_25_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07647_ _13474_/Q _13473_/Q _07647_/C vssd1 vssd1 vccd1 vccd1 _07650_/B sky130_fd_sc_hd__and3_2
XFILLER_25_155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_306 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07578_ _14744_/Q _07629_/A _07577_/Y _07949_/C1 vssd1 vssd1 vccd1 vccd1 _13455_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_90_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09317_ _09554_/A _09317_/B _09317_/C vssd1 vssd1 vccd1 vccd1 _09317_/X sky130_fd_sc_hd__and3_1
XFILLER_40_158 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09248_ _09550_/A1 _09246_/X _09247_/X vssd1 vssd1 vccd1 vccd1 _09252_/B sky130_fd_sc_hd__a21o_1
XFILLER_108_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_4_10_0_clk clkbuf_3_5_0_clk/X vssd1 vssd1 vccd1 vccd1 clkbuf_5_21_0_clk/A
+ sky130_fd_sc_hd__clkbuf_8
X_09179_ _13920_/Q _09178_/X _12481_/A vssd1 vssd1 vccd1 vccd1 _13920_/D sky130_fd_sc_hd__mux2_1
XFILLER_108_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_99 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11210_ _10555_/B _14999_/Q _11237_/S vssd1 vssd1 vccd1 vccd1 _14999_/D sky130_fd_sc_hd__mux2_1
X_12190_ _15286_/Q _15254_/Q _15222_/Q _15153_/Q _12489_/S0 _12465_/S1 vssd1 vssd1
+ vccd1 vccd1 _12191_/B sky130_fd_sc_hd__mux4_1
XFILLER_150_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11141_ _11344_/A _11191_/B vssd1 vssd1 vccd1 vccd1 _11141_/Y sky130_fd_sc_hd__nand2_1
XFILLER_123_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput44 _07180_/X vssd1 vssd1 vccd1 vccd1 ext_address[18] sky130_fd_sc_hd__clkbuf_2
Xoutput55 _07191_/X vssd1 vssd1 vccd1 vccd1 ext_address[29] sky130_fd_sc_hd__clkbuf_2
Xoutput66 _06865_/B vssd1 vssd1 vccd1 vccd1 ext_instruction sky130_fd_sc_hd__clkbuf_2
Xoutput77 _07139_/X vssd1 vssd1 vccd1 vccd1 ext_write_data[19] sky130_fd_sc_hd__clkbuf_2
X_11072_ _11380_/A _11071_/X _11202_/A vssd1 vssd1 vccd1 vccd1 _11072_/Y sky130_fd_sc_hd__o21ai_1
Xoutput88 _07159_/X vssd1 vssd1 vccd1 vccd1 ext_write_data[29] sky130_fd_sc_hd__clkbuf_2
Xoutput99 _07101_/X vssd1 vssd1 vccd1 vccd1 ext_write_strobe[0] sky130_fd_sc_hd__clkbuf_2
XFILLER_163_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10023_ _11877_/A1 _14381_/Q _10028_/S vssd1 vssd1 vccd1 vccd1 _14381_/D sky130_fd_sc_hd__mux2_1
X_14900_ _15536_/CLK _14900_/D vssd1 vssd1 vccd1 vccd1 _14900_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_89_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14831_ _15536_/CLK _14831_/D vssd1 vssd1 vccd1 vccd1 _14831_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_56_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14762_ _15647_/CLK _14762_/D vssd1 vssd1 vccd1 vccd1 _14762_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_3964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11974_ _12273_/A1 _11973_/X _11972_/X _12503_/C1 vssd1 vssd1 vccd1 vccd1 _11975_/C
+ sky130_fd_sc_hd__a211o_1
XTAP_3975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13713_ _15584_/CLK _13713_/D vssd1 vssd1 vccd1 vccd1 _13713_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10925_ _11500_/A _10929_/B vssd1 vssd1 vccd1 vccd1 _10925_/X sky130_fd_sc_hd__and2b_1
X_14693_ _15608_/CLK _14693_/D vssd1 vssd1 vccd1 vccd1 _14693_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13644_ _15372_/CLK _13644_/D vssd1 vssd1 vccd1 vccd1 _13644_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10856_ _14888_/Q _13780_/Q _12878_/S vssd1 vssd1 vccd1 vccd1 _14888_/D sky130_fd_sc_hd__mux2_1
XFILLER_188_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13575_ _14493_/CLK _13575_/D vssd1 vssd1 vccd1 vccd1 _13575_/Q sky130_fd_sc_hd__dfxtp_2
X_10787_ _14819_/Q _15451_/Q _12929_/S vssd1 vssd1 vccd1 vccd1 _14819_/D sky130_fd_sc_hd__mux2_1
XFILLER_13_884 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15314_ _15656_/CLK _15314_/D vssd1 vssd1 vccd1 vccd1 _15314_/Q sky130_fd_sc_hd__dfxtp_2
XPHY_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12526_ _12618_/A1 _12525_/X _12524_/X _12618_/C1 vssd1 vssd1 vccd1 vccd1 _12527_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_184_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15245_ _15277_/CLK _15245_/D vssd1 vssd1 vccd1 vccd1 _15245_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12457_ _12503_/A1 _12456_/X _12455_/X _12503_/C1 vssd1 vssd1 vccd1 vccd1 _12458_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_126_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11408_ _13178_/B _11409_/B vssd1 vssd1 vccd1 vccd1 _11421_/B sky130_fd_sc_hd__nor2_1
X_15176_ _15176_/CLK _15176_/D vssd1 vssd1 vccd1 vccd1 _15176_/Q sky130_fd_sc_hd__dfxtp_1
X_12388_ _12618_/A1 _12387_/X _12386_/X _12618_/C1 vssd1 vssd1 vccd1 vccd1 _12389_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_153_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_1103 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14127_ _15094_/CLK _14127_/D vssd1 vssd1 vccd1 vccd1 _14127_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11339_ _11283_/A _11282_/X _11338_/X vssd1 vssd1 vccd1 vccd1 _11339_/X sky130_fd_sc_hd__o21a_1
XFILLER_98_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14058_ _15328_/CLK _14058_/D vssd1 vssd1 vccd1 vccd1 _14058_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13009_ _07460_/X _13039_/A2 _13008_/X _12944_/A vssd1 vssd1 vccd1 vccd1 _13009_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_67_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06880_ _14514_/Q _06873_/B _14513_/Q _06698_/Y _06871_/B vssd1 vssd1 vccd1 vccd1
+ _06880_/X sky130_fd_sc_hd__a221o_1
XFILLER_39_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08550_ _13609_/Q _08749_/A2 _08750_/B1 _13641_/Q vssd1 vssd1 vccd1 vccd1 _08550_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_82_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07501_ _13350_/A0 _13414_/Q _07501_/S vssd1 vssd1 vccd1 vccd1 _13414_/D sky130_fd_sc_hd__mux2_1
XFILLER_63_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08481_ _09405_/A _08487_/B vssd1 vssd1 vccd1 vccd1 _08481_/X sky130_fd_sc_hd__and2_1
XFILLER_62_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07432_ _14748_/Q _07431_/X _07480_/S vssd1 vssd1 vccd1 vccd1 _07432_/X sky130_fd_sc_hd__mux2_8
XFILLER_23_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07363_ _07363_/A _07363_/B _07363_/C _07363_/D vssd1 vssd1 vccd1 vccd1 _07363_/X
+ sky130_fd_sc_hd__or4_1
X_09102_ _14464_/Q _14432_/Q _13853_/Q _14206_/Q _09438_/S0 _09448_/S1 vssd1 vssd1
+ vccd1 vccd1 _09102_/X sky130_fd_sc_hd__mux4_2
XFILLER_149_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07294_ _07294_/A vssd1 vssd1 vccd1 vccd1 _07294_/Y sky130_fd_sc_hd__inv_2
XFILLER_30_180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_686 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09033_ _08519_/B _09031_/X _09032_/X _08668_/D vssd1 vssd1 vccd1 vccd1 _09033_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_108_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_712 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_892 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09935_ _13322_/A0 _14295_/Q _09958_/S vssd1 vssd1 vccd1 vccd1 _14295_/D sky130_fd_sc_hd__mux2_1
XFILLER_131_244 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09866_ _11852_/A1 _14228_/Q _09892_/S vssd1 vssd1 vccd1 vccd1 _14228_/D sky130_fd_sc_hd__mux2_1
XTAP_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08817_ _14714_/Q _08817_/B vssd1 vssd1 vccd1 vccd1 _08817_/Y sky130_fd_sc_hd__nand2_2
XFILLER_133_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09797_ _14163_/Q _13319_/A0 _09823_/S vssd1 vssd1 vccd1 vccd1 _14163_/D sky130_fd_sc_hd__mux2_1
XFILLER_58_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08748_ _15368_/Q _08748_/A2 _08748_/B1 _14486_/Q vssd1 vssd1 vccd1 vccd1 _08748_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_2515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08679_ _13590_/Q _08691_/A2 _08693_/B1 _13622_/Q vssd1 vssd1 vccd1 vccd1 _08679_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_26_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10710_ _14760_/Q _10709_/X _10710_/S vssd1 vssd1 vccd1 vccd1 _14760_/D sky130_fd_sc_hd__mux2_1
XFILLER_14_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11690_ _13332_/A0 _15121_/Q _11703_/S vssd1 vssd1 vccd1 vccd1 _15121_/D sky130_fd_sc_hd__mux2_1
XTAP_1869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_406 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10641_ _15566_/Q _10706_/B vssd1 vssd1 vccd1 vccd1 _10641_/X sky130_fd_sc_hd__and2_1
XFILLER_13_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13360_ _14463_/Q vssd1 vssd1 vccd1 vccd1 _14463_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_166_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10572_ _10581_/B _10570_/X _10571_/X _10581_/A vssd1 vssd1 vccd1 vccd1 _10572_/X
+ sky130_fd_sc_hd__o211a_1
X_12311_ _13893_/Q _14408_/Q _12614_/S vssd1 vssd1 vccd1 vccd1 _12311_/X sky130_fd_sc_hd__mux2_1
XFILLER_177_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_539 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13291_ _12659_/Y _15623_/Q _13291_/S vssd1 vssd1 vccd1 vccd1 _15623_/D sky130_fd_sc_hd__mux2_1
XFILLER_182_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15030_ _15042_/CLK _15030_/D vssd1 vssd1 vccd1 vccd1 _15030_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_177_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12242_ _13890_/Q _14405_/Q _12246_/S vssd1 vssd1 vccd1 vccd1 _12242_/X sky130_fd_sc_hd__mux2_1
XFILLER_5_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12173_ _13887_/Q _14402_/Q _12246_/S vssd1 vssd1 vccd1 vccd1 _12173_/X sky130_fd_sc_hd__mux2_1
XFILLER_150_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11124_ _11074_/X _11084_/X _11297_/S vssd1 vssd1 vccd1 vccd1 _11124_/X sky130_fd_sc_hd__mux2_1
XFILLER_174_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_1000 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_91 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11055_ _11129_/B vssd1 vssd1 vccd1 vccd1 _11055_/Y sky130_fd_sc_hd__inv_2
XFILLER_67_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10006_ _11860_/A1 _14364_/Q _10028_/S vssd1 vssd1 vccd1 vccd1 _14364_/D sky130_fd_sc_hd__mux2_1
XFILLER_92_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14814_ _15446_/CLK _14814_/D vssd1 vssd1 vccd1 vccd1 _14814_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14745_ _15592_/CLK _14745_/D vssd1 vssd1 vccd1 vccd1 _14745_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_3794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11957_ _15111_/Q _15079_/Q _15652_/Q _13386_/Q _12453_/S _12061_/A vssd1 vssd1 vccd1
+ vccd1 _11957_/X sky130_fd_sc_hd__mux4_1
XFILLER_44_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10908_ _13178_/B _13177_/A vssd1 vssd1 vccd1 vccd1 _10908_/Y sky130_fd_sc_hd__nand2_1
XFILLER_32_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14676_ _15647_/CLK _14676_/D vssd1 vssd1 vccd1 vccd1 _14676_/Q sky130_fd_sc_hd__dfxtp_1
X_11888_ _15108_/Q _15076_/Q _15649_/Q _13383_/Q _12154_/S _11992_/A vssd1 vssd1 vccd1
+ vccd1 _11888_/X sky130_fd_sc_hd__mux4_1
XFILLER_149_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13627_ _13627_/CLK _13627_/D vssd1 vssd1 vccd1 vccd1 _13627_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10839_ _14871_/Q _13797_/Q _12927_/S vssd1 vssd1 vccd1 vccd1 _14871_/D sky130_fd_sc_hd__mux2_1
XFILLER_34_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13558_ _15386_/CLK _13558_/D vssd1 vssd1 vccd1 vccd1 _13558_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_158_675 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_1078 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12509_ _15135_/Q _15103_/Q _15676_/Q _13410_/Q _12522_/S _12521_/A vssd1 vssd1 vccd1
+ vccd1 _12509_/X sky130_fd_sc_hd__mux4_1
X_13489_ _15383_/CLK _13489_/D vssd1 vssd1 vccd1 vccd1 _13489_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_145_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_172_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15228_ _15275_/CLK _15228_/D vssd1 vssd1 vccd1 vccd1 _15228_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_126_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15159_ _15275_/CLK _15159_/D vssd1 vssd1 vccd1 vccd1 _15159_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout108 _13288_/S vssd1 vssd1 vccd1 vccd1 _13282_/S sky130_fd_sc_hd__buf_8
X_07981_ _13561_/Q _07981_/B vssd1 vssd1 vccd1 vccd1 _07981_/X sky130_fd_sc_hd__xor2_1
Xfanout119 _13051_/X vssd1 vssd1 vccd1 vccd1 _13104_/B1 sky130_fd_sc_hd__clkbuf_16
XFILLER_86_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09720_ _13342_/A0 _14090_/Q _09728_/S vssd1 vssd1 vccd1 vccd1 _14090_/D sky130_fd_sc_hd__mux2_1
X_06932_ _06923_/X _06926_/X _06929_/X _06931_/Y vssd1 vssd1 vccd1 vccd1 _06932_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_101_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09651_ _14024_/Q _13340_/A0 _09661_/S vssd1 vssd1 vccd1 vccd1 _14024_/D sky130_fd_sc_hd__mux2_1
XFILLER_110_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06863_ _12828_/A _06863_/B vssd1 vssd1 vccd1 vccd1 _12622_/A sky130_fd_sc_hd__or2_4
X_08602_ _15389_/Q _08748_/A2 _08736_/A2 _13434_/Q vssd1 vssd1 vccd1 vccd1 _08602_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_82_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09582_ _13958_/Q _13338_/A0 _09594_/S vssd1 vssd1 vccd1 vccd1 _13958_/D sky130_fd_sc_hd__mux2_1
X_06794_ _14596_/Q _14595_/Q vssd1 vssd1 vccd1 vccd1 _06796_/B sky130_fd_sc_hd__nor2_1
X_08533_ _13508_/Q _08747_/B1 _08750_/B1 _13643_/Q vssd1 vssd1 vccd1 vccd1 _08533_/X
+ sky130_fd_sc_hd__a22o_1
X_08464_ _14595_/Q _12900_/S _08773_/B _08463_/X vssd1 vssd1 vccd1 vccd1 _13762_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_24_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07415_ _13659_/Q _07483_/A2 _07483_/B1 _14687_/Q _07414_/X vssd1 vssd1 vccd1 vccd1
+ _07415_/X sky130_fd_sc_hd__a221o_1
XFILLER_50_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08395_ _13729_/Q _13140_/S _08394_/X hold8/X vssd1 vssd1 vccd1 vccd1 _13729_/D sky130_fd_sc_hd__a22o_1
XFILLER_148_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07346_ _07312_/X _07314_/Y _07319_/X _07321_/Y vssd1 vssd1 vccd1 vccd1 _07360_/D
+ sky130_fd_sc_hd__o22ai_2
XFILLER_148_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07277_ _15321_/Q _15477_/Q _07340_/S vssd1 vssd1 vccd1 vccd1 _07278_/B sky130_fd_sc_hd__mux2_4
XFILLER_164_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09016_ _14362_/Q _15178_/Q _13817_/Q _14556_/Q _09521_/S _09523_/A1 vssd1 vssd1
+ vccd1 vccd1 _09017_/B sky130_fd_sc_hd__mux4_1
XFILLER_128_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout620 _12545_/S vssd1 vssd1 vccd1 vccd1 _12541_/S sky130_fd_sc_hd__buf_12
Xfanout631 _13242_/A vssd1 vssd1 vccd1 vccd1 _13251_/A sky130_fd_sc_hd__buf_12
X_09918_ _13338_/A0 _14279_/Q _09930_/S vssd1 vssd1 vccd1 vccd1 _14279_/D sky130_fd_sc_hd__mux2_1
Xfanout642 fanout647/X vssd1 vssd1 vccd1 vccd1 _08012_/C1 sky130_fd_sc_hd__clkbuf_8
X_09849_ _14213_/Q _11761_/A0 _09863_/S vssd1 vssd1 vccd1 vccd1 _14213_/D sky130_fd_sc_hd__mux2_1
XFILLER_74_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12860_ _14754_/Q _15388_/Q _12866_/S vssd1 vssd1 vccd1 vccd1 _15388_/D sky130_fd_sc_hd__mux2_1
XFILLER_37_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11811_ _15234_/Q _11877_/A1 _11816_/S vssd1 vssd1 vccd1 vccd1 _15234_/D sky130_fd_sc_hd__mux2_1
XTAP_2334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12791_ _13309_/B _13309_/C _12792_/B vssd1 vssd1 vccd1 vccd1 _12791_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_26_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14530_ _14530_/CLK _14530_/D vssd1 vssd1 vccd1 vccd1 _14530_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11742_ _15171_/Q _13350_/A0 _11742_/S vssd1 vssd1 vccd1 vccd1 _15171_/D sky130_fd_sc_hd__mux2_1
XTAP_2389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_1007 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14461_ _15649_/CLK _14461_/D vssd1 vssd1 vccd1 vccd1 _14461_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11673_ _11881_/A1 _15105_/Q _11675_/S vssd1 vssd1 vccd1 vccd1 _15105_/D sky130_fd_sc_hd__mux2_1
XTAP_1699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13412_ _15678_/CLK _13412_/D vssd1 vssd1 vccd1 vccd1 _13412_/Q sky130_fd_sc_hd__dfxtp_1
X_10624_ _15052_/Q _10714_/A2 _10621_/X _10623_/X vssd1 vssd1 vccd1 vccd1 _10624_/X
+ sky130_fd_sc_hd__o22a_4
X_14392_ _15211_/CLK _14392_/D vssd1 vssd1 vccd1 vccd1 _14392_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_167_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13343_ _13343_/A0 _15673_/Q _13345_/S vssd1 vssd1 vccd1 vccd1 _15673_/D sky130_fd_sc_hd__mux2_1
X_10555_ _10555_/A _10555_/B _10555_/C _10555_/D vssd1 vssd1 vccd1 vccd1 _10556_/D
+ sky130_fd_sc_hd__or4_1
XFILLER_128_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13274_ _15358_/Q _15605_/Q _13309_/A vssd1 vssd1 vccd1 vccd1 _15605_/D sky130_fd_sc_hd__mux2_1
X_10486_ _07237_/A _08225_/Y _10485_/X vssd1 vssd1 vccd1 vccd1 _11561_/A sky130_fd_sc_hd__a21o_4
XFILLER_142_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15013_ _15014_/CLK _15013_/D vssd1 vssd1 vccd1 vccd1 _15013_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12225_ _12218_/X _12220_/X _12222_/X _12224_/X _12501_/C1 vssd1 vssd1 vccd1 vccd1
+ _12225_/X sky130_fd_sc_hd__o221a_1
XFILLER_64_1016 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12156_ _12149_/X _12151_/X _12153_/X _12155_/X _12455_/C1 vssd1 vssd1 vccd1 vccd1
+ _12156_/X sky130_fd_sc_hd__o221a_1
XFILLER_64_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11107_ _11021_/X _11039_/X _11115_/S vssd1 vssd1 vccd1 vccd1 _11107_/X sky130_fd_sc_hd__mux2_2
X_12087_ _12080_/X _12082_/X _12084_/X _12086_/X _12455_/C1 vssd1 vssd1 vccd1 vccd1
+ _12087_/X sky130_fd_sc_hd__o221a_1
XFILLER_1_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11038_ _11025_/A _13202_/B _11249_/B vssd1 vssd1 vccd1 vccd1 _11038_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_77_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12989_ _15476_/Q _10834_/S _13025_/B1 _12988_/X vssd1 vssd1 vccd1 vccd1 _15476_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_92_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14728_ _15552_/CLK _14728_/D vssd1 vssd1 vccd1 vccd1 _14728_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_162_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14659_ _15630_/CLK _14659_/D vssd1 vssd1 vccd1 vccd1 _14659_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_177_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_180_clk clkbuf_5_22_0_clk/X vssd1 vssd1 vccd1 vccd1 _14439_/CLK sky130_fd_sc_hd__clkbuf_16
X_07200_ _15335_/Q _15491_/Q _07335_/S vssd1 vssd1 vccd1 vccd1 _07201_/A sky130_fd_sc_hd__mux2_8
X_08180_ _13677_/Q _10730_/S _08155_/X _08179_/X vssd1 vssd1 vccd1 vccd1 _13677_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_186_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07131_ _07131_/A _07131_/B vssd1 vssd1 vccd1 vccd1 _07131_/X sky130_fd_sc_hd__and2_4
XFILLER_146_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07062_ _07061_/X _14753_/Q _07098_/S vssd1 vssd1 vccd1 vccd1 _13599_/D sky130_fd_sc_hd__mux2_1
XFILLER_145_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07964_ _07964_/A _07964_/B vssd1 vssd1 vccd1 vccd1 _07964_/Y sky130_fd_sc_hd__nand2_1
XFILLER_114_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09703_ _13325_/A0 _14073_/Q _09723_/S vssd1 vssd1 vccd1 vccd1 _14073_/D sky130_fd_sc_hd__mux2_1
X_06915_ _06714_/Y _13464_/Q _06717_/Y _13463_/Q vssd1 vssd1 vccd1 vccd1 _06922_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_96_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07895_ _07897_/B _07894_/X _07903_/A vssd1 vssd1 vccd1 vccd1 _07895_/X sky130_fd_sc_hd__a21bo_1
X_09634_ _14007_/Q _11681_/A0 _09660_/S vssd1 vssd1 vccd1 vccd1 _14007_/D sky130_fd_sc_hd__mux2_1
XFILLER_67_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06846_ _12618_/A1 _14908_/Q _14909_/Q _06672_/Y _06845_/Y vssd1 vssd1 vccd1 vccd1
+ _06846_/X sky130_fd_sc_hd__o221a_1
XFILLER_167_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09565_ _13941_/Q _11854_/A1 _09594_/S vssd1 vssd1 vccd1 vccd1 _13941_/D sky130_fd_sc_hd__mux2_1
X_06777_ input33/X _06865_/B vssd1 vssd1 vccd1 vccd1 _06782_/A sky130_fd_sc_hd__or2_2
XFILLER_82_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08516_ _14612_/Q _14611_/Q _13133_/C _08536_/A vssd1 vssd1 vccd1 vccd1 _08528_/C
+ sky130_fd_sc_hd__o31a_1
X_09496_ _09532_/A _09496_/B vssd1 vssd1 vccd1 vccd1 _09496_/X sky130_fd_sc_hd__or2_1
XFILLER_169_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_404 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08447_ _08490_/A1 _08390_/C _08425_/X _10764_/S vssd1 vssd1 vccd1 vccd1 _08447_/X
+ sky130_fd_sc_hd__a211o_1
Xclkbuf_leaf_171_clk clkbuf_5_23_0_clk/X vssd1 vssd1 vccd1 vccd1 _15300_/CLK sky130_fd_sc_hd__clkbuf_16
X_08378_ _11347_/A _11290_/B vssd1 vssd1 vccd1 vccd1 _08378_/Y sky130_fd_sc_hd__nor2_1
XFILLER_17_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_143_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1095 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07329_ _07329_/A vssd1 vssd1 vccd1 vccd1 _07329_/Y sky130_fd_sc_hd__inv_2
XFILLER_136_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_976 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10340_ _14725_/Q _14918_/Q _10343_/S vssd1 vssd1 vccd1 vccd1 _14725_/D sky130_fd_sc_hd__mux2_1
XFILLER_137_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_935 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10271_ _14656_/Q _14809_/Q _10650_/S vssd1 vssd1 vccd1 vccd1 _14656_/D sky130_fd_sc_hd__mux2_1
XFILLER_117_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12010_ _13944_/Q _13686_/Q _12407_/S vssd1 vssd1 vccd1 vccd1 _12011_/B sky130_fd_sc_hd__mux2_1
XFILLER_3_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout450 _10244_/S vssd1 vssd1 vccd1 vccd1 _10710_/S sky130_fd_sc_hd__buf_12
Xfanout461 _13131_/A vssd1 vssd1 vccd1 vccd1 _09450_/B1 sky130_fd_sc_hd__buf_12
XFILLER_120_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout472 _12168_/A vssd1 vssd1 vccd1 vccd1 _12260_/A sky130_fd_sc_hd__buf_12
X_13961_ _15651_/CLK _13961_/D vssd1 vssd1 vccd1 vccd1 _13961_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout483 _06669_/Y vssd1 vssd1 vccd1 vccd1 _12477_/A1 sky130_fd_sc_hd__clkbuf_16
XFILLER_120_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout494 _15043_/Q vssd1 vssd1 vccd1 vccd1 _08094_/S sky130_fd_sc_hd__clkbuf_16
XFILLER_48_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12912_ _15440_/Q _15626_/Q _12918_/S vssd1 vssd1 vccd1 vccd1 _15440_/D sky130_fd_sc_hd__mux2_1
XFILLER_74_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_1036 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13892_ _15668_/CLK _13892_/D vssd1 vssd1 vccd1 vccd1 _13892_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_185_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15631_ _15632_/CLK _15631_/D vssd1 vssd1 vccd1 vccd1 _15631_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12843_ _14737_/Q _15371_/Q _12871_/S vssd1 vssd1 vccd1 vccd1 _15371_/D sky130_fd_sc_hd__mux2_1
XFILLER_74_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15562_ _15580_/CLK _15562_/D vssd1 vssd1 vccd1 vccd1 _15562_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12774_ _15358_/Q _12765_/B _12773_/X _12788_/C1 vssd1 vssd1 vccd1 vccd1 _15358_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_1430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14513_ _14513_/CLK _14513_/D vssd1 vssd1 vccd1 vccd1 _14513_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11725_ _15154_/Q _13080_/B2 _11741_/S vssd1 vssd1 vccd1 vccd1 _15154_/D sky130_fd_sc_hd__mux2_1
XFILLER_42_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15493_ _15525_/CLK _15493_/D vssd1 vssd1 vccd1 vccd1 _15493_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_162_clk clkbuf_5_19_0_clk/X vssd1 vssd1 vccd1 vccd1 _14225_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_1496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14444_ _15081_/CLK _14444_/D vssd1 vssd1 vccd1 vccd1 _14444_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11656_ _13331_/A0 _15088_/Q _11670_/S vssd1 vssd1 vccd1 vccd1 _15088_/D sky130_fd_sc_hd__mux2_1
XFILLER_156_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_95 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10607_ _15000_/Q _10569_/B _10602_/B _13719_/Q _10732_/C1 vssd1 vssd1 vccd1 vccd1
+ _10607_/X sky130_fd_sc_hd__a221o_1
XFILLER_156_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14375_ _15292_/CLK _14375_/D vssd1 vssd1 vccd1 vccd1 _14375_/Q sky130_fd_sc_hd__dfxtp_1
X_11587_ _11586_/A _11586_/B _11614_/S vssd1 vssd1 vccd1 vccd1 _11587_/X sky130_fd_sc_hd__o21ba_1
XFILLER_155_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_656 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13326_ _13326_/A0 _15656_/Q _13345_/S vssd1 vssd1 vccd1 vccd1 _15656_/D sky130_fd_sc_hd__mux2_1
X_10538_ _11536_/A _13208_/B _11536_/B _11500_/A vssd1 vssd1 vccd1 vccd1 _10538_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_143_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_496 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13257_ _15341_/Q _15588_/Q _13282_/S vssd1 vssd1 vccd1 vccd1 _15588_/D sky130_fd_sc_hd__mux2_1
X_10469_ _10532_/A _10469_/B vssd1 vssd1 vccd1 vccd1 _10470_/D sky130_fd_sc_hd__or2_1
XFILLER_89_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12208_ _14468_/Q _14436_/Q _13857_/Q _14210_/Q _08457_/A _12489_/S1 vssd1 vssd1
+ vccd1 vccd1 _12208_/X sky130_fd_sc_hd__mux4_1
XFILLER_130_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13188_ _15563_/Q _13241_/A2 _13186_/Y _13187_/X vssd1 vssd1 vccd1 vccd1 _15563_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_151_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12139_ _14465_/Q _14433_/Q _13854_/Q _14207_/Q _12472_/S _12465_/S1 vssd1 vssd1
+ vccd1 vccd1 _12139_/X sky130_fd_sc_hd__mux4_1
XFILLER_29_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06700_ _14512_/Q vssd1 vssd1 vccd1 vccd1 _06700_/Y sky130_fd_sc_hd__inv_2
XFILLER_49_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07680_ _07678_/Y _07687_/C _07676_/A vssd1 vssd1 vccd1 vccd1 _07680_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_64_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09350_ _15295_/Q _15263_/Q _15231_/Q _15162_/Q _09521_/S _09523_/A1 vssd1 vssd1
+ vccd1 vccd1 _09350_/X sky130_fd_sc_hd__mux4_1
XFILLER_64_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08301_ _11349_/B _11399_/A vssd1 vssd1 vccd1 vccd1 _11044_/B sky130_fd_sc_hd__and2_1
X_09281_ _12573_/A _09281_/B _09281_/C vssd1 vssd1 vccd1 vccd1 _09281_/X sky130_fd_sc_hd__and3_1
XFILLER_21_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_153_clk clkbuf_5_24_0_clk/X vssd1 vssd1 vccd1 vccd1 _15534_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_127_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08232_ _08232_/A _11344_/A vssd1 vssd1 vccd1 vccd1 _11309_/A sky130_fd_sc_hd__nor2_2
XFILLER_21_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08163_ _08185_/A _08163_/B vssd1 vssd1 vccd1 vccd1 _08163_/X sky130_fd_sc_hd__and2_1
XFILLER_109_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07114_ _14836_/Q _07115_/B _07157_/A vssd1 vssd1 vccd1 vccd1 _07114_/X sky130_fd_sc_hd__and3_4
XFILLER_180_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08094_ input1/X input31/X _08094_/S vssd1 vssd1 vccd1 vccd1 _08095_/B sky130_fd_sc_hd__mux2_1
X_07045_ _14627_/Q _14659_/Q _07078_/S vssd1 vssd1 vccd1 vccd1 _07045_/X sky130_fd_sc_hd__mux2_1
XFILLER_161_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_1044 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_383 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08996_ _08507_/A _08995_/X _08994_/X _09524_/A vssd1 vssd1 vccd1 vccd1 _08996_/X
+ sky130_fd_sc_hd__o211a_1
X_07947_ _13551_/Q _13550_/Q _07946_/D _13552_/Q vssd1 vssd1 vccd1 vccd1 _07947_/Y
+ sky130_fd_sc_hd__a31oi_1
XFILLER_102_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07878_ _13533_/Q _07884_/C _13534_/Q vssd1 vssd1 vccd1 vccd1 _07878_/X sky130_fd_sc_hd__a21o_1
XFILLER_141_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09617_ _13991_/Q _13092_/B2 _09628_/S vssd1 vssd1 vccd1 vccd1 _13991_/D sky130_fd_sc_hd__mux2_1
XFILLER_56_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06829_ _14709_/Q _08817_/B vssd1 vssd1 vccd1 vccd1 _07783_/A sky130_fd_sc_hd__nand2_4
XFILLER_56_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09548_ _13970_/Q _13712_/Q _09557_/S vssd1 vssd1 vccd1 vccd1 _09548_/X sky130_fd_sc_hd__mux2_1
XFILLER_169_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09479_ _14482_/Q _14450_/Q _13871_/Q _14224_/Q _09557_/S _09550_/A1 vssd1 vssd1
+ vccd1 vccd1 _09479_/X sky130_fd_sc_hd__mux4_1
XFILLER_54_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_144_clk clkbuf_5_28_0_clk/X vssd1 vssd1 vccd1 vccd1 _15374_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_169_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11510_ _11536_/B _11537_/A _13233_/A vssd1 vssd1 vccd1 vccd1 _11511_/B sky130_fd_sc_hd__a21o_1
XFILLER_12_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12490_ _12490_/A _12490_/B vssd1 vssd1 vccd1 vccd1 _12490_/X sky130_fd_sc_hd__or2_1
XFILLER_133_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11441_ _11441_/A _11441_/B vssd1 vssd1 vccd1 vccd1 _11441_/X sky130_fd_sc_hd__or2_1
XFILLER_138_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14160_ _15130_/CLK _14160_/D vssd1 vssd1 vccd1 vccd1 _14160_/Q sky130_fd_sc_hd__dfxtp_1
X_11372_ _11375_/B _11375_/C _13165_/B vssd1 vssd1 vccd1 vccd1 _11423_/A sky130_fd_sc_hd__a21bo_2
XFILLER_109_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_103 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13111_ _15523_/Q _10877_/S _13042_/A _13110_/X vssd1 vssd1 vccd1 vccd1 _15523_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_109_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10323_ _14708_/Q _14893_/Q _10735_/S vssd1 vssd1 vccd1 vccd1 _14708_/D sky130_fd_sc_hd__mux2_1
X_14091_ _14542_/CLK _14091_/D vssd1 vssd1 vccd1 vccd1 _14091_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13042_ _13042_/A vssd1 vssd1 vccd1 vccd1 _13042_/Y sky130_fd_sc_hd__inv_2
XFILLER_112_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10254_ _14639_/Q _14792_/Q _10695_/S vssd1 vssd1 vccd1 vccd1 _14639_/D sky130_fd_sc_hd__mux2_1
XFILLER_121_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10185_ _11838_/A1 _14569_/Q _10197_/S vssd1 vssd1 vccd1 vccd1 _14569_/D sky130_fd_sc_hd__mux2_1
XFILLER_59_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout280 _11309_/A vssd1 vssd1 vccd1 vccd1 _11351_/C1 sky130_fd_sc_hd__clkbuf_16
X_14993_ _15584_/CLK _14993_/D vssd1 vssd1 vccd1 vccd1 _14993_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout291 _07484_/X vssd1 vssd1 vccd1 vccd1 _13346_/A0 sky130_fd_sc_hd__buf_6
XFILLER_115_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_40 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_248 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13944_ _15081_/CLK _13944_/D vssd1 vssd1 vccd1 vccd1 _13944_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_911 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13875_ _15665_/CLK _13875_/D vssd1 vssd1 vccd1 vccd1 _13875_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_46_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15614_ _15647_/CLK _15614_/D vssd1 vssd1 vccd1 vccd1 _15614_/Q sky130_fd_sc_hd__dfxtp_1
X_12826_ _15366_/Q _12827_/B vssd1 vssd1 vccd1 vccd1 _12833_/B sky130_fd_sc_hd__nand2_1
XFILLER_188_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12757_ _13600_/Q _12756_/X _12785_/B vssd1 vssd1 vccd1 vccd1 _12757_/X sky130_fd_sc_hd__mux2_1
XTAP_1260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15545_ _15670_/CLK _15545_/D vssd1 vssd1 vccd1 vccd1 _15545_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_43_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_135_clk clkbuf_5_29_0_clk/X vssd1 vssd1 vccd1 vccd1 _13569_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_1282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11708_ _13350_/A0 _15139_/Q _11708_/S vssd1 vssd1 vccd1 vccd1 _15139_/D sky130_fd_sc_hd__mux2_1
X_15476_ _15501_/CLK _15476_/D vssd1 vssd1 vccd1 vccd1 _15476_/Q sky130_fd_sc_hd__dfxtp_1
X_12688_ _15347_/Q _12688_/B vssd1 vssd1 vccd1 vccd1 _12689_/B sky130_fd_sc_hd__nor2_1
X_14427_ _15211_/CLK _14427_/D vssd1 vssd1 vccd1 vccd1 _14427_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11639_ _11639_/A _11639_/B vssd1 vssd1 vccd1 vccd1 _11640_/B sky130_fd_sc_hd__xnor2_1
XFILLER_128_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14358_ _15275_/CLK _14358_/D vssd1 vssd1 vccd1 vccd1 _14358_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_772 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13309_ _13309_/A _13309_/B _13309_/C vssd1 vssd1 vccd1 vccd1 _13309_/X sky130_fd_sc_hd__or3_1
XFILLER_144_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14289_ _15526_/CLK _14289_/D vssd1 vssd1 vccd1 vccd1 _14289_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08850_ _13873_/Q _11816_/A1 _08851_/S vssd1 vssd1 vccd1 vccd1 _13873_/D sky130_fd_sc_hd__mux2_1
XFILLER_112_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07801_ _13514_/Q _13513_/Q vssd1 vssd1 vccd1 vccd1 _07802_/D sky130_fd_sc_hd__and2_1
XFILLER_69_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08781_ _13809_/Q _10892_/B _08775_/X vssd1 vssd1 vccd1 vccd1 _13809_/D sky130_fd_sc_hd__a21o_1
XFILLER_84_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_632 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07732_ _07732_/A _07732_/B _07732_/C vssd1 vssd1 vccd1 vccd1 _07739_/C sky130_fd_sc_hd__and3_2
XFILLER_38_665 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07663_ _14734_/Q _07777_/A _07662_/Y _08016_/C1 vssd1 vssd1 vccd1 vccd1 _13477_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_37_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09402_ _14027_/Q _13995_/Q _09407_/S vssd1 vssd1 vccd1 vccd1 _09402_/X sky130_fd_sc_hd__mux2_1
XFILLER_164_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07594_ _13459_/Q _07603_/C _13460_/Q vssd1 vssd1 vccd1 vccd1 _07594_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_53_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_5_31_0_clk clkbuf_5_31_0_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_5_31_0_clk/X
+ sky130_fd_sc_hd__clkbuf_8
X_09333_ _08510_/B _09329_/X _09332_/X _09328_/X vssd1 vssd1 vccd1 vccd1 _09346_/B
+ sky130_fd_sc_hd__a211o_1
Xclkbuf_leaf_126_clk clkbuf_5_31_0_clk/X vssd1 vssd1 vccd1 vccd1 _14506_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_179_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09264_ _14246_/Q _14278_/Q _14310_/Q _14342_/Q _09557_/S _09550_/A1 vssd1 vssd1
+ vccd1 vccd1 _09264_/X sky130_fd_sc_hd__mux4_1
XFILLER_139_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08215_ _13706_/Q _13344_/A0 _08216_/S vssd1 vssd1 vccd1 vccd1 _13706_/D sky130_fd_sc_hd__mux2_1
XFILLER_21_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09195_ _09449_/A1 _09193_/X _09194_/X _09449_/B2 vssd1 vssd1 vccd1 vccd1 _09195_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_146_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08146_ _08145_/S _06765_/Y _08151_/S vssd1 vssd1 vccd1 vccd1 _08146_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_107_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08077_ _15204_/Q _13645_/Q _08085_/S vssd1 vssd1 vccd1 vccd1 _08078_/A sky130_fd_sc_hd__mux2_1
XFILLER_106_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_1019 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07028_ _07027_/X _13588_/Q _12764_/S vssd1 vssd1 vccd1 vccd1 _07028_/X sky130_fd_sc_hd__mux2_1
XFILLER_121_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_565 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08979_ _13943_/Q _13685_/Q _09230_/S vssd1 vssd1 vccd1 vccd1 _08979_/X sky130_fd_sc_hd__mux2_1
XFILLER_88_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11990_ _12500_/A1 _11989_/X _12260_/A vssd1 vssd1 vccd1 vccd1 _11990_/X sky130_fd_sc_hd__a21o_1
XFILLER_91_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10941_ _14955_/Q _10940_/X _10944_/B vssd1 vssd1 vccd1 vccd1 _14955_/D sky130_fd_sc_hd__mux2_1
XFILLER_44_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13660_ _14703_/CLK _13660_/D vssd1 vssd1 vccd1 vccd1 _13660_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10872_ _13734_/Q _14904_/Q _13140_/S vssd1 vssd1 vccd1 vccd1 _14904_/D sky130_fd_sc_hd__mux2_1
XFILLER_72_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12611_ _12615_/A1 _12610_/X _12617_/S vssd1 vssd1 vccd1 vccd1 _12611_/X sky130_fd_sc_hd__a21o_1
X_13591_ _15453_/CLK _13591_/D vssd1 vssd1 vccd1 vccd1 _13591_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_117_clk _15447_/CLK vssd1 vssd1 vccd1 vccd1 _15378_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_71_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15330_ _15500_/CLK _15330_/D vssd1 vssd1 vccd1 vccd1 _15330_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12542_ _12592_/A1 _12541_/X _12536_/A vssd1 vssd1 vccd1 vccd1 _12542_/X sky130_fd_sc_hd__a21o_1
XPHY_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15261_ _15293_/CLK _15261_/D vssd1 vssd1 vccd1 vccd1 _15261_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_75 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12473_ _12477_/A1 _12472_/X _12490_/A vssd1 vssd1 vccd1 vccd1 _12473_/X sky130_fd_sc_hd__a21o_1
X_14212_ _15108_/CLK _14212_/D vssd1 vssd1 vccd1 vccd1 _14212_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11424_ _11404_/A _11423_/X _11422_/X vssd1 vssd1 vccd1 vccd1 _11425_/B sky130_fd_sc_hd__a21oi_4
X_15192_ _15192_/CLK _15192_/D vssd1 vssd1 vccd1 vccd1 _15192_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_8 _08970_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14143_ _14530_/CLK _14143_/D vssd1 vssd1 vccd1 vccd1 _14143_/Q sky130_fd_sc_hd__dfxtp_1
X_11355_ _10555_/C _07146_/S _11641_/S vssd1 vssd1 vccd1 vccd1 _15043_/D sky130_fd_sc_hd__mux2_1
XFILLER_153_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10306_ _14691_/Q _14876_/Q _10650_/S vssd1 vssd1 vccd1 vccd1 _14691_/D sky130_fd_sc_hd__mux2_1
X_14074_ _15276_/CLK _14074_/D vssd1 vssd1 vccd1 vccd1 _14074_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11286_ _15032_/Q wire438/X _11284_/X _11285_/X vssd1 vssd1 vccd1 vccd1 _15032_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_112_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13025_ _15488_/Q _13105_/A2 _13025_/B1 _13024_/X vssd1 vssd1 vccd1 vccd1 _15488_/D
+ sky130_fd_sc_hd__a22o_1
X_10237_ _14622_/Q _14775_/Q _10650_/S vssd1 vssd1 vccd1 vccd1 _14622_/D sky130_fd_sc_hd__mux2_1
XFILLER_94_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10168_ _11854_/A1 _14552_/Q _10197_/S vssd1 vssd1 vccd1 vccd1 _14552_/D sky130_fd_sc_hd__mux2_1
XFILLER_86_61 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_695 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_226 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14976_ _15020_/CLK _14976_/D vssd1 vssd1 vccd1 vccd1 _14976_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10099_ _14717_/Q _10099_/B _10099_/C vssd1 vssd1 vccd1 vccd1 _10099_/X sky130_fd_sc_hd__and3_4
XFILLER_75_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_602 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13927_ _15667_/CLK _13927_/D vssd1 vssd1 vccd1 vccd1 _13927_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_74_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13858_ _15332_/CLK _13858_/D vssd1 vssd1 vccd1 vccd1 _13858_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_616 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12809_ _15363_/Q _12765_/B _12808_/X _12809_/C1 vssd1 vssd1 vccd1 vccd1 _15363_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_50_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_108_clk clkbuf_5_26_0_clk/X vssd1 vssd1 vccd1 vccd1 _15630_/CLK sky130_fd_sc_hd__clkbuf_16
X_13789_ _15385_/CLK _13789_/D vssd1 vssd1 vccd1 vccd1 _13789_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_96_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_852 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15528_ _15536_/CLK _15528_/D vssd1 vssd1 vccd1 vccd1 _15528_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_187_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_1024 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15459_ _15645_/CLK _15459_/D vssd1 vssd1 vccd1 vccd1 _15459_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08000_ _13566_/Q _08006_/D vssd1 vssd1 vccd1 vccd1 _08000_/X sky130_fd_sc_hd__or2_1
XFILLER_175_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09951_ _11838_/A1 _14311_/Q _09963_/S vssd1 vssd1 vccd1 vccd1 _14311_/D sky130_fd_sc_hd__mux2_1
XFILLER_171_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08902_ _09130_/A _08895_/X _08898_/X _09450_/B1 vssd1 vssd1 vccd1 vccd1 _08902_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_44_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09882_ _11868_/A1 _14244_/Q _09892_/S vssd1 vssd1 vccd1 vccd1 _14244_/D sky130_fd_sc_hd__mux2_1
XTAP_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08833_ _13856_/Q _13078_/B2 _08846_/S vssd1 vssd1 vccd1 vccd1 _13856_/D sky130_fd_sc_hd__mux2_1
XFILLER_100_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1039 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08764_ _08754_/A _14613_/Q _08778_/D vssd1 vssd1 vccd1 vccd1 _08764_/X sky130_fd_sc_hd__a21o_1
XFILLER_39_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07715_ _13491_/Q _07712_/B _13492_/Q vssd1 vssd1 vccd1 vccd1 _07715_/Y sky130_fd_sc_hd__a21oi_1
XTAP_2708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08695_ _13798_/Q _08573_/S _08692_/X _08694_/X vssd1 vssd1 vccd1 vccd1 _13798_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_65_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07646_ _13473_/Q _07647_/C _13474_/Q vssd1 vssd1 vccd1 vccd1 _07646_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_54_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07577_ _07575_/Y _07588_/D _07629_/A vssd1 vssd1 vccd1 vccd1 _07577_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_15_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09316_ _08519_/A _09314_/X _09315_/X vssd1 vssd1 vccd1 vccd1 _09317_/C sky130_fd_sc_hd__a21o_1
XFILLER_15_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_1078 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09247_ _13892_/Q _09522_/A2 _08512_/B _14407_/Q _08507_/A vssd1 vssd1 vccd1 vccd1
+ _09247_/X sky130_fd_sc_hd__a221o_1
X_09178_ _09162_/X _09165_/X _09172_/X _09177_/X vssd1 vssd1 vccd1 vccd1 _09178_/X
+ sky130_fd_sc_hd__o22a_2
XFILLER_181_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08129_ input2/X input10/X _08145_/S vssd1 vssd1 vccd1 vccd1 _08129_/X sky130_fd_sc_hd__mux2_1
XFILLER_108_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_467 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11140_ _11298_/A _11058_/A _11129_/Y vssd1 vssd1 vccd1 vccd1 _11191_/B sky130_fd_sc_hd__a21oi_2
XFILLER_123_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput45 _07181_/X vssd1 vssd1 vccd1 vccd1 ext_address[19] sky130_fd_sc_hd__clkbuf_2
Xoutput56 _07164_/X vssd1 vssd1 vccd1 vccd1 ext_address[2] sky130_fd_sc_hd__clkbuf_2
Xoutput67 _07108_/X vssd1 vssd1 vccd1 vccd1 ext_write_data[0] sky130_fd_sc_hd__clkbuf_2
XFILLER_150_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput78 _07109_/X vssd1 vssd1 vccd1 vccd1 ext_write_data[1] sky130_fd_sc_hd__clkbuf_2
X_11071_ _11298_/A _11067_/X _11070_/X _11048_/Y _11069_/X vssd1 vssd1 vccd1 vccd1
+ _11071_/X sky130_fd_sc_hd__o221a_1
Xoutput89 _07110_/X vssd1 vssd1 vccd1 vccd1 ext_write_data[2] sky130_fd_sc_hd__clkbuf_2
X_10022_ _11876_/A1 _14380_/Q _10028_/S vssd1 vssd1 vccd1 vccd1 _14380_/D sky130_fd_sc_hd__mux2_1
XFILLER_103_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14830_ _15462_/CLK _14830_/D vssd1 vssd1 vccd1 vccd1 _14830_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_102_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14761_ _15638_/CLK _14761_/D vssd1 vssd1 vccd1 vccd1 _14761_/Q sky130_fd_sc_hd__dfxtp_4
X_11973_ _11956_/X _11957_/X _12582_/A vssd1 vssd1 vccd1 vccd1 _11973_/X sky130_fd_sc_hd__mux2_1
XTAP_3954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10924_ _14945_/Q _10929_/B _10923_/Y _13202_/B vssd1 vssd1 vccd1 vccd1 _14945_/D
+ sky130_fd_sc_hd__o22a_1
X_13712_ _15301_/CLK _13712_/D vssd1 vssd1 vccd1 vccd1 _13712_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14692_ _15608_/CLK _14692_/D vssd1 vssd1 vccd1 vccd1 _14692_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_186_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10855_ _14887_/Q _13781_/Q _12927_/S vssd1 vssd1 vccd1 vccd1 _14887_/D sky130_fd_sc_hd__mux2_1
XFILLER_44_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13643_ _14517_/CLK _13643_/D vssd1 vssd1 vccd1 vccd1 _13643_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_176_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13574_ _13803_/CLK _13574_/D vssd1 vssd1 vccd1 vccd1 _13574_/Q sky130_fd_sc_hd__dfxtp_4
X_10786_ _14818_/Q _15450_/Q _12929_/S vssd1 vssd1 vccd1 vccd1 _14818_/D sky130_fd_sc_hd__mux2_1
XFILLER_158_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15313_ _15510_/CLK _15313_/D vssd1 vssd1 vccd1 vccd1 _15313_/Q sky130_fd_sc_hd__dfxtp_1
X_12525_ _12508_/X _12509_/X _12617_/S vssd1 vssd1 vccd1 vccd1 _12525_/X sky130_fd_sc_hd__mux2_1
XPHY_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15244_ _15244_/CLK _15244_/D vssd1 vssd1 vccd1 vccd1 _15244_/Q sky130_fd_sc_hd__dfxtp_1
X_12456_ _12439_/X _12440_/X _12502_/S vssd1 vssd1 vccd1 vccd1 _12456_/X sky130_fd_sc_hd__mux2_1
XFILLER_184_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11407_ _13177_/A _11407_/B vssd1 vssd1 vccd1 vccd1 _11409_/B sky130_fd_sc_hd__xor2_1
X_15175_ _15212_/CLK _15175_/D vssd1 vssd1 vccd1 vccd1 _15175_/Q sky130_fd_sc_hd__dfxtp_1
X_12387_ _12370_/X _12371_/X _12617_/S vssd1 vssd1 vccd1 vccd1 _12387_/X sky130_fd_sc_hd__mux2_1
XFILLER_126_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_871 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14126_ _15676_/CLK _14126_/D vssd1 vssd1 vccd1 vccd1 _14126_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11338_ _11048_/Y _11313_/X _11337_/X _11351_/C1 vssd1 vssd1 vccd1 vccd1 _11338_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_113_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14057_ _15654_/CLK _14057_/D vssd1 vssd1 vccd1 vccd1 _14057_/Q sky130_fd_sc_hd__dfxtp_1
X_11269_ _11283_/A _08348_/X _11268_/Y _08233_/B vssd1 vssd1 vccd1 vccd1 _11269_/X
+ sky130_fd_sc_hd__o211a_1
X_13008_ _10684_/X _14883_/Q _13038_/S vssd1 vssd1 vccd1 vccd1 _13008_/X sky130_fd_sc_hd__mux2_4
XFILLER_140_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14959_ _15582_/CLK _14959_/D vssd1 vssd1 vccd1 vccd1 _14959_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07500_ _14765_/Q _07499_/X _07500_/S vssd1 vssd1 vccd1 vccd1 _07500_/X sky130_fd_sc_hd__mux2_8
XFILLER_165_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08480_ _13770_/Q _12900_/S _08479_/X vssd1 vssd1 vccd1 vccd1 _13770_/D sky130_fd_sc_hd__o21a_1
XFILLER_23_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07431_ _13663_/Q _07483_/A2 _07483_/B1 _14691_/Q _07430_/X vssd1 vssd1 vccd1 vccd1
+ _07431_/X sky130_fd_sc_hd__a221o_1
XFILLER_62_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07362_ _07362_/A _07362_/B vssd1 vssd1 vccd1 vccd1 _07363_/D sky130_fd_sc_hd__nand2_1
XFILLER_188_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09101_ _09437_/A1 _09100_/X _09099_/X _09405_/A vssd1 vssd1 vccd1 vccd1 _09101_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_188_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07293_ _13917_/Q _15504_/Q _07339_/S vssd1 vssd1 vccd1 vccd1 _07294_/A sky130_fd_sc_hd__mux2_8
XFILLER_30_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09032_ _14524_/Q _14137_/Q _14169_/Q _14105_/Q _09521_/S _09523_/A1 vssd1 vssd1
+ vccd1 vccd1 _09032_/X sky130_fd_sc_hd__mux4_1
XFILLER_136_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_176_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_724 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_148 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09934_ _13321_/A0 _14294_/Q _09963_/S vssd1 vssd1 vccd1 vccd1 _14294_/D sky130_fd_sc_hd__mux2_1
XFILLER_131_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09865_ _11851_/A _09964_/B vssd1 vssd1 vccd1 vccd1 _09865_/Y sky130_fd_sc_hd__nand2b_4
XFILLER_131_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08816_ _13350_/A0 _13842_/Q _08816_/S vssd1 vssd1 vccd1 vccd1 _13842_/D sky130_fd_sc_hd__mux2_1
XTAP_3206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09796_ _13318_/D _10132_/B vssd1 vssd1 vccd1 vccd1 _09796_/Y sky130_fd_sc_hd__nor2_8
XTAP_3217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08747_ _13541_/Q _08747_/A2 _08747_/B1 _13477_/Q _08746_/X vssd1 vssd1 vccd1 vccd1
+ _08751_/B sky130_fd_sc_hd__a221o_2
XTAP_2505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08678_ _13423_/Q _08690_/B1 _08693_/A2 _14496_/Q vssd1 vssd1 vccd1 vccd1 _08678_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_27_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07629_ _07629_/A _07629_/B vssd1 vssd1 vccd1 vccd1 _07629_/Y sky130_fd_sc_hd__nand2_1
XFILLER_26_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10640_ _14746_/Q _10639_/X _10650_/S vssd1 vssd1 vccd1 vccd1 _14746_/D sky130_fd_sc_hd__mux2_1
XFILLER_146_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10571_ _14928_/Q _13713_/Q _14927_/Q vssd1 vssd1 vccd1 vccd1 _10571_/X sky130_fd_sc_hd__or3b_1
XFILLER_158_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12310_ _12383_/A _12310_/B vssd1 vssd1 vccd1 vccd1 _12310_/X sky130_fd_sc_hd__and2_1
XFILLER_155_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13290_ _12651_/X _15622_/Q _13291_/S vssd1 vssd1 vccd1 vccd1 _15622_/D sky130_fd_sc_hd__mux2_1
XFILLER_166_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12241_ _12452_/A _12241_/B vssd1 vssd1 vccd1 vccd1 _12241_/X sky130_fd_sc_hd__and2_1
XFILLER_154_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12172_ _12452_/A _12172_/B vssd1 vssd1 vccd1 vccd1 _12172_/X sky130_fd_sc_hd__and2_1
XFILLER_174_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11123_ _10350_/Y _11375_/B _11122_/X _11371_/A vssd1 vssd1 vccd1 vccd1 _11185_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_27_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11054_ _13251_/A _13251_/B vssd1 vssd1 vccd1 vccd1 _11129_/B sky130_fd_sc_hd__nand2_4
XFILLER_114_1012 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10005_ _12967_/A1 _14363_/Q _10028_/S vssd1 vssd1 vccd1 vccd1 _14363_/D sky130_fd_sc_hd__mux2_1
XFILLER_76_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_911 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14813_ _15446_/CLK _14813_/D vssd1 vssd1 vccd1 vccd1 _14813_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14744_ _15608_/CLK _14744_/D vssd1 vssd1 vccd1 vccd1 _14744_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_3784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11956_ _14521_/Q _14134_/Q _14166_/Q _14102_/Q _12079_/S _12080_/A vssd1 vssd1 vccd1
+ vccd1 _11956_/X sky130_fd_sc_hd__mux4_1
XTAP_3795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10907_ _14936_/Q _10951_/B _10906_/Y _11399_/A vssd1 vssd1 vccd1 vccd1 _14936_/D
+ sky130_fd_sc_hd__o22a_1
X_11887_ _14518_/Q _14131_/Q _14163_/Q _14099_/Q _11993_/S _12253_/S1 vssd1 vssd1
+ vccd1 vccd1 _11887_/X sky130_fd_sc_hd__mux4_1
X_14675_ _15622_/CLK _14675_/D vssd1 vssd1 vccd1 vccd1 _14675_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13626_ _15383_/CLK _13626_/D vssd1 vssd1 vccd1 vccd1 _13626_/Q sky130_fd_sc_hd__dfxtp_1
X_10838_ _14870_/Q _13798_/Q _12910_/S vssd1 vssd1 vccd1 vccd1 _14870_/D sky130_fd_sc_hd__mux2_1
XFILLER_20_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_1051 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13557_ _15386_/CLK _13557_/D vssd1 vssd1 vccd1 vccd1 _13557_/Q sky130_fd_sc_hd__dfxtp_1
X_10769_ _14801_/Q _15433_/Q _12932_/S vssd1 vssd1 vccd1 vccd1 _14801_/D sky130_fd_sc_hd__mux2_1
XFILLER_8_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12508_ _14545_/Q _14158_/Q _14190_/Q _14126_/Q _12522_/S _12521_/A vssd1 vssd1 vccd1
+ vccd1 _12508_/X sky130_fd_sc_hd__mux4_1
X_13488_ _14495_/CLK _13488_/D vssd1 vssd1 vccd1 vccd1 _13488_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_146_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_163 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15227_ _15259_/CLK _15227_/D vssd1 vssd1 vccd1 vccd1 _15227_/Q sky130_fd_sc_hd__dfxtp_1
X_12439_ _14542_/Q _14155_/Q _14187_/Q _14123_/Q _12453_/S _12452_/A vssd1 vssd1 vccd1
+ vccd1 _12439_/X sky130_fd_sc_hd__mux4_1
XFILLER_59_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15158_ _15259_/CLK _15158_/D vssd1 vssd1 vccd1 vccd1 _15158_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14109_ _15674_/CLK _14109_/D vssd1 vssd1 vccd1 vccd1 _14109_/Q sky130_fd_sc_hd__dfxtp_1
X_07980_ _14753_/Q _07971_/A _07979_/X _07987_/C1 vssd1 vssd1 vccd1 vccd1 _13560_/D
+ sky130_fd_sc_hd__o211a_1
X_15089_ _15331_/CLK _15089_/D vssd1 vssd1 vccd1 vccd1 _15089_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout109 _13288_/S vssd1 vssd1 vccd1 vccd1 _13291_/S sky130_fd_sc_hd__buf_12
XFILLER_101_407 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06931_ _06931_/A _06931_/B vssd1 vssd1 vccd1 vccd1 _06931_/Y sky130_fd_sc_hd__nand2_1
XFILLER_110_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09650_ _14023_/Q _13092_/B2 _09661_/S vssd1 vssd1 vccd1 vccd1 _14023_/D sky130_fd_sc_hd__mux2_1
XFILLER_80_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06862_ _12640_/S _12785_/B vssd1 vssd1 vccd1 vccd1 _06863_/B sky130_fd_sc_hd__nand2_2
XFILLER_55_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08601_ _13530_/Q _08683_/A2 _08750_/B1 _13633_/Q _08600_/X vssd1 vssd1 vccd1 vccd1
+ _08605_/B sky130_fd_sc_hd__a221o_1
XFILLER_95_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09581_ _13957_/Q _13337_/A0 _09594_/S vssd1 vssd1 vccd1 vccd1 _13957_/D sky130_fd_sc_hd__mux2_1
X_06793_ _14587_/Q _06789_/B _08391_/B _08421_/A vssd1 vssd1 vccd1 vccd1 _06799_/A
+ sky130_fd_sc_hd__o211ai_2
XFILLER_94_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08532_ _08538_/A _08532_/B vssd1 vssd1 vccd1 vccd1 _08532_/Y sky130_fd_sc_hd__nor2_8
XFILLER_70_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08463_ _13762_/Q _12900_/S _08426_/X vssd1 vssd1 vccd1 vccd1 _08463_/X sky130_fd_sc_hd__o21a_1
XFILLER_168_407 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07414_ _14655_/Q _07474_/B _07482_/C vssd1 vssd1 vccd1 vccd1 _07414_/X sky130_fd_sc_hd__and3_1
X_08394_ _08469_/A _08390_/X _08400_/C _13138_/S vssd1 vssd1 vccd1 vccd1 _08394_/X
+ sky130_fd_sc_hd__o31a_2
X_07345_ _07343_/X _07344_/X _07360_/B vssd1 vssd1 vccd1 vccd1 _07345_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_177_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_30_clk clkbuf_5_6_0_clk/X vssd1 vssd1 vccd1 vccd1 _15501_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_137_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07276_ _10360_/A vssd1 vssd1 vccd1 vccd1 _07278_/A sky130_fd_sc_hd__inv_2
XFILLER_176_495 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09015_ _13912_/Q _10877_/S _09014_/X vssd1 vssd1 vccd1 vccd1 _13912_/D sky130_fd_sc_hd__a21o_1
XFILLER_145_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout610 _12470_/S vssd1 vssd1 vccd1 vccd1 _12453_/S sky130_fd_sc_hd__buf_12
Xfanout621 _12612_/S vssd1 vssd1 vccd1 vccd1 _12614_/S sky130_fd_sc_hd__buf_12
X_09917_ _07448_/X _14278_/Q _09930_/S vssd1 vssd1 vccd1 vccd1 _14278_/D sky130_fd_sc_hd__mux2_1
Xfanout632 _13739_/Q vssd1 vssd1 vccd1 vccd1 _13242_/A sky130_fd_sc_hd__clkbuf_16
Xfanout643 _07965_/C1 vssd1 vssd1 vccd1 vccd1 _07949_/C1 sky130_fd_sc_hd__buf_8
XFILLER_86_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_97_clk clkbuf_5_24_0_clk/X vssd1 vssd1 vccd1 vccd1 _15623_/CLK sky130_fd_sc_hd__clkbuf_16
X_09848_ _14212_/Q _11868_/A1 _09858_/S vssd1 vssd1 vccd1 vccd1 _14212_/D sky130_fd_sc_hd__mux2_1
XTAP_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09779_ _14146_/Q _13082_/B2 _09790_/S vssd1 vssd1 vccd1 vccd1 _14146_/D sky130_fd_sc_hd__mux2_1
XTAP_2302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11810_ _15233_/Q _11876_/A1 _11816_/S vssd1 vssd1 vccd1 vccd1 _15233_/D sky130_fd_sc_hd__mux2_1
XTAP_2324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12790_ _15360_/Q _12789_/C _15361_/Q vssd1 vssd1 vccd1 vccd1 _13309_/C sky130_fd_sc_hd__a21oi_1
XTAP_2335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_379 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11741_ _15170_/Q _13349_/A0 _11741_/S vssd1 vssd1 vccd1 vccd1 _15170_/D sky130_fd_sc_hd__mux2_1
XTAP_2368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14460_ _15178_/CLK _14460_/D vssd1 vssd1 vccd1 vccd1 _14460_/Q sky130_fd_sc_hd__dfxtp_1
X_11672_ _11847_/A1 _15104_/Q _11675_/S vssd1 vssd1 vccd1 vccd1 _15104_/D sky130_fd_sc_hd__mux2_1
XTAP_1678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10623_ _14971_/Q _10718_/A2 _10722_/B1 _14939_/Q _10622_/X vssd1 vssd1 vccd1 vccd1
+ _10623_/X sky130_fd_sc_hd__a221o_1
X_13411_ _15677_/CLK _13411_/D vssd1 vssd1 vccd1 vccd1 _13411_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14391_ _15077_/CLK _14391_/D vssd1 vssd1 vccd1 vccd1 _14391_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_21_clk clkbuf_5_3_0_clk/X vssd1 vssd1 vccd1 vccd1 _15315_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_6_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13342_ _13342_/A0 _15672_/Q _13350_/S vssd1 vssd1 vccd1 vccd1 _15672_/D sky130_fd_sc_hd__mux2_1
XFILLER_127_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10554_ _10554_/A _10554_/B vssd1 vssd1 vccd1 vccd1 _10555_/D sky130_fd_sc_hd__and2_1
XFILLER_182_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13273_ _15357_/Q _15604_/Q _13309_/A vssd1 vssd1 vccd1 vccd1 _15604_/D sky130_fd_sc_hd__mux2_1
X_10485_ _10520_/A1 _13784_/Q _13752_/Q _10520_/B2 vssd1 vssd1 vccd1 vccd1 _10485_/X
+ sky130_fd_sc_hd__a22o_1
X_15012_ _15577_/CLK _15012_/D vssd1 vssd1 vccd1 vccd1 _15012_/Q sky130_fd_sc_hd__dfxtp_1
X_12224_ _12477_/A1 _12223_/X _12500_/B1 vssd1 vssd1 vccd1 vccd1 _12224_/X sky130_fd_sc_hd__a21o_1
XFILLER_108_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12155_ _12500_/A1 _12154_/X _12500_/B1 vssd1 vssd1 vccd1 vccd1 _12155_/X sky130_fd_sc_hd__a21o_1
XFILLER_64_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_939 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11106_ _11347_/A _11156_/B _11105_/X vssd1 vssd1 vccd1 vccd1 _11181_/B sky130_fd_sc_hd__o21ai_2
XFILLER_1_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12086_ _12500_/A1 _12085_/X _12468_/A1 vssd1 vssd1 vccd1 vccd1 _12086_/X sky130_fd_sc_hd__a21o_1
XFILLER_68_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_88_clk clkbuf_5_13_0_clk/X vssd1 vssd1 vccd1 vccd1 _14892_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_110_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11037_ _11037_/A _11500_/A vssd1 vssd1 vccd1 vccd1 _11249_/B sky130_fd_sc_hd__and2_1
XFILLER_37_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12988_ _13080_/B2 _13024_/A2 _12987_/X _13024_/B2 vssd1 vssd1 vccd1 vccd1 _12988_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_3592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14727_ _15552_/CLK _14727_/D vssd1 vssd1 vccd1 vccd1 _14727_/Q sky130_fd_sc_hd__dfxtp_1
X_11939_ _12615_/B1 _11936_/X _12616_/C1 vssd1 vssd1 vccd1 vccd1 _11939_/X sky130_fd_sc_hd__o21a_1
XFILLER_162_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14658_ _15446_/CLK _14658_/D vssd1 vssd1 vccd1 vccd1 _14658_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13609_ _15647_/CLK _13609_/D vssd1 vssd1 vccd1 vccd1 _13609_/Q sky130_fd_sc_hd__dfxtp_2
X_14589_ _14612_/CLK _14589_/D vssd1 vssd1 vccd1 vccd1 _14589_/Q sky130_fd_sc_hd__dfxtp_2
Xclkbuf_leaf_12_clk clkbuf_5_2_0_clk/X vssd1 vssd1 vccd1 vccd1 _15286_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_119_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07130_ _14845_/Q _14837_/Q _08150_/S vssd1 vssd1 vccd1 vccd1 _07131_/B sky130_fd_sc_hd__mux2_1
XFILLER_146_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07061_ _07060_/X _13599_/Q _12728_/S vssd1 vssd1 vccd1 vccd1 _07061_/X sky130_fd_sc_hd__mux2_1
XFILLER_146_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07963_ _07973_/D _07963_/B vssd1 vssd1 vccd1 vccd1 _07964_/B sky130_fd_sc_hd__nand2b_1
XFILLER_59_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_79_clk clkbuf_5_15_0_clk/X vssd1 vssd1 vccd1 vccd1 _15606_/CLK sky130_fd_sc_hd__clkbuf_16
X_06914_ _15390_/Q _07621_/A _15389_/Q _06711_/Y vssd1 vssd1 vccd1 vccd1 _06920_/B
+ sky130_fd_sc_hd__a22o_1
X_09702_ _11857_/A1 _14072_/Q _09728_/S vssd1 vssd1 vccd1 vccd1 _14072_/D sky130_fd_sc_hd__mux2_1
XFILLER_114_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07894_ _13537_/Q _07900_/C _13538_/Q vssd1 vssd1 vccd1 vccd1 _07894_/X sky130_fd_sc_hd__a21o_1
XFILLER_56_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09633_ _14006_/Q _11680_/A0 _09660_/S vssd1 vssd1 vccd1 vccd1 _14006_/D sky130_fd_sc_hd__mux2_1
X_06845_ _12379_/A _06845_/B vssd1 vssd1 vccd1 vccd1 _06845_/Y sky130_fd_sc_hd__nand2_1
XFILLER_55_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09564_ _13940_/Q _11853_/A1 _09594_/S vssd1 vssd1 vccd1 vccd1 _13940_/D sky130_fd_sc_hd__mux2_1
X_06776_ _07188_/S vssd1 vssd1 vccd1 vccd1 _06865_/B sky130_fd_sc_hd__inv_4
XFILLER_130_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08515_ _14613_/Q _14614_/Q vssd1 vssd1 vccd1 vccd1 _13133_/C sky130_fd_sc_hd__nand2_1
X_09495_ _14385_/Q _15201_/Q _13840_/Q _14579_/Q _09512_/S _08494_/B vssd1 vssd1 vccd1
+ vccd1 _09496_/B sky130_fd_sc_hd__mux4_1
XFILLER_51_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08446_ _13753_/Q _12906_/S _08426_/B _08445_/X vssd1 vssd1 vccd1 vccd1 _13753_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_11_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08377_ _08337_/X _08376_/X _11297_/S vssd1 vssd1 vccd1 vccd1 _11290_/B sky130_fd_sc_hd__mux2_1
XFILLER_23_298 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07328_ _15307_/Q _15463_/Q _07335_/S vssd1 vssd1 vccd1 vccd1 _07329_/A sky130_fd_sc_hd__mux2_4
XFILLER_139_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07259_ _07261_/A _07261_/B _07256_/X _07258_/Y vssd1 vssd1 vccd1 vccd1 _07270_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_165_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_487 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10270_ _14655_/Q _14808_/Q _10630_/S vssd1 vssd1 vccd1 vccd1 _14655_/D sky130_fd_sc_hd__mux2_1
XFILLER_180_958 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout440 _07374_/X vssd1 vssd1 vccd1 vccd1 _07499_/B1 sky130_fd_sc_hd__buf_12
Xfanout451 _10695_/S vssd1 vssd1 vccd1 vccd1 _10285_/S sky130_fd_sc_hd__clkbuf_16
Xfanout462 _06675_/Y vssd1 vssd1 vccd1 vccd1 _09445_/C1 sky130_fd_sc_hd__buf_12
XFILLER_93_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout473 _12168_/A vssd1 vssd1 vccd1 vccd1 _12582_/A sky130_fd_sc_hd__buf_12
XFILLER_48_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13960_ _15304_/CLK _13960_/D vssd1 vssd1 vccd1 vccd1 _13960_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout484 _12615_/A1 vssd1 vssd1 vccd1 vccd1 _12592_/A1 sky130_fd_sc_hd__buf_12
XFILLER_171_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout495 _15043_/Q vssd1 vssd1 vccd1 vccd1 _08150_/S sky130_fd_sc_hd__buf_12
XFILLER_47_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12911_ _15439_/Q _15625_/Q _12918_/S vssd1 vssd1 vccd1 vccd1 _15439_/D sky130_fd_sc_hd__mux2_1
XFILLER_47_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13891_ _15665_/CLK _13891_/D vssd1 vssd1 vccd1 vccd1 _13891_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_1048 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15630_ _15630_/CLK _15630_/D vssd1 vssd1 vccd1 vccd1 _15630_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12842_ _14736_/Q _15370_/Q _12871_/S vssd1 vssd1 vccd1 vccd1 _15370_/D sky130_fd_sc_hd__mux2_1
XFILLER_73_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15561_ _15570_/CLK _15561_/D vssd1 vssd1 vccd1 vccd1 _15561_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12773_ _06861_/Y _12770_/X _12771_/X _12772_/X vssd1 vssd1 vccd1 vccd1 _12773_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_15_744 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14512_ _15397_/CLK _14512_/D vssd1 vssd1 vccd1 vccd1 _14512_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11724_ _15153_/Q _13332_/A0 _11741_/S vssd1 vssd1 vccd1 vccd1 _15153_/D sky130_fd_sc_hd__mux2_1
XTAP_1475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15492_ _15499_/CLK _15492_/D vssd1 vssd1 vccd1 vccd1 _15492_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11655_ _13074_/B2 _15087_/Q _11670_/S vssd1 vssd1 vccd1 vccd1 _15087_/D sky130_fd_sc_hd__mux2_1
X_14443_ _15300_/CLK _14443_/D vssd1 vssd1 vccd1 vccd1 _14443_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_175_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10606_ _15559_/Q _10731_/B vssd1 vssd1 vccd1 vccd1 _10606_/X sky130_fd_sc_hd__and2_1
X_11586_ _11586_/A _11586_/B vssd1 vssd1 vccd1 vccd1 _11586_/Y sky130_fd_sc_hd__nand2_1
X_14374_ _15291_/CLK _14374_/D vssd1 vssd1 vccd1 vccd1 _14374_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_167_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10537_ _10537_/A _10537_/B _10537_/C vssd1 vssd1 vccd1 vccd1 _10548_/B sky130_fd_sc_hd__or3_1
X_13325_ _13325_/A0 _15655_/Q _13350_/S vssd1 vssd1 vccd1 vccd1 _15655_/D sky130_fd_sc_hd__mux2_1
XFILLER_128_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10468_ _11598_/A _13233_/B vssd1 vssd1 vccd1 vccd1 _10469_/B sky130_fd_sc_hd__and2b_1
X_13256_ _15340_/Q _15587_/Q _13282_/S vssd1 vssd1 vccd1 vccd1 _15587_/D sky130_fd_sc_hd__mux2_1
XFILLER_142_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12207_ _14242_/Q _14274_/Q _14306_/Q _14338_/Q _12489_/S0 _12489_/S1 vssd1 vssd1
+ vccd1 vccd1 _12207_/X sky130_fd_sc_hd__mux4_1
X_13187_ _13229_/A _11440_/A _13219_/S vssd1 vssd1 vccd1 vccd1 _13187_/X sky130_fd_sc_hd__o21a_1
XFILLER_69_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10399_ _10399_/A _10399_/B vssd1 vssd1 vccd1 vccd1 _10556_/A sky130_fd_sc_hd__or2_1
XFILLER_111_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12138_ _14239_/Q _14271_/Q _14303_/Q _14335_/Q _12472_/S _12465_/S1 vssd1 vssd1
+ vccd1 vccd1 _12138_/X sky130_fd_sc_hd__mux4_1
XFILLER_69_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12069_ _14236_/Q _14268_/Q _14300_/Q _14332_/Q _12470_/S _12080_/A vssd1 vssd1 vccd1
+ vccd1 _12069_/X sky130_fd_sc_hd__mux4_1
XFILLER_38_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_1_clk clkbuf_5_0_0_clk/X vssd1 vssd1 vccd1 vccd1 _15284_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_84_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08300_ _13719_/Q _08232_/A _11351_/C1 _08299_/X vssd1 vssd1 vccd1 vccd1 _13719_/D
+ sky130_fd_sc_hd__a22o_1
X_09280_ _08510_/B _09276_/X _09279_/X _09275_/X vssd1 vssd1 vccd1 vccd1 _09281_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_166_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08231_ _07322_/X _10457_/A2 _08229_/X vssd1 vssd1 vccd1 vccd1 _08231_/X sky130_fd_sc_hd__a21o_4
XFILLER_166_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08162_ _13668_/Q _10285_/S _08155_/X _08161_/X vssd1 vssd1 vccd1 vccd1 _13668_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_158_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07113_ _14835_/Q _07115_/B _07157_/A vssd1 vssd1 vccd1 vccd1 _07113_/X sky130_fd_sc_hd__and3_4
X_08093_ _08154_/B _08093_/B vssd1 vssd1 vccd1 vccd1 _08093_/Y sky130_fd_sc_hd__nand2b_2
XFILLER_109_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07044_ _07043_/X _14747_/Q _07077_/S vssd1 vssd1 vccd1 vccd1 _13593_/D sky130_fd_sc_hd__mux2_1
XFILLER_118_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_1031 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08995_ _15278_/Q _15246_/Q _15214_/Q _15145_/Q _09005_/S _09511_/S1 vssd1 vssd1
+ vccd1 vccd1 _08995_/X sky130_fd_sc_hd__mux4_1
XFILLER_47_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07946_ _13552_/Q _13551_/Q _13550_/Q _07946_/D vssd1 vssd1 vccd1 vccd1 _07961_/C
+ sky130_fd_sc_hd__and4_4
XFILLER_75_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07877_ _07884_/C _07884_/D vssd1 vssd1 vccd1 vccd1 _07881_/B sky130_fd_sc_hd__nand2_1
X_09616_ _13990_/Q _11838_/A1 _09628_/S vssd1 vssd1 vccd1 vccd1 _13990_/D sky130_fd_sc_hd__mux2_1
X_06828_ _14730_/Q _14709_/Q _12640_/S vssd1 vssd1 vccd1 vccd1 _08036_/A sky130_fd_sc_hd__and3_2
XFILLER_44_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06759_ input17/X vssd1 vssd1 vccd1 vccd1 _06759_/Y sky130_fd_sc_hd__inv_2
X_09547_ _08497_/A _09545_/X _09546_/X _08507_/Y _13049_/A1 vssd1 vssd1 vccd1 vccd1
+ _09547_/X sky130_fd_sc_hd__a221o_1
XFILLER_24_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09478_ _14256_/Q _14288_/Q _14320_/Q _14352_/Q _09551_/S _09553_/A1 vssd1 vssd1
+ vccd1 vccd1 _09478_/X sky130_fd_sc_hd__mux4_1
XFILLER_180_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08429_ _14612_/Q _08390_/C _08425_/X _10764_/S vssd1 vssd1 vccd1 vccd1 _08429_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_156_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11440_ _11440_/A _11440_/B vssd1 vssd1 vccd1 vccd1 _11440_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_11_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_780 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11371_ _11371_/A _11371_/B vssd1 vssd1 vccd1 vccd1 _11375_/C sky130_fd_sc_hd__or2_1
XFILLER_164_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13110_ _13032_/X _13118_/A2 _13114_/B1 _13110_/B2 vssd1 vssd1 vccd1 vccd1 _13110_/X
+ sky130_fd_sc_hd__a22o_1
X_10322_ _14707_/Q _14892_/Q _10730_/S vssd1 vssd1 vccd1 vccd1 _14707_/D sky130_fd_sc_hd__mux2_1
XFILLER_30_1071 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14090_ _15328_/CLK _14090_/D vssd1 vssd1 vccd1 vccd1 _14090_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_124_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13041_ _08501_/A _08724_/B _10877_/S vssd1 vssd1 vccd1 vccd1 _13041_/Y sky130_fd_sc_hd__a21oi_4
X_10253_ _14638_/Q _14791_/Q _10285_/S vssd1 vssd1 vccd1 vccd1 _14638_/D sky130_fd_sc_hd__mux2_1
X_10184_ _11870_/A1 _14568_/Q _10197_/S vssd1 vssd1 vccd1 vccd1 _14568_/D sky130_fd_sc_hd__mux2_1
XFILLER_59_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14992_ _15582_/CLK _14992_/D vssd1 vssd1 vccd1 vccd1 _14992_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout270 _08513_/Y vssd1 vssd1 vccd1 vccd1 _08693_/A2 sky130_fd_sc_hd__buf_8
XFILLER_19_302 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout292 _07484_/X vssd1 vssd1 vccd1 vccd1 _11879_/A1 sky130_fd_sc_hd__buf_4
X_13943_ _15665_/CLK _13943_/D vssd1 vssd1 vccd1 vccd1 _13943_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13874_ _14485_/CLK _13874_/D vssd1 vssd1 vccd1 vccd1 _13874_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_74_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15613_ _15613_/CLK _15613_/D vssd1 vssd1 vccd1 vccd1 _15613_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12825_ _15365_/Q _12759_/B _12824_/X _12832_/C1 vssd1 vssd1 vccd1 vccd1 _15365_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_27_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15544_ _15544_/CLK _15544_/D vssd1 vssd1 vccd1 vccd1 _15544_/Q sky130_fd_sc_hd__dfxtp_1
X_12756_ _15063_/Q _12755_/X _12834_/B vssd1 vssd1 vccd1 vccd1 _12756_/X sky130_fd_sc_hd__mux2_1
XTAP_1261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11707_ _11816_/A1 _15138_/Q _11708_/S vssd1 vssd1 vccd1 vccd1 _15138_/D sky130_fd_sc_hd__mux2_1
XTAP_1294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15475_ _15520_/CLK _15475_/D vssd1 vssd1 vccd1 vccd1 _15475_/Q sky130_fd_sc_hd__dfxtp_1
X_12687_ _15347_/Q _12688_/B vssd1 vssd1 vccd1 vccd1 _12701_/C sky130_fd_sc_hd__and2_2
XFILLER_147_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_922 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14426_ _15284_/CLK _14426_/D vssd1 vssd1 vccd1 vccd1 _14426_/Q sky130_fd_sc_hd__dfxtp_1
X_11638_ _13242_/A _10530_/B _11632_/B vssd1 vssd1 vccd1 vccd1 _11639_/B sky130_fd_sc_hd__o21ai_1
XFILLER_156_730 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14357_ _15077_/CLK _14357_/D vssd1 vssd1 vccd1 vccd1 _14357_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11569_ _11561_/A _11569_/B _13218_/A _11569_/D vssd1 vssd1 vccd1 vccd1 _11589_/C
+ sky130_fd_sc_hd__and4b_1
XFILLER_144_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_402 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13308_ _15640_/Q _12783_/X _13316_/S vssd1 vssd1 vccd1 vccd1 _15640_/D sky130_fd_sc_hd__mux2_1
Xmax_cap437 wire438/X vssd1 vssd1 vccd1 vccd1 _11302_/A sky130_fd_sc_hd__buf_4
XFILLER_170_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14288_ _14482_/CLK _14288_/D vssd1 vssd1 vccd1 vccd1 _14288_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_157_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13239_ _06769_/Y wire360/X _11610_/A vssd1 vssd1 vccd1 vccd1 _13239_/X sky130_fd_sc_hd__o21a_1
XFILLER_41_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07800_ _14738_/Q _07816_/A _07799_/Y _08084_/C1 vssd1 vssd1 vccd1 vccd1 _13513_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_69_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08780_ _08910_/S _08779_/X _10892_/B _13808_/Q vssd1 vssd1 vccd1 vccd1 _13808_/D
+ sky130_fd_sc_hd__a2bb2o_1
X_07731_ _13496_/Q _13495_/Q _13494_/Q _13493_/Q vssd1 vssd1 vccd1 vccd1 _07732_/C
+ sky130_fd_sc_hd__and4_1
XFILLER_65_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07662_ _07777_/A _07662_/B vssd1 vssd1 vccd1 vccd1 _07662_/Y sky130_fd_sc_hd__nand2_1
XFILLER_93_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09401_ _09406_/S1 _09399_/X _09400_/X vssd1 vssd1 vccd1 vccd1 _09405_/B sky130_fd_sc_hd__a21o_1
X_07593_ _14748_/Q _07607_/A _07592_/Y _07965_/C1 vssd1 vssd1 vccd1 vccd1 _13459_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_53_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09332_ _14475_/Q _09536_/A2 _09331_/X _13125_/B vssd1 vssd1 vccd1 vccd1 _09332_/X
+ sky130_fd_sc_hd__a211o_1
X_09263_ _08507_/A _09262_/X _09261_/X _09524_/A vssd1 vssd1 vccd1 vccd1 _09263_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_33_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08214_ _13705_/Q _11876_/A1 _08216_/S vssd1 vssd1 vccd1 vccd1 _13705_/D sky130_fd_sc_hd__mux2_1
XFILLER_14_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09194_ _14532_/Q _14145_/Q _14177_/Q _14113_/Q _09190_/S _09429_/S1 vssd1 vssd1
+ vccd1 vccd1 _09194_/X sky130_fd_sc_hd__mux4_1
XFILLER_147_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08145_ input6/X input15/X _08145_/S vssd1 vssd1 vccd1 vccd1 _08145_/X sky130_fd_sc_hd__mux2_1
XFILLER_135_903 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08076_ _14734_/Q _08083_/A _08075_/X _08084_/C1 vssd1 vssd1 vccd1 vccd1 _13644_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_134_435 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07027_ _14621_/Q _14653_/Q _07078_/S vssd1 vssd1 vccd1 vccd1 _07027_/X sky130_fd_sc_hd__mux2_1
XFILLER_136_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08978_ _09449_/B2 _08976_/X _08977_/X _09449_/A1 _06676_/A vssd1 vssd1 vccd1 vccd1
+ _08978_/X sky130_fd_sc_hd__a221o_1
X_07929_ _13547_/Q _07935_/D vssd1 vssd1 vccd1 vccd1 _07929_/X sky130_fd_sc_hd__or2_1
XFILLER_57_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10940_ _11598_/A _13233_/B vssd1 vssd1 vccd1 vccd1 _10940_/X sky130_fd_sc_hd__or2_1
XFILLER_45_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10871_ _13038_/S _13735_/Q _10871_/S vssd1 vssd1 vccd1 vccd1 _14903_/D sky130_fd_sc_hd__mux2_1
XPHY_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12610_ _13906_/Q _14421_/Q _12612_/S vssd1 vssd1 vccd1 vccd1 _12610_/X sky130_fd_sc_hd__mux2_1
XFILLER_71_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13590_ _15453_/CLK _13590_/D vssd1 vssd1 vccd1 vccd1 _13590_/Q sky130_fd_sc_hd__dfxtp_2
XPHY_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12541_ _13903_/Q _14418_/Q _12541_/S vssd1 vssd1 vccd1 vccd1 _12541_/X sky130_fd_sc_hd__mux2_1
XFILLER_12_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15260_ _15275_/CLK _15260_/D vssd1 vssd1 vccd1 vccd1 _15260_/Q sky130_fd_sc_hd__dfxtp_1
X_12472_ _13900_/Q _14415_/Q _12472_/S vssd1 vssd1 vccd1 vccd1 _12472_/X sky130_fd_sc_hd__mux2_1
XFILLER_185_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_87 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14211_ _15332_/CLK _14211_/D vssd1 vssd1 vccd1 vccd1 _14211_/Q sky130_fd_sc_hd__dfxtp_1
X_11423_ _11423_/A _11423_/B _11423_/C _11423_/D vssd1 vssd1 vccd1 vccd1 _11423_/X
+ sky130_fd_sc_hd__and4_2
X_15191_ _15292_/CLK _15191_/D vssd1 vssd1 vccd1 vccd1 _15191_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_9 _09054_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14142_ _15253_/CLK _14142_/D vssd1 vssd1 vccd1 vccd1 _14142_/Q sky130_fd_sc_hd__dfxtp_1
X_11354_ _14929_/D _14928_/D _14927_/D vssd1 vssd1 vccd1 vccd1 _11354_/X sky130_fd_sc_hd__or3_2
XFILLER_180_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10305_ _14690_/Q _14875_/Q _10650_/S vssd1 vssd1 vccd1 vccd1 _14690_/D sky130_fd_sc_hd__mux2_1
XFILLER_4_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14073_ _15178_/CLK _14073_/D vssd1 vssd1 vccd1 vccd1 _14073_/Q sky130_fd_sc_hd__dfxtp_1
X_11285_ _11283_/A _11380_/A _08290_/X _08232_/A vssd1 vssd1 vccd1 vccd1 _11285_/X
+ sky130_fd_sc_hd__a31o_1
X_10236_ _14621_/Q _14774_/Q _10285_/S vssd1 vssd1 vccd1 vccd1 _14621_/D sky130_fd_sc_hd__mux2_1
X_13024_ _13104_/B2 _13024_/A2 _13023_/X _13024_/B2 vssd1 vssd1 vccd1 vccd1 _13024_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_67_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10167_ _11853_/A1 _14551_/Q _10197_/S vssd1 vssd1 vccd1 vccd1 _14551_/D sky130_fd_sc_hd__mux2_1
XFILLER_117_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14975_ _15577_/CLK _14975_/D vssd1 vssd1 vccd1 vccd1 _14975_/Q sky130_fd_sc_hd__dfxtp_1
X_10098_ _10098_/A _10098_/B vssd1 vssd1 vccd1 vccd1 _10099_/C sky130_fd_sc_hd__nor2_1
XFILLER_48_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13926_ _15077_/CLK _13926_/D vssd1 vssd1 vccd1 vccd1 _13926_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_35_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13857_ _14468_/CLK _13857_/D vssd1 vssd1 vccd1 vccd1 _13857_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12808_ _06861_/Y _12805_/X _12806_/X _12807_/X vssd1 vssd1 vccd1 vccd1 _12808_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_62_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13788_ _14495_/CLK _13788_/D vssd1 vssd1 vccd1 vccd1 _13788_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_31_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15527_ _15527_/CLK _15527_/D vssd1 vssd1 vccd1 vccd1 _15527_/Q sky130_fd_sc_hd__dfxtp_4
X_12739_ _15354_/Q _12745_/C vssd1 vssd1 vccd1 vccd1 _12739_/X sky130_fd_sc_hd__xor2_1
XTAP_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_302 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_1088 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15458_ _15644_/CLK _15458_/D vssd1 vssd1 vccd1 vccd1 _15458_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14409_ _15127_/CLK _14409_/D vssd1 vssd1 vccd1 vccd1 _14409_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15389_ _15389_/CLK _15389_/D vssd1 vssd1 vccd1 vccd1 _15389_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09950_ _13337_/A0 _14310_/Q _09963_/S vssd1 vssd1 vccd1 vccd1 _14310_/D sky130_fd_sc_hd__mux2_1
XFILLER_89_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08901_ _09449_/A1 _08899_/X _08900_/X _09449_/B2 vssd1 vssd1 vccd1 vccd1 _08901_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_98_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09881_ _13334_/A0 _14243_/Q _09892_/S vssd1 vssd1 vccd1 vccd1 _14243_/D sky130_fd_sc_hd__mux2_1
XFILLER_170_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08832_ _13855_/Q _11689_/A0 _08846_/S vssd1 vssd1 vccd1 vccd1 _13855_/D sky130_fd_sc_hd__mux2_1
XTAP_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08763_ _08778_/D _08762_/X _06808_/X vssd1 vssd1 vccd1 vccd1 _08763_/X sky130_fd_sc_hd__o21a_1
XFILLER_85_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07714_ _14748_/Q _07713_/A _07713_/Y _07949_/C1 vssd1 vssd1 vccd1 vccd1 _13491_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_122_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08694_ _13549_/Q _08747_/A2 _08693_/X _08722_/A vssd1 vssd1 vccd1 vccd1 _08694_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_65_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07645_ _14762_/Q _07644_/A _07644_/Y _08016_/C1 vssd1 vssd1 vccd1 vccd1 _13473_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_80_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07576_ _13455_/Q _13452_/Q _07576_/C _07576_/D vssd1 vssd1 vccd1 vccd1 _07588_/D
+ sky130_fd_sc_hd__and4_2
X_09315_ _14087_/Q _13123_/B _09519_/B1 _14055_/Q _09543_/A vssd1 vssd1 vccd1 vccd1
+ _09315_/X sky130_fd_sc_hd__a221o_1
XFILLER_139_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09246_ _13956_/Q _13698_/Q _09557_/S vssd1 vssd1 vccd1 vccd1 _09246_/X sky130_fd_sc_hd__mux2_1
XFILLER_178_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09177_ _09421_/A1 _09173_/X _09176_/X vssd1 vssd1 vccd1 vccd1 _09177_/X sky130_fd_sc_hd__a21o_1
XFILLER_31_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08128_ _13658_/Q _10285_/S _08119_/X _08127_/X vssd1 vssd1 vccd1 vccd1 _13658_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_181_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_766 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08059_ _14752_/Q _13630_/Q _08072_/S vssd1 vssd1 vccd1 vccd1 _13630_/D sky130_fd_sc_hd__mux2_1
XFILLER_107_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput46 _07182_/X vssd1 vssd1 vccd1 vccd1 ext_address[20] sky130_fd_sc_hd__clkbuf_2
Xoutput57 _07192_/X vssd1 vssd1 vccd1 vccd1 ext_address[30] sky130_fd_sc_hd__clkbuf_2
X_11070_ _10987_/B _10998_/Y _11088_/S vssd1 vssd1 vccd1 vccd1 _11070_/X sky130_fd_sc_hd__mux2_2
XFILLER_0_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput68 _07121_/X vssd1 vssd1 vccd1 vccd1 ext_write_data[10] sky130_fd_sc_hd__clkbuf_2
Xoutput79 _07141_/X vssd1 vssd1 vccd1 vccd1 ext_write_data[20] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10021_ _13098_/B2 _14379_/Q _10029_/S vssd1 vssd1 vccd1 vccd1 _14379_/D sky130_fd_sc_hd__mux2_1
XFILLER_131_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_89 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14760_ _15591_/CLK _14760_/D vssd1 vssd1 vccd1 vccd1 _14760_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_3944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11972_ _11965_/X _11967_/X _11969_/X _11971_/X _12455_/C1 vssd1 vssd1 vccd1 vccd1
+ _11972_/X sky130_fd_sc_hd__o221a_1
XFILLER_17_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13711_ _15679_/CLK _13711_/D vssd1 vssd1 vccd1 vccd1 _13711_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10923_ _11496_/B _10929_/B vssd1 vssd1 vccd1 vccd1 _10923_/Y sky130_fd_sc_hd__nand2_1
XFILLER_44_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14691_ _15592_/CLK _14691_/D vssd1 vssd1 vccd1 vccd1 _14691_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13642_ _13642_/CLK _13642_/D vssd1 vssd1 vccd1 vccd1 _13642_/Q sky130_fd_sc_hd__dfxtp_1
X_10854_ _14886_/Q _13782_/Q _12927_/S vssd1 vssd1 vccd1 vccd1 _14886_/D sky130_fd_sc_hd__mux2_1
XFILLER_13_820 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13573_ _13803_/CLK _13573_/D vssd1 vssd1 vccd1 vccd1 _13573_/Q sky130_fd_sc_hd__dfxtp_1
X_10785_ _14817_/Q _15449_/Q _12928_/S vssd1 vssd1 vccd1 vccd1 _14817_/D sky130_fd_sc_hd__mux2_1
XPHY_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15312_ _15517_/CLK _15312_/D vssd1 vssd1 vccd1 vccd1 _15312_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12524_ _12517_/X _12519_/X _12521_/X _12523_/X _08405_/C vssd1 vssd1 vccd1 vccd1
+ _12524_/X sky130_fd_sc_hd__o221a_1
XPHY_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15243_ _15275_/CLK _15243_/D vssd1 vssd1 vccd1 vccd1 _15243_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_184_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12455_ _12448_/X _12450_/X _12452_/X _12454_/X _12455_/C1 vssd1 vssd1 vccd1 vccd1
+ _12455_/X sky130_fd_sc_hd__o221a_1
X_11406_ _11414_/A _11437_/A _11414_/C _11414_/D _13251_/A vssd1 vssd1 vccd1 vccd1
+ _11407_/B sky130_fd_sc_hd__a41o_1
X_15174_ _15275_/CLK _15174_/D vssd1 vssd1 vccd1 vccd1 _15174_/Q sky130_fd_sc_hd__dfxtp_1
X_12386_ _12379_/X _12381_/X _12383_/X _12385_/X _08405_/C vssd1 vssd1 vccd1 vccd1
+ _12386_/X sky130_fd_sc_hd__o221a_1
XFILLER_125_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14125_ _15675_/CLK _14125_/D vssd1 vssd1 vccd1 vccd1 _14125_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11337_ _11053_/S _11324_/Y _11336_/Y _11307_/A vssd1 vssd1 vccd1 vccd1 _11337_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_181_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14056_ _15334_/CLK _14056_/D vssd1 vssd1 vccd1 vccd1 _14056_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_5_30_0_clk clkbuf_5_31_0_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_5_30_0_clk/X
+ sky130_fd_sc_hd__clkbuf_8
X_11268_ _11283_/A _11323_/B vssd1 vssd1 vccd1 vccd1 _11268_/Y sky130_fd_sc_hd__nand2_1
XFILLER_79_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13007_ _15482_/Q _13093_/A2 _13116_/C _13006_/X vssd1 vssd1 vccd1 vccd1 _15482_/D
+ sky130_fd_sc_hd__a22o_1
X_10219_ input14/X _08487_/A _13282_/S vssd1 vssd1 vccd1 vccd1 _14604_/D sky130_fd_sc_hd__mux2_1
X_11199_ _11199_/A _11199_/B vssd1 vssd1 vccd1 vccd1 _11199_/Y sky130_fd_sc_hd__nor2_1
XFILLER_95_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14958_ _15021_/CLK _14958_/D vssd1 vssd1 vccd1 vccd1 _14958_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_94_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13909_ _15523_/CLK _13909_/D vssd1 vssd1 vccd1 vccd1 _13909_/Q sky130_fd_sc_hd__dfxtp_1
X_14889_ _15644_/CLK _14889_/D vssd1 vssd1 vccd1 vccd1 _14889_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07430_ _14659_/Q _07474_/B _07482_/C vssd1 vssd1 vccd1 vccd1 _07430_/X sky130_fd_sc_hd__and3_1
XFILLER_23_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_572 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07361_ _07352_/A _07352_/B _07331_/Y _07332_/X _07344_/X vssd1 vssd1 vccd1 vccd1
+ _07362_/B sky130_fd_sc_hd__o221a_1
XFILLER_188_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09100_ _15283_/Q _15251_/Q _15219_/Q _15150_/Q _09444_/S _09446_/A1 vssd1 vssd1
+ vccd1 vccd1 _09100_/X sky130_fd_sc_hd__mux4_1
X_07292_ _07292_/A _07292_/B vssd1 vssd1 vccd1 vccd1 _07348_/A sky130_fd_sc_hd__nor2_1
XFILLER_30_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09031_ _15114_/Q _15082_/Q _15655_/Q _13389_/Q _09521_/S _09523_/A1 vssd1 vssd1
+ vccd1 vccd1 _09031_/X sky130_fd_sc_hd__mux4_1
XFILLER_175_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09933_ _13320_/A0 _14293_/Q _09963_/S vssd1 vssd1 vccd1 vccd1 _14293_/D sky130_fd_sc_hd__mux2_1
XTAP_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09864_ _08817_/Y _11743_/C _13318_/C vssd1 vssd1 vccd1 vccd1 _09964_/B sky130_fd_sc_hd__and3b_4
XFILLER_100_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08815_ _11816_/A1 _13841_/Q _08816_/S vssd1 vssd1 vccd1 vccd1 _13841_/D sky130_fd_sc_hd__mux2_1
XTAP_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_856 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09795_ _14162_/Q _11883_/A1 _09795_/S vssd1 vssd1 vccd1 vccd1 _14162_/D sky130_fd_sc_hd__mux2_1
XFILLER_100_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08746_ _13445_/Q _08746_/A2 _08523_/Y _13644_/Q vssd1 vssd1 vccd1 vccd1 _08746_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_2506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08677_ _13519_/Q _08683_/A2 _08685_/A2 _13551_/Q _08676_/X vssd1 vssd1 vccd1 vccd1
+ _08681_/B sky130_fd_sc_hd__a221o_1
XTAP_1805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07628_ _13469_/Q _07655_/A vssd1 vssd1 vccd1 vccd1 _07629_/B sky130_fd_sc_hd__xnor2_1
XTAP_1838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07559_ _13451_/Q _13450_/Q _13449_/Q _07559_/D vssd1 vssd1 vccd1 vccd1 _07576_/C
+ sky130_fd_sc_hd__and4_4
XFILLER_50_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10570_ _15026_/Q _14731_/Q _14927_/Q vssd1 vssd1 vccd1 vccd1 _10570_/X sky130_fd_sc_hd__mux2_1
XFILLER_10_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09229_ _09234_/S1 _09227_/X _09228_/X vssd1 vssd1 vccd1 vccd1 _09229_/X sky130_fd_sc_hd__a21o_1
XFILLER_181_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12240_ _13954_/Q _13696_/Q _12246_/S vssd1 vssd1 vccd1 vccd1 _12241_/B sky130_fd_sc_hd__mux2_1
XFILLER_5_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_256_clk clkbuf_5_0_0_clk/X vssd1 vssd1 vccd1 vccd1 _15176_/CLK sky130_fd_sc_hd__clkbuf_16
X_12171_ _13951_/Q _13693_/Q _12246_/S vssd1 vssd1 vccd1 vccd1 _12172_/B sky130_fd_sc_hd__mux2_1
XFILLER_150_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11122_ _11076_/X _11080_/X _11252_/A vssd1 vssd1 vccd1 vccd1 _11122_/X sky130_fd_sc_hd__mux2_1
XFILLER_174_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11053_ _10955_/B _10963_/Y _11053_/S vssd1 vssd1 vccd1 vccd1 _11053_/X sky130_fd_sc_hd__mux2_1
XFILLER_77_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10004_ _13325_/A0 _14362_/Q _10029_/S vssd1 vssd1 vccd1 vccd1 _14362_/D sky130_fd_sc_hd__mux2_1
XFILLER_114_1024 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14812_ _15630_/CLK _14812_/D vssd1 vssd1 vccd1 vccd1 _14812_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_208 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14743_ _15592_/CLK _14743_/D vssd1 vssd1 vccd1 vccd1 _14743_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_91_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11955_ _14457_/Q _14425_/Q _13846_/Q _14199_/Q _12079_/S _12268_/A vssd1 vssd1 vccd1
+ vccd1 _11955_/X sky130_fd_sc_hd__mux4_1
XFILLER_45_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10906_ _11414_/C _10951_/B vssd1 vssd1 vccd1 vccd1 _10906_/Y sky130_fd_sc_hd__nand2_1
XFILLER_178_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14674_ _15645_/CLK _14674_/D vssd1 vssd1 vccd1 vccd1 _14674_/Q sky130_fd_sc_hd__dfxtp_1
X_11886_ _14454_/Q _14422_/Q _13843_/Q _14196_/Q _12154_/S _12253_/S1 vssd1 vssd1
+ vccd1 vccd1 _11886_/X sky130_fd_sc_hd__mux4_1
XFILLER_32_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13625_ _15379_/CLK _13625_/D vssd1 vssd1 vccd1 vccd1 _13625_/Q sky130_fd_sc_hd__dfxtp_1
X_10837_ _14869_/Q _13799_/Q _12906_/S vssd1 vssd1 vccd1 vccd1 _14869_/D sky130_fd_sc_hd__mux2_1
XFILLER_158_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13556_ _13627_/CLK _13556_/D vssd1 vssd1 vccd1 vccd1 _13556_/Q sky130_fd_sc_hd__dfxtp_1
X_10768_ _14800_/Q _15432_/Q _12932_/S vssd1 vssd1 vccd1 vccd1 _14800_/D sky130_fd_sc_hd__mux2_1
XFILLER_12_171 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12507_ _14481_/Q _14449_/Q _13870_/Q _14223_/Q _12522_/S _12521_/A vssd1 vssd1 vccd1
+ vccd1 _12507_/X sky130_fd_sc_hd__mux4_1
XFILLER_160_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13487_ _15377_/CLK _13487_/D vssd1 vssd1 vccd1 vccd1 _13487_/Q sky130_fd_sc_hd__dfxtp_2
X_10699_ _15067_/Q _10714_/A2 _10696_/X _10698_/X vssd1 vssd1 vccd1 vccd1 _10699_/X
+ sky130_fd_sc_hd__o22a_2
XFILLER_8_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15226_ _15226_/CLK _15226_/D vssd1 vssd1 vccd1 vccd1 _15226_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12438_ _14478_/Q _14446_/Q _13867_/Q _14220_/Q _12453_/S _12452_/A vssd1 vssd1 vccd1
+ vccd1 _12438_/X sky130_fd_sc_hd__mux4_1
XFILLER_126_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_247_clk clkbuf_5_4_0_clk/X vssd1 vssd1 vccd1 vccd1 _15285_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_141_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15157_ _15666_/CLK _15157_/D vssd1 vssd1 vccd1 vccd1 _15157_/Q sky130_fd_sc_hd__dfxtp_1
X_12369_ _14475_/Q _14443_/Q _13864_/Q _14217_/Q _12522_/S _12521_/A vssd1 vssd1 vccd1
+ vccd1 _12369_/X sky130_fd_sc_hd__mux4_1
XFILLER_99_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14108_ _15663_/CLK _14108_/D vssd1 vssd1 vccd1 vccd1 _14108_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15088_ _15088_/CLK _15088_/D vssd1 vssd1 vccd1 vccd1 _15088_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14039_ _15108_/CLK _14039_/D vssd1 vssd1 vccd1 vccd1 _14039_/Q sky130_fd_sc_hd__dfxtp_1
X_06930_ _06690_/Y _13475_/Q _06693_/Y _13474_/Q _06884_/X vssd1 vssd1 vccd1 vccd1
+ _06931_/B sky130_fd_sc_hd__o221a_1
XFILLER_67_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06861_ _12647_/B _06861_/B vssd1 vssd1 vccd1 vccd1 _06861_/Y sky130_fd_sc_hd__nor2_8
XFILLER_94_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08600_ _13466_/Q _08684_/A2 _08691_/B1 _13498_/Q vssd1 vssd1 vccd1 vccd1 _08600_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_67_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09580_ _13956_/Q _11761_/A0 _09594_/S vssd1 vssd1 vccd1 vccd1 _13956_/D sky130_fd_sc_hd__mux2_1
XFILLER_67_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06792_ _14589_/Q _08465_/B vssd1 vssd1 vccd1 vccd1 _09829_/B sky130_fd_sc_hd__and2_2
XFILLER_83_859 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08531_ _13125_/B _13125_/A _08531_/C vssd1 vssd1 vccd1 vccd1 _08531_/Y sky130_fd_sc_hd__nor3_2
XFILLER_82_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08462_ _14596_/Q _12878_/S _08773_/B _08461_/X vssd1 vssd1 vccd1 vccd1 _13761_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_23_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07413_ _13328_/A0 _13392_/Q _07481_/S vssd1 vssd1 vccd1 vccd1 _13392_/D sky130_fd_sc_hd__mux2_1
XFILLER_168_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08393_ _14587_/Q _08421_/B vssd1 vssd1 vccd1 vccd1 _08400_/C sky130_fd_sc_hd__nor2_2
XFILLER_177_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07344_ _07322_/X _07324_/Y _07339_/X _07341_/Y vssd1 vssd1 vccd1 vccd1 _07344_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_177_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07275_ _13922_/Q _15509_/Q _07339_/S vssd1 vssd1 vccd1 vccd1 _10360_/A sky130_fd_sc_hd__mux2_4
XFILLER_163_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09014_ _12573_/A _09014_/B _09014_/C vssd1 vssd1 vccd1 vccd1 _09014_/X sky130_fd_sc_hd__and3_4
XFILLER_129_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_238_clk clkbuf_5_5_0_clk/X vssd1 vssd1 vccd1 vccd1 _15244_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_105_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout600 _14599_/Q vssd1 vssd1 vccd1 vccd1 fanout600/X sky130_fd_sc_hd__buf_12
Xfanout611 _08457_/A vssd1 vssd1 vccd1 vccd1 _12470_/S sky130_fd_sc_hd__buf_12
XFILLER_137_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09916_ _11761_/A0 _14277_/Q _09930_/S vssd1 vssd1 vccd1 vccd1 _14277_/D sky130_fd_sc_hd__mux2_1
Xfanout622 _12545_/S vssd1 vssd1 vccd1 vccd1 _12612_/S sky130_fd_sc_hd__buf_12
Xfanout633 _13739_/Q vssd1 vssd1 vccd1 vccd1 _13236_/A sky130_fd_sc_hd__buf_8
Xfanout644 _07965_/C1 vssd1 vssd1 vccd1 vccd1 _08002_/C1 sky130_fd_sc_hd__buf_8
XTAP_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09847_ _14211_/Q _13334_/A0 _09858_/S vssd1 vssd1 vccd1 vccd1 _14211_/D sky130_fd_sc_hd__mux2_1
XFILLER_101_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_964 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09778_ _14145_/Q _13333_/A0 _09790_/S vssd1 vssd1 vccd1 vccd1 _14145_/D sky130_fd_sc_hd__mux2_1
XTAP_3026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08729_ _13583_/Q _08749_/A2 _08538_/Y _15371_/Q vssd1 vssd1 vccd1 vccd1 _08729_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_73_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11740_ _15169_/Q _11881_/A1 _11742_/S vssd1 vssd1 vccd1 vccd1 _15169_/D sky130_fd_sc_hd__mux2_1
XTAP_1624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11671_ _13346_/A0 _15103_/Q _11675_/S vssd1 vssd1 vccd1 vccd1 _15103_/D sky130_fd_sc_hd__mux2_1
XFILLER_168_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13410_ _15676_/CLK _13410_/D vssd1 vssd1 vccd1 vccd1 _13410_/Q sky130_fd_sc_hd__dfxtp_1
X_10622_ _15003_/Q _10717_/A2 _10652_/B _13722_/Q _10717_/C1 vssd1 vssd1 vccd1 vccd1
+ _10622_/X sky130_fd_sc_hd__a221o_1
X_14390_ _15665_/CLK _14390_/D vssd1 vssd1 vccd1 vccd1 _14390_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_168_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13341_ _13341_/A0 _15671_/Q _13345_/S vssd1 vssd1 vccd1 vccd1 _15671_/D sky130_fd_sc_hd__mux2_1
XFILLER_182_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10553_ _11356_/B _13159_/B vssd1 vssd1 vccd1 vccd1 _10554_/B sky130_fd_sc_hd__nand2_1
XFILLER_167_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13272_ _15356_/Q _15603_/Q _13288_/S vssd1 vssd1 vccd1 vccd1 _15603_/D sky130_fd_sc_hd__mux2_1
XFILLER_143_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10484_ _11536_/A _13208_/B vssd1 vssd1 vccd1 vccd1 _10528_/A sky130_fd_sc_hd__xnor2_1
XFILLER_182_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15011_ _15577_/CLK _15011_/D vssd1 vssd1 vccd1 vccd1 _15011_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_229_clk clkbuf_5_6_0_clk/X vssd1 vssd1 vccd1 vccd1 _15233_/CLK sky130_fd_sc_hd__clkbuf_16
X_12223_ _14081_/Q _14049_/Q _12476_/S vssd1 vssd1 vccd1 vccd1 _12223_/X sky130_fd_sc_hd__mux2_1
XFILLER_5_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12154_ _14078_/Q _14046_/Q _12154_/S vssd1 vssd1 vccd1 vccd1 _12154_/X sky130_fd_sc_hd__mux2_1
XFILLER_78_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11105_ _11129_/A _11105_/B vssd1 vssd1 vccd1 vccd1 _11105_/X sky130_fd_sc_hd__or2_1
XFILLER_151_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12085_ _14075_/Q _14043_/Q _12269_/S vssd1 vssd1 vccd1 vccd1 _12085_/X sky130_fd_sc_hd__mux2_1
XFILLER_1_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11036_ _11036_/A _11036_/B vssd1 vssd1 vccd1 vccd1 _11036_/Y sky130_fd_sc_hd__nor2_1
XFILLER_103_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12987_ _10649_/X _14876_/Q _13029_/S vssd1 vssd1 vccd1 vccd1 _12987_/X sky130_fd_sc_hd__mux2_8
XTAP_3560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14726_ _15552_/CLK _14726_/D vssd1 vssd1 vccd1 vccd1 _14726_/Q sky130_fd_sc_hd__dfxtp_1
X_11938_ _12536_/A _11938_/B vssd1 vssd1 vccd1 vccd1 _11938_/X sky130_fd_sc_hd__or2_1
XFILLER_17_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14657_ _15628_/CLK _14657_/D vssd1 vssd1 vccd1 vccd1 _14657_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_178_739 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11869_ _15290_/Q _13336_/A0 _11883_/S vssd1 vssd1 vccd1 vccd1 _15290_/D sky130_fd_sc_hd__mux2_1
XFILLER_159_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13608_ _15375_/CLK _13608_/D vssd1 vssd1 vccd1 vccd1 _13608_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_159_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14588_ _14612_/CLK _14588_/D vssd1 vssd1 vccd1 vccd1 _14588_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_159_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13539_ _13642_/CLK _13539_/D vssd1 vssd1 vccd1 vccd1 _13539_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_71_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07060_ _14632_/Q _14664_/Q _07078_/S vssd1 vssd1 vccd1 vccd1 _07060_/X sky130_fd_sc_hd__mux2_1
XFILLER_145_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15209_ _15209_/CLK _15209_/D vssd1 vssd1 vccd1 vccd1 _15209_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07962_ _13555_/Q _07961_/C _07961_/D _13556_/Q vssd1 vssd1 vccd1 vccd1 _07963_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_87_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09701_ _11681_/A0 _14071_/Q _09723_/S vssd1 vssd1 vccd1 vccd1 _14071_/D sky130_fd_sc_hd__mux2_1
X_06913_ _07621_/A _15390_/Q _13468_/Q _06918_/A vssd1 vssd1 vccd1 vccd1 _06920_/A
+ sky130_fd_sc_hd__a2bb2o_1
X_07893_ _07900_/C _07900_/D vssd1 vssd1 vccd1 vccd1 _07897_/B sky130_fd_sc_hd__nand2_1
XFILLER_114_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09632_ _14005_/Q _11854_/A1 _09661_/S vssd1 vssd1 vccd1 vccd1 _14005_/D sky130_fd_sc_hd__mux2_1
XFILLER_55_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06844_ _08405_/B _06680_/Y _06842_/X _06843_/Y vssd1 vssd1 vccd1 vccd1 _06844_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_56_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09563_ _13939_/Q _13319_/A0 _09589_/S vssd1 vssd1 vccd1 vccd1 _13939_/D sky130_fd_sc_hd__mux2_1
XFILLER_55_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06775_ _14924_/Q _06775_/B _10561_/C vssd1 vssd1 vccd1 vccd1 _06775_/Y sky130_fd_sc_hd__nor3_2
XFILLER_167_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08514_ _13444_/Q _08736_/A2 _08748_/B1 _14517_/Q vssd1 vssd1 vccd1 vccd1 _08514_/X
+ sky130_fd_sc_hd__a22o_1
X_09494_ _13935_/Q _09493_/X _12573_/A vssd1 vssd1 vccd1 vccd1 _13935_/D sky130_fd_sc_hd__mux2_1
XFILLER_23_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08445_ _08487_/A _08390_/C _08425_/X _10764_/S vssd1 vssd1 vccd1 vccd1 _08445_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_168_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08376_ _08355_/Y _08375_/Y _11259_/S vssd1 vssd1 vccd1 vccd1 _08376_/X sky130_fd_sc_hd__mux2_1
XFILLER_177_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07327_ _07327_/A vssd1 vssd1 vccd1 vccd1 _07327_/Y sky130_fd_sc_hd__inv_2
XFILLER_176_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07258_ _07258_/A vssd1 vssd1 vccd1 vccd1 _07258_/Y sky130_fd_sc_hd__inv_2
XFILLER_164_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07189_ _15363_/Q _15070_/Q _07193_/S vssd1 vssd1 vccd1 vccd1 _07189_/X sky130_fd_sc_hd__mux2_2
XFILLER_3_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout430 _08497_/A vssd1 vssd1 vccd1 vccd1 _08519_/B sky130_fd_sc_hd__buf_12
Xfanout441 _07500_/S vssd1 vssd1 vccd1 vccd1 _07480_/S sky130_fd_sc_hd__buf_12
XFILLER_87_940 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout452 _10630_/S vssd1 vssd1 vccd1 vccd1 _10695_/S sky130_fd_sc_hd__buf_8
Xfanout463 _06675_/Y vssd1 vssd1 vccd1 vccd1 _09437_/A1 sky130_fd_sc_hd__buf_12
Xfanout474 _12548_/S vssd1 vssd1 vccd1 vccd1 _12168_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_58_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout485 _06669_/Y vssd1 vssd1 vccd1 vccd1 _12615_/A1 sky130_fd_sc_hd__buf_12
X_12910_ _15438_/Q _15624_/Q _12910_/S vssd1 vssd1 vccd1 vccd1 _15438_/D sky130_fd_sc_hd__mux2_1
XFILLER_19_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout496 _08145_/S vssd1 vssd1 vccd1 vccd1 _08133_/S sky130_fd_sc_hd__buf_8
XFILLER_111_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13890_ _15088_/CLK _13890_/D vssd1 vssd1 vccd1 vccd1 _13890_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12841_ _14735_/Q _15369_/Q _12871_/S vssd1 vssd1 vccd1 vccd1 _15369_/D sky130_fd_sc_hd__mux2_1
XTAP_2111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15560_ _15587_/CLK _15560_/D vssd1 vssd1 vccd1 vccd1 _15560_/Q sky130_fd_sc_hd__dfxtp_1
X_12772_ _13435_/Q _12647_/B _08030_/Y _13602_/Q _12743_/A vssd1 vssd1 vccd1 vccd1
+ _12772_/X sky130_fd_sc_hd__a221o_1
XTAP_2155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14511_ _14511_/CLK _14511_/D vssd1 vssd1 vccd1 vccd1 _14511_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11723_ _15152_/Q _13331_/A0 _11741_/S vssd1 vssd1 vccd1 vccd1 _15152_/D sky130_fd_sc_hd__mux2_1
XTAP_1454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15491_ _15499_/CLK _15491_/D vssd1 vssd1 vccd1 vccd1 _15491_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14442_ _15669_/CLK _14442_/D vssd1 vssd1 vccd1 vccd1 _14442_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11654_ _13329_/A0 _15086_/Q _11670_/S vssd1 vssd1 vccd1 vccd1 _15086_/D sky130_fd_sc_hd__mux2_1
XFILLER_174_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10605_ _14739_/Q _10604_/X _10730_/S vssd1 vssd1 vccd1 vccd1 _14739_/D sky130_fd_sc_hd__mux2_1
X_14373_ _14373_/CLK _14373_/D vssd1 vssd1 vccd1 vccd1 _14373_/Q sky130_fd_sc_hd__dfxtp_1
X_11585_ _11585_/A _11585_/B vssd1 vssd1 vccd1 vccd1 _11586_/B sky130_fd_sc_hd__nor2_2
XFILLER_127_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13324_ _13324_/A0 _15654_/Q _13350_/S vssd1 vssd1 vccd1 vccd1 _15654_/D sky130_fd_sc_hd__mux2_1
XFILLER_6_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10536_ _11616_/A _13242_/B _10534_/X _10535_/X _10442_/Y vssd1 vssd1 vccd1 vccd1
+ _10537_/C sky130_fd_sc_hd__o221a_1
XFILLER_171_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13255_ _15339_/Q _15586_/Q _13291_/S vssd1 vssd1 vccd1 vccd1 _15586_/D sky130_fd_sc_hd__mux2_1
X_10467_ _13233_/B _11598_/A vssd1 vssd1 vccd1 vccd1 _10532_/A sky130_fd_sc_hd__and2b_1
XFILLER_6_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12206_ _15319_/Q _13105_/A2 _12205_/X vssd1 vssd1 vccd1 vccd1 _15319_/D sky130_fd_sc_hd__a21o_1
XFILLER_124_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13186_ _13229_/A _11440_/A _11476_/B vssd1 vssd1 vccd1 vccd1 _13186_/Y sky130_fd_sc_hd__a21oi_1
X_10398_ _11399_/A _11414_/C vssd1 vssd1 vccd1 vccd1 _10399_/B sky130_fd_sc_hd__xnor2_1
XFILLER_2_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12137_ _15316_/Q _13105_/A2 _12136_/X vssd1 vssd1 vccd1 vccd1 _15316_/D sky130_fd_sc_hd__a21o_1
XFILLER_123_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12068_ _15313_/Q _13081_/A2 _12067_/X vssd1 vssd1 vccd1 vccd1 _15313_/D sky130_fd_sc_hd__a21o_1
XFILLER_49_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11019_ _11025_/A _13208_/B vssd1 vssd1 vccd1 vccd1 _11249_/A sky130_fd_sc_hd__and2_1
XTAP_4080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14709_ _15615_/CLK _14709_/D vssd1 vssd1 vccd1 vccd1 _14709_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_20_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08230_ _07322_/X _10457_/A2 _08229_/X vssd1 vssd1 vccd1 vccd1 _08230_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_60_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08161_ _08185_/A _08161_/B vssd1 vssd1 vccd1 vccd1 _08161_/X sky130_fd_sc_hd__and2_1
XFILLER_174_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07112_ _14834_/Q _07115_/B _07163_/A vssd1 vssd1 vccd1 vccd1 _07112_/X sky130_fd_sc_hd__and3_2
XFILLER_174_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08092_ input8/X input17/X _08145_/S vssd1 vssd1 vccd1 vccd1 _08154_/B sky130_fd_sc_hd__mux2_1
XFILLER_162_904 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_978 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07043_ _07042_/X _13593_/Q _12728_/S vssd1 vssd1 vccd1 vccd1 _07043_/X sky130_fd_sc_hd__mux2_1
XFILLER_146_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08994_ _09532_/A _08994_/B vssd1 vssd1 vccd1 vccd1 _08994_/X sky130_fd_sc_hd__or2_1
XFILLER_87_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_558 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07945_ _14744_/Q _07964_/A _07944_/Y vssd1 vssd1 vccd1 vccd1 _13551_/D sky130_fd_sc_hd__o21a_1
XFILLER_69_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07876_ _13534_/Q _13533_/Q vssd1 vssd1 vccd1 vccd1 _07884_/D sky130_fd_sc_hd__and2_1
XFILLER_141_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09615_ _13989_/Q _13337_/A0 _09628_/S vssd1 vssd1 vccd1 vccd1 _13989_/D sky130_fd_sc_hd__mux2_1
X_06827_ _14730_/Q _12640_/S vssd1 vssd1 vccd1 vccd1 _08817_/B sky130_fd_sc_hd__and2_4
XFILLER_43_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09546_ _14259_/Q _14291_/Q _14323_/Q _14355_/Q _09469_/S _09546_/S1 vssd1 vssd1
+ vccd1 vccd1 _09546_/X sky130_fd_sc_hd__mux4_1
X_06758_ _13738_/Q vssd1 vssd1 vccd1 vccd1 _06758_/Y sky130_fd_sc_hd__inv_2
XFILLER_36_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09477_ _13123_/A _09474_/X _09476_/X _09554_/A vssd1 vssd1 vccd1 vccd1 _09477_/X
+ sky130_fd_sc_hd__o211a_1
X_06689_ _14516_/Q vssd1 vssd1 vccd1 vccd1 _06874_/A sky130_fd_sc_hd__inv_2
XFILLER_24_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08428_ _13744_/Q _12906_/S _08426_/B _08427_/X vssd1 vssd1 vccd1 vccd1 _13744_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_141_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08359_ _08282_/X _08358_/X _11329_/A vssd1 vssd1 vccd1 vccd1 _08359_/X sky130_fd_sc_hd__mux2_2
XFILLER_177_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11370_ _15045_/Q _11641_/S _11369_/X vssd1 vssd1 vccd1 vccd1 _15045_/D sky130_fd_sc_hd__a21bo_1
XFILLER_180_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_263 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10321_ _14706_/Q _14891_/Q _10730_/S vssd1 vssd1 vccd1 vccd1 _14706_/D sky130_fd_sc_hd__mux2_1
XFILLER_30_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13040_ _15493_/Q _10892_/B _13116_/C _13039_/X vssd1 vssd1 vccd1 vccd1 _15493_/D
+ sky130_fd_sc_hd__a22o_1
X_10252_ _14637_/Q _14790_/Q _10710_/S vssd1 vssd1 vccd1 vccd1 _14637_/D sky130_fd_sc_hd__mux2_1
XFILLER_1_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10183_ _11761_/A0 _14567_/Q _10197_/S vssd1 vssd1 vccd1 vccd1 _14567_/D sky130_fd_sc_hd__mux2_1
XFILLER_105_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14991_ _15582_/CLK _14991_/D vssd1 vssd1 vccd1 vccd1 _14991_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout260 _07370_/X vssd1 vssd1 vccd1 vccd1 _07501_/S sky130_fd_sc_hd__buf_12
Xfanout271 _08510_/X vssd1 vssd1 vccd1 vccd1 _08736_/A2 sky130_fd_sc_hd__buf_12
XFILLER_8_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout282 _11883_/A1 vssd1 vssd1 vccd1 vccd1 _13350_/A0 sky130_fd_sc_hd__buf_6
XFILLER_75_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13942_ _15202_/CLK _13942_/D vssd1 vssd1 vccd1 vccd1 _13942_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout293 _13104_/B2 vssd1 vssd1 vccd1 vccd1 _13345_/A0 sky130_fd_sc_hd__buf_6
XFILLER_115_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13873_ _14420_/CLK _13873_/D vssd1 vssd1 vccd1 vccd1 _13873_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15612_ _15612_/CLK _15612_/D vssd1 vssd1 vccd1 vccd1 _15612_/Q sky130_fd_sc_hd__dfxtp_1
X_12824_ _06861_/Y _12821_/X _12822_/X _12823_/X vssd1 vssd1 vccd1 vccd1 _12824_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_61_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15543_ _15543_/CLK _15543_/D vssd1 vssd1 vccd1 vccd1 _15543_/Q sky130_fd_sc_hd__dfxtp_1
X_12755_ _12767_/C _12755_/B vssd1 vssd1 vccd1 vccd1 _12755_/X sky130_fd_sc_hd__and2b_1
XTAP_1240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11706_ _11881_/A1 _15137_/Q _11708_/S vssd1 vssd1 vccd1 vccd1 _15137_/D sky130_fd_sc_hd__mux2_1
XTAP_1284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15474_ _15501_/CLK _15474_/D vssd1 vssd1 vccd1 vccd1 _15474_/Q sky130_fd_sc_hd__dfxtp_1
X_12686_ _15346_/Q _12765_/B _12685_/X _12809_/C1 vssd1 vssd1 vccd1 vccd1 _15346_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_1295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14425_ _15244_/CLK _14425_/D vssd1 vssd1 vccd1 vccd1 _14425_/Q sky130_fd_sc_hd__dfxtp_1
X_11637_ _11633_/A _11633_/B _11635_/A _11635_/B vssd1 vssd1 vccd1 vccd1 _11640_/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_30_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14356_ _15172_/CLK _14356_/D vssd1 vssd1 vccd1 vccd1 _14356_/Q sky130_fd_sc_hd__dfxtp_1
X_11568_ _11567_/X _15065_/Q _11614_/S vssd1 vssd1 vccd1 vccd1 _15065_/D sky130_fd_sc_hd__mux2_1
XFILLER_183_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13307_ _15639_/Q _12778_/B _13316_/S vssd1 vssd1 vccd1 vccd1 _15639_/D sky130_fd_sc_hd__mux2_1
XFILLER_155_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10519_ _10519_/A _10519_/B vssd1 vssd1 vccd1 vccd1 _10528_/D sky130_fd_sc_hd__or2_1
XFILLER_155_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14287_ _15199_/CLK _14287_/D vssd1 vssd1 vccd1 vccd1 _14287_/Q sky130_fd_sc_hd__dfxtp_1
X_11499_ _11500_/A _11500_/B vssd1 vssd1 vccd1 vccd1 _11501_/A sky130_fd_sc_hd__nand2_1
X_13238_ _13236_/Y _13237_/X _15579_/Q _13214_/B vssd1 vssd1 vccd1 vccd1 _15579_/D
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_130_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13169_ _13251_/A _13168_/B _13219_/S _11380_/A vssd1 vssd1 vccd1 vccd1 _13169_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_34_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_355 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07730_ _13495_/Q _07727_/B _13496_/Q vssd1 vssd1 vccd1 vccd1 _07730_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_38_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07661_ _13477_/Q _07665_/C vssd1 vssd1 vccd1 vccd1 _07662_/B sky130_fd_sc_hd__xnor2_1
XFILLER_19_870 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09400_ _13899_/Q _09445_/A2 _09522_/B1 _14414_/Q _09445_/C1 vssd1 vssd1 vccd1 vccd1
+ _09400_/X sky130_fd_sc_hd__a221o_1
X_07592_ _07607_/A _07592_/B vssd1 vssd1 vccd1 vccd1 _07592_/Y sky130_fd_sc_hd__nand2_1
X_09331_ _14443_/Q _08540_/B _13130_/C1 _09330_/X vssd1 vssd1 vccd1 vccd1 _09331_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_34_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09262_ _15291_/Q _15259_/Q _15227_/Q _15158_/Q _09484_/S _09550_/A1 vssd1 vssd1
+ vccd1 vccd1 _09262_/X sky130_fd_sc_hd__mux4_1
XFILLER_138_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08213_ _13704_/Q _13342_/A0 _08221_/S vssd1 vssd1 vccd1 vccd1 _13704_/D sky130_fd_sc_hd__mux2_1
XFILLER_178_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09193_ _15122_/Q _15090_/Q _15663_/Q _13397_/Q _09190_/S _09429_/S1 vssd1 vssd1
+ vccd1 vccd1 _09193_/X sky130_fd_sc_hd__mux4_1
XFILLER_140_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08144_ _13662_/Q _10610_/S _08119_/X _08143_/X vssd1 vssd1 vccd1 vccd1 _13662_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_162_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08075_ _08078_/B _08075_/B _08083_/A vssd1 vssd1 vccd1 vccd1 _08075_/X sky130_fd_sc_hd__or3b_1
XFILLER_161_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07026_ _07025_/X _14741_/Q _07098_/S vssd1 vssd1 vccd1 vccd1 _13587_/D sky130_fd_sc_hd__mux2_1
XFILLER_136_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08977_ _14458_/Q _14426_/Q _13847_/Q _14200_/Q _09225_/S0 _09225_/S1 vssd1 vssd1
+ vccd1 vccd1 _08977_/X sky130_fd_sc_hd__mux4_1
XFILLER_29_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07928_ _13547_/Q _07935_/D vssd1 vssd1 vccd1 vccd1 _07932_/B sky130_fd_sc_hd__nand2_1
XFILLER_29_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07859_ _13528_/Q _13527_/Q _07858_/D _13529_/Q vssd1 vssd1 vccd1 vccd1 _07859_/Y
+ sky130_fd_sc_hd__a31oi_1
XFILLER_16_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_23 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10870_ _14902_/Q _13736_/Q _12904_/S vssd1 vssd1 vccd1 vccd1 _14902_/D sky130_fd_sc_hd__mux2_1
XPHY_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09529_ _08668_/D _09525_/X _09528_/X _09524_/X vssd1 vssd1 vccd1 vccd1 _09539_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_43_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12540_ _12540_/A _12540_/B vssd1 vssd1 vccd1 vccd1 _12540_/X sky130_fd_sc_hd__and2_1
XFILLER_24_383 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12471_ _12498_/A _12471_/B vssd1 vssd1 vccd1 vccd1 _12471_/X sky130_fd_sc_hd__and2_1
XFILLER_12_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_336 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14210_ _14468_/CLK _14210_/D vssd1 vssd1 vccd1 vccd1 _14210_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_99 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11422_ _11404_/A _11402_/Y _11423_/D _11421_/X _11410_/B vssd1 vssd1 vccd1 vccd1
+ _11422_/X sky130_fd_sc_hd__a32o_2
XFILLER_172_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15190_ _15291_/CLK _15190_/D vssd1 vssd1 vccd1 vccd1 _15190_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_165_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14141_ _15674_/CLK _14141_/D vssd1 vssd1 vccd1 vccd1 _14141_/Q sky130_fd_sc_hd__dfxtp_1
X_11353_ _08388_/X _11303_/A _11352_/Y vssd1 vssd1 vccd1 vccd1 _15042_/D sky130_fd_sc_hd__o21ai_1
XFILLER_165_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10304_ _14689_/Q _14874_/Q _10650_/S vssd1 vssd1 vccd1 vccd1 _14689_/D sky130_fd_sc_hd__mux2_1
X_14072_ _15295_/CLK _14072_/D vssd1 vssd1 vccd1 vccd1 _14072_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_141_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_243 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11284_ _11347_/A _11282_/X _11283_/X _08233_/B vssd1 vssd1 vccd1 vccd1 _11284_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_180_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_108 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13023_ _10709_/X _14888_/Q _13029_/S vssd1 vssd1 vccd1 vccd1 _13023_/X sky130_fd_sc_hd__mux2_4
X_10235_ _14620_/Q _14773_/Q _10343_/S vssd1 vssd1 vccd1 vccd1 _14620_/D sky130_fd_sc_hd__mux2_1
XFILLER_134_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10166_ _11852_/A1 _14550_/Q _10192_/S vssd1 vssd1 vccd1 vccd1 _14550_/D sky130_fd_sc_hd__mux2_1
XFILLER_86_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14974_ _14988_/CLK _14974_/D vssd1 vssd1 vccd1 vccd1 _14974_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10097_ _14453_/Q _11883_/A1 _10097_/S vssd1 vssd1 vccd1 vccd1 _14453_/D sky130_fd_sc_hd__mux2_1
X_13925_ _14439_/CLK _13925_/D vssd1 vssd1 vccd1 vccd1 _13925_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_90_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13856_ _15235_/CLK _13856_/D vssd1 vssd1 vccd1 vccd1 _13856_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12807_ _13440_/Q _12647_/B _08030_/Y _13607_/Q _12743_/A vssd1 vssd1 vccd1 vccd1
+ _12807_/X sky130_fd_sc_hd__a221o_2
XFILLER_90_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13787_ _15389_/CLK _13787_/D vssd1 vssd1 vccd1 vccd1 _13787_/Q sky130_fd_sc_hd__dfxtp_4
X_10999_ _10999_/A _10999_/B vssd1 vssd1 vccd1 vccd1 _10999_/Y sky130_fd_sc_hd__nor2_1
X_12738_ _15353_/Q _12765_/B _12737_/X _12809_/C1 vssd1 vssd1 vccd1 vccd1 _15353_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15526_ _15526_/CLK _15526_/D vssd1 vssd1 vccd1 vccd1 _15526_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_176_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15457_ _15643_/CLK _15457_/D vssd1 vssd1 vccd1 vccd1 _15457_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_175_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12669_ _13588_/Q _12668_/X _12763_/S vssd1 vssd1 vccd1 vccd1 _12669_/X sky130_fd_sc_hd__mux2_1
X_14408_ _15094_/CLK _14408_/D vssd1 vssd1 vccd1 vccd1 _14408_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15388_ _15389_/CLK _15388_/D vssd1 vssd1 vccd1 vccd1 _15388_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_571 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14339_ _15306_/CLK _14339_/D vssd1 vssd1 vccd1 vccd1 _14339_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_143_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08900_ _14518_/Q _14131_/Q _14163_/Q _14099_/Q _09132_/S _08988_/A1 vssd1 vssd1
+ vccd1 vccd1 _08900_/X sky130_fd_sc_hd__mux4_1
XFILLER_143_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09880_ _13080_/B2 _14242_/Q _09892_/S vssd1 vssd1 vccd1 vccd1 _14242_/D sky130_fd_sc_hd__mux2_1
XTAP_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08831_ _13854_/Q _13330_/A0 _08846_/S vssd1 vssd1 vccd1 vccd1 _13854_/D sky130_fd_sc_hd__mux2_1
XTAP_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08762_ _14597_/Q _08756_/B _08410_/Y _14596_/Q _14613_/Q vssd1 vssd1 vccd1 vccd1
+ _08762_/X sky130_fd_sc_hd__o221a_1
XFILLER_39_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07713_ _07713_/A _07713_/B vssd1 vssd1 vccd1 vccd1 _07713_/Y sky130_fd_sc_hd__nand2_1
XFILLER_72_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08693_ _14494_/Q _08693_/A2 _08693_/B1 _13620_/Q _08690_/X vssd1 vssd1 vccd1 vccd1
+ _08693_/X sky130_fd_sc_hd__a221o_1
XFILLER_38_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07644_ _07644_/A _07644_/B vssd1 vssd1 vccd1 vccd1 _07644_/Y sky130_fd_sc_hd__nand2_1
XFILLER_65_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07575_ _13455_/Q _07575_/B vssd1 vssd1 vccd1 vccd1 _07575_/Y sky130_fd_sc_hd__nor2_1
XFILLER_25_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09314_ _14023_/Q _13991_/Q _09481_/S vssd1 vssd1 vccd1 vccd1 _09314_/X sky130_fd_sc_hd__mux2_1
XFILLER_22_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09245_ _08510_/B _09243_/X _09244_/X _08519_/B _13049_/A1 vssd1 vssd1 vccd1 vccd1
+ _09245_/X sky130_fd_sc_hd__a221o_1
X_09176_ _15121_/Q _09536_/A2 _13130_/B1 _15089_/Q _09175_/X vssd1 vssd1 vccd1 vccd1
+ _09176_/X sky130_fd_sc_hd__a221o_1
XFILLER_182_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08127_ _08093_/B _08125_/X _08126_/Y _08121_/X vssd1 vssd1 vccd1 vccd1 _08127_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_147_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08058_ _14751_/Q _13629_/Q _08066_/S vssd1 vssd1 vccd1 vccd1 _13629_/D sky130_fd_sc_hd__mux2_1
XFILLER_135_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput36 _07172_/X vssd1 vssd1 vccd1 vccd1 ext_address[10] sky130_fd_sc_hd__clkbuf_2
XFILLER_1_714 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput47 _07183_/X vssd1 vssd1 vccd1 vccd1 ext_address[21] sky130_fd_sc_hd__clkbuf_2
X_07009_ _14615_/Q _14647_/Q _07096_/S vssd1 vssd1 vccd1 vccd1 _07009_/X sky130_fd_sc_hd__mux2_1
Xoutput58 _07193_/X vssd1 vssd1 vccd1 vccd1 ext_address[31] sky130_fd_sc_hd__clkbuf_2
XFILLER_122_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput69 _07123_/X vssd1 vssd1 vccd1 vccd1 ext_write_data[11] sky130_fd_sc_hd__clkbuf_2
XFILLER_62_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10020_ _11874_/A1 _14378_/Q _10029_/S vssd1 vssd1 vccd1 vccd1 _14378_/D sky130_fd_sc_hd__mux2_1
XFILLER_163_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11971_ _12500_/A1 _11970_/X _12468_/A1 vssd1 vssd1 vccd1 vccd1 _11971_/X sky130_fd_sc_hd__a21o_1
XFILLER_17_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13710_ _15651_/CLK _13710_/D vssd1 vssd1 vccd1 vccd1 _13710_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_1083 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10922_ _14944_/Q _10356_/A _10944_/B vssd1 vssd1 vccd1 vccd1 _14944_/D sky130_fd_sc_hd__mux2_1
XTAP_3978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14690_ _15608_/CLK _14690_/D vssd1 vssd1 vccd1 vccd1 _14690_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13641_ _15397_/CLK _13641_/D vssd1 vssd1 vccd1 vccd1 _13641_/Q sky130_fd_sc_hd__dfxtp_1
X_10853_ _14885_/Q _13783_/Q _12927_/S vssd1 vssd1 vccd1 vccd1 _14885_/D sky130_fd_sc_hd__mux2_1
XFILLER_112_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13572_ _13642_/CLK _13572_/D vssd1 vssd1 vccd1 vccd1 _13572_/Q sky130_fd_sc_hd__dfxtp_1
X_10784_ _14816_/Q _15448_/Q _12928_/S vssd1 vssd1 vccd1 vccd1 _14816_/D sky130_fd_sc_hd__mux2_1
XFILLER_24_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15311_ _15523_/CLK _15311_/D vssd1 vssd1 vccd1 vccd1 _15311_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12523_ _12615_/A1 _12522_/X _08405_/B vssd1 vssd1 vccd1 vccd1 _12523_/X sky130_fd_sc_hd__a21o_1
XPHY_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15242_ _15676_/CLK _15242_/D vssd1 vssd1 vccd1 vccd1 _15242_/Q sky130_fd_sc_hd__dfxtp_1
X_12454_ _12477_/A1 _12453_/X _12468_/A1 vssd1 vssd1 vccd1 vccd1 _12454_/X sky130_fd_sc_hd__a21o_1
XFILLER_126_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11405_ _11404_/Y _15049_/Q _11641_/S vssd1 vssd1 vccd1 vccd1 _15049_/D sky130_fd_sc_hd__mux2_1
X_15173_ _15650_/CLK _15173_/D vssd1 vssd1 vccd1 vccd1 _15173_/Q sky130_fd_sc_hd__dfxtp_1
X_12385_ _12615_/A1 _12384_/X _12615_/B1 vssd1 vssd1 vccd1 vccd1 _12385_/X sky130_fd_sc_hd__a21o_1
XFILLER_125_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14124_ _15674_/CLK _14124_/D vssd1 vssd1 vccd1 vccd1 _14124_/Q sky130_fd_sc_hd__dfxtp_1
X_11336_ _11007_/B _11013_/X _11053_/S vssd1 vssd1 vccd1 vccd1 _11336_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_154_1019 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14055_ _15292_/CLK _14055_/D vssd1 vssd1 vccd1 vccd1 _14055_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11267_ _08386_/X _11266_/X _11297_/S vssd1 vssd1 vccd1 vccd1 _11323_/B sky130_fd_sc_hd__mux2_1
X_13006_ _13092_/B2 _13039_/A2 _13005_/X _12944_/A vssd1 vssd1 vccd1 vccd1 _13006_/X
+ sky130_fd_sc_hd__a22o_1
X_10218_ input13/X _08910_/S _13291_/S vssd1 vssd1 vccd1 vccd1 _14603_/D sky130_fd_sc_hd__mux2_1
XFILLER_67_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11198_ _14991_/Q _11202_/A _11170_/X _11197_/Y vssd1 vssd1 vccd1 vccd1 _14991_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_121_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10149_ _14534_/Q _13335_/A0 _10159_/S vssd1 vssd1 vccd1 vccd1 _14534_/D sky130_fd_sc_hd__mux2_1
X_14957_ _15580_/CLK _14957_/D vssd1 vssd1 vccd1 vccd1 _14957_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13908_ _15499_/CLK _13908_/D vssd1 vssd1 vccd1 vccd1 _13908_/Q sky130_fd_sc_hd__dfxtp_1
X_14888_ _14888_/CLK _14888_/D vssd1 vssd1 vccd1 vccd1 _14888_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13839_ _15259_/CLK _13839_/D vssd1 vssd1 vccd1 vccd1 _13839_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07360_ _07360_/A _07360_/B _07360_/C _07360_/D vssd1 vssd1 vccd1 vccd1 _07363_/C
+ sky130_fd_sc_hd__or4_1
XFILLER_15_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15509_ _15520_/CLK _15509_/D vssd1 vssd1 vccd1 vccd1 _15509_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_175_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07291_ _15318_/Q _15474_/Q _07340_/S vssd1 vssd1 vccd1 vccd1 _07292_/B sky130_fd_sc_hd__mux2_8
XFILLER_176_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09030_ _09523_/A1 _09028_/X _09029_/X vssd1 vssd1 vccd1 vccd1 _09030_/X sky130_fd_sc_hd__a21o_1
XFILLER_129_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_572 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_891 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09932_ _11852_/A1 _14292_/Q _09958_/S vssd1 vssd1 vccd1 vccd1 _14292_/D sky130_fd_sc_hd__mux2_1
XFILLER_131_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09863_ _14227_/Q _11883_/A1 _09863_/S vssd1 vssd1 vccd1 vccd1 _14227_/D sky130_fd_sc_hd__mux2_1
XFILLER_86_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08814_ _11881_/A1 _13840_/Q _08816_/S vssd1 vssd1 vccd1 vccd1 _13840_/D sky130_fd_sc_hd__mux2_1
XTAP_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09794_ _14161_/Q _13349_/A0 _09795_/S vssd1 vssd1 vccd1 vccd1 _14161_/D sky130_fd_sc_hd__mux2_1
XFILLER_100_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08745_ _13805_/Q _08744_/X _12900_/S vssd1 vssd1 vccd1 vccd1 _13805_/D sky130_fd_sc_hd__mux2_1
XFILLER_26_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08676_ _13455_/Q _08684_/A2 _08691_/B1 _13487_/Q vssd1 vssd1 vccd1 vccd1 _08676_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_38_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07627_ _14757_/Q _07629_/A _07626_/Y _08002_/C1 vssd1 vssd1 vccd1 vccd1 _13468_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_1828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07558_ _14739_/Q _07651_/A _07557_/Y _07938_/C1 vssd1 vssd1 vccd1 vccd1 _13450_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_179_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07489_ _13347_/A0 _13411_/Q _07501_/S vssd1 vssd1 vccd1 vccd1 _13411_/D sky130_fd_sc_hd__mux2_1
XFILLER_107_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09228_ _14083_/Q _09231_/A2 _09403_/B1 _14051_/Q _09391_/A vssd1 vssd1 vccd1 vccd1
+ _09228_/X sky130_fd_sc_hd__a221o_1
XFILLER_42_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09159_ _15286_/Q _15254_/Q _15222_/Q _15153_/Q _09444_/S _09446_/A1 vssd1 vssd1
+ vccd1 vccd1 _09159_/X sky130_fd_sc_hd__mux4_1
XFILLER_107_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12170_ _12503_/A1 _12165_/X _12168_/X _12169_/X _08449_/A vssd1 vssd1 vccd1 vccd1
+ _12182_/B sky130_fd_sc_hd__a221o_1
XFILLER_101_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11121_ _11371_/A _11371_/B vssd1 vssd1 vccd1 vccd1 _11375_/B sky130_fd_sc_hd__nand2_1
XFILLER_89_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11052_ _14963_/Q _11202_/A _11051_/X vssd1 vssd1 vccd1 vccd1 _14963_/D sky130_fd_sc_hd__o21a_1
XFILLER_150_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10003_ _11857_/A1 _14361_/Q _10029_/S vssd1 vssd1 vccd1 vccd1 _14361_/D sky130_fd_sc_hd__mux2_1
XFILLER_27_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14811_ _15446_/CLK _14811_/D vssd1 vssd1 vccd1 vccd1 _14811_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_97_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14742_ _15607_/CLK _14742_/D vssd1 vssd1 vccd1 vccd1 _14742_/Q sky130_fd_sc_hd__dfxtp_4
X_11954_ _14231_/Q _14263_/Q _14295_/Q _14327_/Q _12079_/S _12268_/A vssd1 vssd1 vccd1
+ vccd1 _11954_/X sky130_fd_sc_hd__mux4_1
XTAP_3764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10905_ _14935_/Q _10951_/B _10904_/Y _13171_/B vssd1 vssd1 vccd1 vccd1 _14935_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_44_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14673_ _15644_/CLK _14673_/D vssd1 vssd1 vccd1 vccd1 _14673_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_192_clk clkbuf_5_20_0_clk/X vssd1 vssd1 vccd1 vccd1 _15275_/CLK sky130_fd_sc_hd__clkbuf_16
X_11885_ _14228_/Q _14260_/Q _14292_/Q _14324_/Q _11993_/S _12253_/S1 vssd1 vssd1
+ vccd1 vccd1 _11885_/X sky130_fd_sc_hd__mux4_1
XFILLER_60_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13624_ _15381_/CLK _13624_/D vssd1 vssd1 vccd1 vccd1 _13624_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10836_ _14868_/Q _13800_/Q _12878_/S vssd1 vssd1 vccd1 vccd1 _14868_/D sky130_fd_sc_hd__mux2_1
XFILLER_186_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13555_ _13627_/CLK _13555_/D vssd1 vssd1 vccd1 vccd1 _13555_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_158_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10767_ _15431_/Q _14799_/Q _13129_/A vssd1 vssd1 vccd1 vccd1 _14799_/D sky130_fd_sc_hd__mux2_1
XFILLER_40_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12506_ _14255_/Q _14287_/Q _14319_/Q _14351_/Q _08405_/A _12521_/A vssd1 vssd1 vccd1
+ vccd1 _12506_/X sky130_fd_sc_hd__mux4_1
X_13486_ _14495_/CLK _13486_/D vssd1 vssd1 vccd1 vccd1 _13486_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_12_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_1029 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10698_ _14986_/Q _10733_/A2 _10733_/B1 _14954_/Q _10697_/X vssd1 vssd1 vccd1 vccd1
+ _10698_/X sky130_fd_sc_hd__a221o_1
XFILLER_139_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15225_ _15289_/CLK _15225_/D vssd1 vssd1 vccd1 vccd1 _15225_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_173_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12437_ _14252_/Q _14284_/Q _14316_/Q _14348_/Q _12453_/S _12452_/A vssd1 vssd1 vccd1
+ vccd1 _12437_/X sky130_fd_sc_hd__mux4_1
XFILLER_173_659 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15156_ _15289_/CLK _15156_/D vssd1 vssd1 vccd1 vccd1 _15156_/Q sky130_fd_sc_hd__dfxtp_1
X_12368_ _14249_/Q _14281_/Q _14313_/Q _14345_/Q _12522_/S _12521_/A vssd1 vssd1 vccd1
+ vccd1 _12368_/X sky130_fd_sc_hd__mux4_1
XFILLER_154_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14107_ _15212_/CLK _14107_/D vssd1 vssd1 vccd1 vccd1 _14107_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11319_ _11047_/Y _11288_/X _11318_/X _08249_/Y _11344_/A vssd1 vssd1 vccd1 vccd1
+ _11319_/X sky130_fd_sc_hd__a221o_1
X_15087_ _15660_/CLK _15087_/D vssd1 vssd1 vccd1 vccd1 _15087_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12299_ _14246_/Q _14278_/Q _14310_/Q _14342_/Q _12612_/S _12383_/A vssd1 vssd1 vccd1
+ vccd1 _12299_/X sky130_fd_sc_hd__mux4_1
X_14038_ _15244_/CLK _14038_/D vssd1 vssd1 vccd1 vccd1 _14038_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06860_ _14730_/Q _14729_/Q vssd1 vssd1 vccd1 vccd1 _12763_/S sky130_fd_sc_hd__nand2_8
XFILLER_94_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06791_ _14589_/Q _06791_/B vssd1 vssd1 vccd1 vccd1 _08391_/B sky130_fd_sc_hd__or2_1
XFILLER_94_175 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08530_ _08531_/C _08530_/B vssd1 vssd1 vccd1 vccd1 _08530_/Y sky130_fd_sc_hd__nor2_8
X_08461_ _13761_/Q _12878_/S _08426_/X vssd1 vssd1 vccd1 vccd1 _08461_/X sky130_fd_sc_hd__o21a_1
XFILLER_24_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_183_clk clkbuf_5_21_0_clk/X vssd1 vssd1 vccd1 vccd1 _15259_/CLK sky130_fd_sc_hd__clkbuf_16
X_07412_ _14743_/Q _07411_/X _07480_/S vssd1 vssd1 vccd1 vccd1 _07412_/X sky130_fd_sc_hd__mux2_8
XFILLER_50_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08392_ _08392_/A _08392_/B vssd1 vssd1 vccd1 vccd1 _08421_/B sky130_fd_sc_hd__nand2_1
XFILLER_148_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07343_ _07327_/A _07329_/Y _07337_/X _07362_/A _07360_/C vssd1 vssd1 vccd1 vccd1
+ _07343_/X sky130_fd_sc_hd__a311o_1
XFILLER_137_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07274_ _07274_/A _07274_/B _07274_/C _07273_/X vssd1 vssd1 vccd1 vccd1 _07363_/A
+ sky130_fd_sc_hd__or4b_2
XFILLER_177_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09013_ _08668_/D _09009_/X _09012_/X _09008_/X vssd1 vssd1 vccd1 vccd1 _09014_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_136_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout601 _12379_/A vssd1 vssd1 vccd1 vccd1 _12521_/A sky130_fd_sc_hd__buf_12
XFILLER_144_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout612 _08457_/A vssd1 vssd1 vccd1 vccd1 _12489_/S0 sky130_fd_sc_hd__buf_12
XFILLER_132_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09915_ _11868_/A1 _14276_/Q _09925_/S vssd1 vssd1 vccd1 vccd1 _14276_/D sky130_fd_sc_hd__mux2_1
Xfanout623 _14598_/Q vssd1 vssd1 vccd1 vccd1 _12545_/S sky130_fd_sc_hd__buf_12
XFILLER_99_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout634 _13229_/A vssd1 vssd1 vccd1 vccd1 _13233_/A sky130_fd_sc_hd__buf_6
Xfanout645 _07965_/C1 vssd1 vssd1 vccd1 vccd1 _07987_/C1 sky130_fd_sc_hd__buf_6
X_09846_ _14210_/Q _13080_/B2 _09858_/S vssd1 vssd1 vccd1 vccd1 _14210_/D sky130_fd_sc_hd__mux2_1
XTAP_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09777_ _14144_/Q _13332_/A0 _09790_/S vssd1 vssd1 vccd1 vccd1 _14144_/D sky130_fd_sc_hd__mux2_1
XTAP_3016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06989_ _08392_/A _08390_/C _06988_/A vssd1 vssd1 vccd1 vccd1 _09829_/C sky130_fd_sc_hd__a21o_1
XTAP_3027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08728_ _13512_/Q _08750_/A2 _08747_/A2 _13544_/Q vssd1 vssd1 vccd1 vccd1 _08728_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_3049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08659_ _08722_/A _08659_/B _08659_/C vssd1 vssd1 vccd1 vccd1 _08659_/X sky130_fd_sc_hd__or3_4
XFILLER_26_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_174_clk clkbuf_5_23_0_clk/X vssd1 vssd1 vccd1 vccd1 _15203_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_15_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_234 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11670_ _13345_/A0 _15102_/Q _11670_/S vssd1 vssd1 vccd1 vccd1 _15102_/D sky130_fd_sc_hd__mux2_1
XFILLER_187_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10621_ _15562_/Q _10706_/B vssd1 vssd1 vccd1 vccd1 _10621_/X sky130_fd_sc_hd__and2_1
XFILLER_168_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13340_ _13340_/A0 _15670_/Q _13350_/S vssd1 vssd1 vccd1 vccd1 _15670_/D sky130_fd_sc_hd__mux2_1
XFILLER_10_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10552_ _11356_/B _13159_/B vssd1 vssd1 vccd1 vccd1 _10554_/A sky130_fd_sc_hd__or2_1
XFILLER_155_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13271_ _15355_/Q _15602_/Q _13288_/S vssd1 vssd1 vccd1 vccd1 _15602_/D sky130_fd_sc_hd__mux2_1
XFILLER_5_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10483_ _10483_/A _10483_/B vssd1 vssd1 vccd1 vccd1 _13208_/B sky130_fd_sc_hd__or2_4
XFILLER_10_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15010_ _15577_/CLK _15010_/D vssd1 vssd1 vccd1 vccd1 _15010_/Q sky130_fd_sc_hd__dfxtp_1
X_12222_ _12498_/A _12222_/B vssd1 vssd1 vccd1 vccd1 _12222_/X sky130_fd_sc_hd__and2_1
XFILLER_142_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12153_ _12268_/A _12153_/B vssd1 vssd1 vccd1 vccd1 _12153_/X sky130_fd_sc_hd__and2_1
XFILLER_162_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11104_ _11115_/S _11015_/X _11094_/Y vssd1 vssd1 vccd1 vccd1 _11105_/B sky130_fd_sc_hd__a21o_1
X_12084_ _12268_/A _12084_/B vssd1 vssd1 vccd1 vccd1 _12084_/X sky130_fd_sc_hd__and2_1
XFILLER_111_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11035_ _11033_/Y _11034_/Y _11330_/A vssd1 vssd1 vccd1 vccd1 _11035_/X sky130_fd_sc_hd__mux2_1
XFILLER_94_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12986_ _15475_/Q _10834_/S _13025_/B1 _12985_/X vssd1 vssd1 vccd1 vccd1 _15475_/D
+ sky130_fd_sc_hd__a22o_1
XTAP_3561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14725_ _15552_/CLK _14725_/D vssd1 vssd1 vccd1 vccd1 _14725_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11937_ _15275_/Q _15243_/Q _15211_/Q _15142_/Q _12543_/S _12544_/A vssd1 vssd1 vccd1
+ vccd1 _11938_/B sky130_fd_sc_hd__mux4_1
XFILLER_45_584 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_165_clk clkbuf_5_22_0_clk/X vssd1 vssd1 vccd1 vccd1 _15334_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_60_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14656_ _15628_/CLK _14656_/D vssd1 vssd1 vccd1 vccd1 _14656_/Q sky130_fd_sc_hd__dfxtp_1
X_11868_ _15289_/Q _11868_/A1 _11878_/S vssd1 vssd1 vccd1 vccd1 _15289_/D sky130_fd_sc_hd__mux2_1
XFILLER_60_576 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13607_ _15375_/CLK _13607_/D vssd1 vssd1 vccd1 vccd1 _13607_/Q sky130_fd_sc_hd__dfxtp_1
X_10819_ _14851_/Q _07242_/X _12885_/S vssd1 vssd1 vccd1 vccd1 _14851_/D sky130_fd_sc_hd__mux2_1
XFILLER_20_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11799_ _15222_/Q _13332_/A0 _11816_/S vssd1 vssd1 vccd1 vccd1 _15222_/D sky130_fd_sc_hd__mux2_1
X_14587_ _14649_/CLK _14587_/D vssd1 vssd1 vccd1 vccd1 _14587_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_118_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13538_ _13642_/CLK _13538_/D vssd1 vssd1 vccd1 vccd1 _13538_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_185_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13469_ _14510_/CLK _13469_/D vssd1 vssd1 vccd1 vccd1 _13469_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_174_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15208_ _15208_/CLK _15208_/D vssd1 vssd1 vccd1 vccd1 _15208_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_142_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15139_ _15326_/CLK _15139_/D vssd1 vssd1 vccd1 vccd1 _15139_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_141_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07961_ _13556_/Q _13555_/Q _07961_/C _07961_/D vssd1 vssd1 vccd1 vccd1 _07973_/D
+ sky130_fd_sc_hd__and4_2
XFILLER_99_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09700_ _11680_/A0 _14070_/Q _09723_/S vssd1 vssd1 vccd1 vccd1 _14070_/D sky130_fd_sc_hd__mux2_1
X_06912_ _06719_/Y _13462_/Q _06919_/A _13461_/Q vssd1 vssd1 vccd1 vccd1 _06923_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_110_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07892_ _13538_/Q _13537_/Q vssd1 vssd1 vccd1 vccd1 _07900_/D sky130_fd_sc_hd__and2_1
XFILLER_114_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09631_ _14004_/Q _11853_/A1 _09661_/S vssd1 vssd1 vccd1 vccd1 _14004_/D sky130_fd_sc_hd__mux2_1
X_06843_ _08405_/A _14905_/Q vssd1 vssd1 vccd1 vccd1 _06843_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_55_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09562_ _10032_/A _13318_/D vssd1 vssd1 vccd1 vccd1 _09562_/Y sky130_fd_sc_hd__nor2_8
XFILLER_167_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06774_ _14897_/Q _14898_/Q vssd1 vssd1 vccd1 vccd1 _10561_/C sky130_fd_sc_hd__nor2_2
X_08513_ _08513_/A _08537_/A vssd1 vssd1 vccd1 vccd1 _08513_/Y sky130_fd_sc_hd__nor2_8
X_09493_ _09477_/X _09480_/X _09487_/X _09492_/X vssd1 vssd1 vccd1 vccd1 _09493_/X
+ sky130_fd_sc_hd__o22a_1
Xclkbuf_leaf_156_clk clkbuf_5_19_0_clk/X vssd1 vssd1 vccd1 vccd1 _15489_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_169_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08444_ _13752_/Q _12878_/S _08426_/X _08443_/X vssd1 vssd1 vccd1 vccd1 _13752_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_24_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08375_ _10991_/B _10990_/A vssd1 vssd1 vccd1 vccd1 _08375_/Y sky130_fd_sc_hd__nor2_1
XFILLER_165_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07326_ _13908_/Q _15495_/Q _07334_/S vssd1 vssd1 vccd1 vccd1 _07327_/A sky130_fd_sc_hd__mux2_8
XFILLER_176_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07257_ _15322_/Q _15478_/Q _07340_/S vssd1 vssd1 vccd1 vccd1 _07258_/A sky130_fd_sc_hd__mux2_8
XFILLER_137_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07188_ _15362_/Q _15069_/Q _07188_/S vssd1 vssd1 vccd1 vccd1 _07188_/X sky130_fd_sc_hd__mux2_8
XFILLER_151_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout420 _10731_/B vssd1 vssd1 vccd1 vccd1 _10706_/B sky130_fd_sc_hd__buf_8
XFILLER_48_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout431 _10481_/B vssd1 vssd1 vccd1 vccd1 _10523_/A2 sky130_fd_sc_hd__buf_12
Xfanout442 _07373_/X vssd1 vssd1 vccd1 vccd1 _07500_/S sky130_fd_sc_hd__buf_12
Xfanout453 _10244_/S vssd1 vssd1 vccd1 vccd1 _10630_/S sky130_fd_sc_hd__buf_8
XFILLER_63_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout464 _13123_/A vssd1 vssd1 vccd1 vccd1 _08507_/A sky130_fd_sc_hd__buf_12
XFILLER_86_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout475 _12502_/S vssd1 vssd1 vccd1 vccd1 _12490_/A sky130_fd_sc_hd__buf_12
XFILLER_86_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout486 _07334_/S vssd1 vssd1 vccd1 vccd1 _07339_/S sky130_fd_sc_hd__buf_12
XFILLER_171_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09829_ _13120_/S _09829_/B _09829_/C vssd1 vssd1 vccd1 vccd1 _09829_/X sky130_fd_sc_hd__or3_1
XFILLER_100_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout497 _15043_/Q vssd1 vssd1 vccd1 vccd1 _08145_/S sky130_fd_sc_hd__buf_6
XFILLER_100_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12840_ _14734_/Q _15368_/Q _12871_/S vssd1 vssd1 vccd1 vccd1 _15368_/D sky130_fd_sc_hd__mux2_1
XFILLER_73_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12771_ _15065_/Q _12834_/B vssd1 vssd1 vccd1 vccd1 _12771_/X sky130_fd_sc_hd__or2_1
XTAP_1400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_147_clk clkbuf_5_25_0_clk/X vssd1 vssd1 vccd1 vccd1 _15429_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_27_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14510_ _14510_/CLK _14510_/D vssd1 vssd1 vccd1 vccd1 _14510_/Q sky130_fd_sc_hd__dfxtp_2
X_11722_ _15151_/Q _13330_/A0 _11741_/S vssd1 vssd1 vccd1 vccd1 _15151_/D sky130_fd_sc_hd__mux2_1
XFILLER_14_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15490_ _15526_/CLK _15490_/D vssd1 vssd1 vccd1 vccd1 _15490_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14441_ _14537_/CLK _14441_/D vssd1 vssd1 vccd1 vccd1 _14441_/Q sky130_fd_sc_hd__dfxtp_1
X_11653_ _13328_/A0 _15085_/Q _11670_/S vssd1 vssd1 vccd1 vccd1 _15085_/D sky130_fd_sc_hd__mux2_1
XFILLER_42_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10604_ _10601_/X _10602_/X _10603_/X _10734_/A2 _15048_/Q vssd1 vssd1 vccd1 vccd1
+ _10604_/X sky130_fd_sc_hd__o32a_4
XFILLER_174_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14372_ _14470_/CLK _14372_/D vssd1 vssd1 vccd1 vccd1 _14372_/Q sky130_fd_sc_hd__dfxtp_1
X_11584_ _11584_/A _11584_/B vssd1 vssd1 vccd1 vccd1 _11585_/B sky130_fd_sc_hd__nor2_1
XFILLER_7_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13323_ _13323_/A0 _15653_/Q _13345_/S vssd1 vssd1 vccd1 vccd1 _15653_/D sky130_fd_sc_hd__mux2_1
X_10535_ _11616_/A _13242_/B _10462_/B vssd1 vssd1 vccd1 vccd1 _10535_/X sky130_fd_sc_hd__a21bo_1
XFILLER_127_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_182_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13254_ _15338_/Q _15585_/Q _13291_/S vssd1 vssd1 vccd1 vccd1 _15585_/D sky130_fd_sc_hd__mux2_1
XFILLER_127_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_92 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10466_ _07208_/A _10523_/A2 _10465_/X vssd1 vssd1 vccd1 vccd1 _13233_/B sky130_fd_sc_hd__a21o_4
XFILLER_50_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12205_ _12481_/A _12205_/B _12205_/C vssd1 vssd1 vccd1 vccd1 _12205_/X sky130_fd_sc_hd__and3_1
XFILLER_108_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13185_ _13183_/Y _13184_/X _15562_/Q _13241_/A2 vssd1 vssd1 vccd1 vccd1 _15562_/D
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_135_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10397_ _07312_/X _10457_/A2 _10396_/X vssd1 vssd1 vccd1 vccd1 _11414_/C sky130_fd_sc_hd__a21oi_4
XFILLER_97_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12136_ _12481_/A _12136_/B _12136_/C vssd1 vssd1 vccd1 vccd1 _12136_/X sky130_fd_sc_hd__and3_1
XFILLER_145_91 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12067_ _12596_/A _12067_/B _12067_/C vssd1 vssd1 vccd1 vccd1 _12067_/X sky130_fd_sc_hd__and3_1
XFILLER_1_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11018_ _11037_/A _11521_/A vssd1 vssd1 vccd1 vccd1 _11020_/A sky130_fd_sc_hd__and2_1
XFILLER_92_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_138_clk clkbuf_5_29_0_clk/X vssd1 vssd1 vccd1 vccd1 _15199_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_3391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12969_ _10619_/X _14870_/Q _13029_/S vssd1 vssd1 vccd1 vccd1 _12969_/X sky130_fd_sc_hd__mux2_4
XFILLER_73_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14708_ _15646_/CLK _14708_/D vssd1 vssd1 vccd1 vccd1 _14708_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14639_ _15645_/CLK _14639_/D vssd1 vssd1 vccd1 vccd1 _14639_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_159_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08160_ _13667_/Q _10285_/S _08155_/X _08159_/X vssd1 vssd1 vccd1 vccd1 _13667_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_158_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07111_ _14833_/Q _07115_/B _07163_/A vssd1 vssd1 vccd1 vccd1 _07111_/X sky130_fd_sc_hd__and3_4
X_08091_ _14765_/Q _08083_/A _08090_/Y vssd1 vssd1 vccd1 vccd1 _13648_/D sky130_fd_sc_hd__o21a_1
XFILLER_9_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07042_ _14626_/Q _14658_/Q _07078_/S vssd1 vssd1 vccd1 vccd1 _07042_/X sky130_fd_sc_hd__mux2_1
XFILLER_106_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08993_ _14361_/Q _15177_/Q _13816_/Q _14555_/Q _09005_/S _09523_/A1 vssd1 vssd1
+ vccd1 vccd1 _08994_/B sky130_fd_sc_hd__mux4_1
XFILLER_87_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07944_ _07964_/A _07943_/X input35/X vssd1 vssd1 vccd1 vccd1 _07944_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_130_879 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07875_ _14758_/Q _07874_/A _07874_/Y _08002_/C1 vssd1 vssd1 vccd1 vccd1 _13533_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_18_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09614_ _13988_/Q _11761_/A0 _09628_/S vssd1 vssd1 vccd1 vccd1 _13988_/D sky130_fd_sc_hd__mux2_1
X_06826_ _08078_/B _08085_/S vssd1 vssd1 vccd1 vccd1 _12647_/B sky130_fd_sc_hd__nand2b_4
XFILLER_84_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09545_ _14485_/Q _14453_/Q _13874_/Q _14227_/Q _09469_/S _09546_/S1 vssd1 vssd1
+ vccd1 vccd1 _09545_/X sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_129_clk clkbuf_5_31_0_clk/X vssd1 vssd1 vccd1 vccd1 _14510_/CLK sky130_fd_sc_hd__clkbuf_16
X_06757_ _13445_/Q vssd1 vssd1 vccd1 vccd1 _06757_/Y sky130_fd_sc_hd__inv_2
XFILLER_110_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09476_ _09543_/A _09476_/B vssd1 vssd1 vccd1 vccd1 _09476_/X sky130_fd_sc_hd__or2_1
XFILLER_70_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06688_ _13476_/Q vssd1 vssd1 vccd1 vccd1 _06688_/Y sky130_fd_sc_hd__inv_2
X_08427_ _14613_/Q _08390_/C _08425_/X _10764_/S vssd1 vssd1 vccd1 vccd1 _08427_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_180_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08358_ _08318_/X _08357_/Y _11297_/S vssd1 vssd1 vccd1 vccd1 _08358_/X sky130_fd_sc_hd__mux2_1
XFILLER_50_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07309_ _07351_/A _07350_/C _07350_/B vssd1 vssd1 vccd1 vccd1 _07309_/X sky130_fd_sc_hd__o21a_1
X_08289_ _08273_/X _08288_/X _11088_/S vssd1 vssd1 vccd1 vccd1 _08289_/X sky130_fd_sc_hd__mux2_1
XFILLER_164_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10320_ _14705_/Q _14890_/Q _10735_/S vssd1 vssd1 vccd1 vccd1 _14705_/D sky130_fd_sc_hd__mux2_1
XFILLER_125_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10251_ _14636_/Q _14789_/Q _10695_/S vssd1 vssd1 vccd1 vccd1 _14636_/D sky130_fd_sc_hd__mux2_1
XFILLER_106_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10182_ _11868_/A1 _14566_/Q _10192_/S vssd1 vssd1 vccd1 vccd1 _14566_/D sky130_fd_sc_hd__mux2_1
XFILLER_59_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout250 _08521_/Y vssd1 vssd1 vccd1 vccd1 _08683_/A2 sky130_fd_sc_hd__clkbuf_16
X_14990_ _15021_/CLK _14990_/D vssd1 vssd1 vccd1 vccd1 _14990_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout261 _07193_/S vssd1 vssd1 vccd1 vccd1 _07188_/S sky130_fd_sc_hd__buf_12
Xfanout272 _08510_/X vssd1 vssd1 vccd1 vccd1 _08690_/B1 sky130_fd_sc_hd__buf_6
X_13941_ _14537_/CLK _13941_/D vssd1 vssd1 vccd1 vccd1 _13941_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout283 _07500_/X vssd1 vssd1 vccd1 vccd1 _11883_/A1 sky130_fd_sc_hd__buf_6
Xfanout294 _07480_/X vssd1 vssd1 vccd1 vccd1 _13104_/B2 sky130_fd_sc_hd__buf_8
XFILLER_74_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13872_ _15526_/CLK _13872_/D vssd1 vssd1 vccd1 vccd1 _13872_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15611_ _15623_/CLK _15611_/D vssd1 vssd1 vccd1 vccd1 _15611_/Q sky130_fd_sc_hd__dfxtp_1
X_12823_ _13442_/Q _12647_/B _08030_/Y _13609_/Q _12743_/A vssd1 vssd1 vccd1 vccd1
+ _12823_/X sky130_fd_sc_hd__a221o_1
XFILLER_15_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15542_ _15542_/CLK _15542_/D vssd1 vssd1 vccd1 vccd1 _15542_/Q sky130_fd_sc_hd__dfxtp_1
X_12754_ _15356_/Q _12754_/B vssd1 vssd1 vccd1 vccd1 _12755_/B sky130_fd_sc_hd__or2_1
XTAP_1241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11705_ _11847_/A1 _15136_/Q _11708_/S vssd1 vssd1 vccd1 vccd1 _15136_/D sky130_fd_sc_hd__mux2_1
XTAP_1274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12685_ _12737_/A _12685_/B vssd1 vssd1 vccd1 vccd1 _12685_/X sky130_fd_sc_hd__or2_1
XTAP_1285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15473_ _15508_/CLK _15473_/D vssd1 vssd1 vccd1 vccd1 _15473_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14424_ _15668_/CLK _14424_/D vssd1 vssd1 vccd1 vccd1 _14424_/Q sky130_fd_sc_hd__dfxtp_1
X_11636_ _11635_/X _15073_/Q _11641_/S vssd1 vssd1 vccd1 vccd1 _15073_/D sky130_fd_sc_hd__mux2_1
XFILLER_187_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_175_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11567_ _11576_/C _11567_/B vssd1 vssd1 vccd1 vccd1 _11567_/X sky130_fd_sc_hd__xor2_1
XFILLER_11_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14355_ _15203_/CLK _14355_/D vssd1 vssd1 vccd1 vccd1 _14355_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_183_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10518_ _11536_/C _11521_/A vssd1 vssd1 vccd1 vccd1 _10519_/B sky130_fd_sc_hd__and2_1
X_13306_ _15638_/Q _12770_/B _13316_/S vssd1 vssd1 vccd1 vccd1 _15638_/D sky130_fd_sc_hd__mux2_1
XFILLER_183_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14286_ _15332_/CLK _14286_/D vssd1 vssd1 vccd1 vccd1 _14286_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11498_ _11536_/B _11498_/B vssd1 vssd1 vccd1 vccd1 _11500_/B sky130_fd_sc_hd__xnor2_1
XFILLER_109_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13237_ _13236_/A _13236_/B _13214_/B _11600_/A vssd1 vssd1 vccd1 vccd1 _13237_/X
+ sky130_fd_sc_hd__a211o_1
X_10449_ _10520_/A1 _13782_/Q _13750_/Q _10520_/B2 vssd1 vssd1 vccd1 vccd1 _10449_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_97_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13168_ _13251_/A _13168_/B vssd1 vssd1 vccd1 vccd1 _13168_/Y sky130_fd_sc_hd__nand2_1
XFILLER_97_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12119_ _12115_/X _12116_/X _12490_/A vssd1 vssd1 vccd1 vccd1 _12119_/X sky130_fd_sc_hd__mux2_1
XFILLER_111_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13099_ _15517_/Q _13139_/S _13042_/A _13098_/X vssd1 vssd1 vccd1 vccd1 _15517_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_27_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07660_ _10099_/B _07660_/B vssd1 vssd1 vccd1 vccd1 _07736_/A sky130_fd_sc_hd__nand2_8
XFILLER_93_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_882 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07591_ _13459_/Q _07603_/C vssd1 vssd1 vccd1 vccd1 _07592_/B sky130_fd_sc_hd__xnor2_1
XFILLER_25_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09330_ _13864_/Q _14217_/Q _09469_/S vssd1 vssd1 vccd1 vccd1 _09330_/X sky130_fd_sc_hd__mux2_1
XFILLER_80_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_362 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09261_ _09543_/A _09261_/B vssd1 vssd1 vccd1 vccd1 _09261_/X sky130_fd_sc_hd__or2_1
XFILLER_60_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08212_ _13703_/Q _11874_/A1 _08216_/S vssd1 vssd1 vccd1 vccd1 _13703_/D sky130_fd_sc_hd__mux2_1
X_09192_ _09427_/A1 _09190_/X _09191_/X vssd1 vssd1 vccd1 vccd1 _09192_/X sky130_fd_sc_hd__a21o_1
XFILLER_159_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08143_ _08093_/B _08141_/X _08142_/Y _08121_/X vssd1 vssd1 vccd1 vccd1 _08143_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_174_551 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08074_ _08074_/A _08074_/B vssd1 vssd1 vccd1 vccd1 _08083_/A sky130_fd_sc_hd__nand2_4
XFILLER_119_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07025_ _07024_/X _13587_/Q _12662_/S vssd1 vssd1 vccd1 vccd1 _07025_/X sky130_fd_sc_hd__mux2_1
XFILLER_162_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08976_ _14232_/Q _14264_/Q _14296_/Q _14328_/Q _09225_/S0 _09225_/S1 vssd1 vssd1
+ vccd1 vccd1 _08976_/X sky130_fd_sc_hd__mux4_1
XFILLER_76_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07927_ _14739_/Q _08012_/A2 _07926_/Y _08084_/C1 vssd1 vssd1 vccd1 vccd1 _13546_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_130_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07858_ _13529_/Q _13528_/Q _13527_/Q _07858_/D vssd1 vssd1 vccd1 vccd1 _07869_/D
+ sky130_fd_sc_hd__and4_2
XFILLER_57_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06809_ _08465_/B _06808_/X _15615_/Q vssd1 vssd1 vccd1 vccd1 _06809_/X sky130_fd_sc_hd__o21a_1
XFILLER_28_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_424 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07789_ _07816_/A _07789_/B vssd1 vssd1 vccd1 vccd1 _07789_/Y sky130_fd_sc_hd__nand2_1
XFILLER_45_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09528_ _15106_/Q _08540_/B _09527_/X _08501_/A vssd1 vssd1 vccd1 vccd1 _09528_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_169_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09459_ _09546_/S1 _09457_/X _09458_/X vssd1 vssd1 vccd1 vccd1 _09459_/X sky130_fd_sc_hd__a21o_1
XPHY_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12470_ _13964_/Q _13706_/Q _12470_/S vssd1 vssd1 vccd1 vccd1 _12471_/B sky130_fd_sc_hd__mux2_1
XFILLER_131_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11421_ _11421_/A _11421_/B vssd1 vssd1 vccd1 vccd1 _11421_/X sky130_fd_sc_hd__or2_1
XFILLER_138_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14140_ _15658_/CLK _14140_/D vssd1 vssd1 vccd1 vccd1 _14140_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_165_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11352_ _15042_/Q _08232_/A _11347_/Y _11351_/X vssd1 vssd1 vccd1 vccd1 _11352_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_125_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10303_ _14688_/Q _14873_/Q _10615_/S vssd1 vssd1 vccd1 vccd1 _14688_/D sky130_fd_sc_hd__mux2_1
X_14071_ _15253_/CLK _14071_/D vssd1 vssd1 vccd1 vccd1 _14071_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_106_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11283_ _11283_/A _11283_/B vssd1 vssd1 vccd1 vccd1 _11283_/X sky130_fd_sc_hd__or2_1
XFILLER_180_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13022_ _15487_/Q _13119_/S _13025_/B1 _13021_/X vssd1 vssd1 vccd1 vccd1 _15487_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_79_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10234_ _14619_/Q _14772_/Q _10610_/S vssd1 vssd1 vccd1 vccd1 _14619_/D sky130_fd_sc_hd__mux2_1
XFILLER_3_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10165_ _14714_/Q _14716_/Q _11710_/A _11743_/C vssd1 vssd1 vccd1 vccd1 _10165_/X
+ sky130_fd_sc_hd__or4_4
XFILLER_126_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14973_ _15021_/CLK _14973_/D vssd1 vssd1 vccd1 vccd1 _14973_/Q sky130_fd_sc_hd__dfxtp_1
X_10096_ _14452_/Q _13349_/A0 _10097_/S vssd1 vssd1 vccd1 vccd1 _14452_/D sky130_fd_sc_hd__mux2_1
XFILLER_59_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13924_ _15666_/CLK _13924_/D vssd1 vssd1 vccd1 vccd1 _13924_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_142_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13855_ _14530_/CLK _13855_/D vssd1 vssd1 vccd1 vccd1 _13855_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_74_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12806_ _15070_/Q _12834_/B vssd1 vssd1 vccd1 vccd1 _12806_/X sky130_fd_sc_hd__or2_1
XFILLER_90_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13786_ _15393_/CLK _13786_/D vssd1 vssd1 vccd1 vccd1 _13786_/Q sky130_fd_sc_hd__dfxtp_4
X_10998_ _11356_/C _11399_/A _08316_/B vssd1 vssd1 vccd1 vccd1 _10998_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_90_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15525_ _15525_/CLK _15525_/D vssd1 vssd1 vccd1 vccd1 _15525_/Q sky130_fd_sc_hd__dfxtp_1
X_12737_ _12737_/A _12737_/B vssd1 vssd1 vccd1 vccd1 _12737_/X sky130_fd_sc_hd__or2_1
XTAP_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15456_ _15643_/CLK _15456_/D vssd1 vssd1 vccd1 vccd1 _15456_/Q sky130_fd_sc_hd__dfxtp_1
X_12668_ _15051_/Q _12667_/Y _12792_/B vssd1 vssd1 vccd1 vccd1 _12668_/X sky130_fd_sc_hd__mux2_1
XFILLER_175_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14407_ _15668_/CLK _14407_/D vssd1 vssd1 vccd1 vccd1 _14407_/Q sky130_fd_sc_hd__dfxtp_1
X_11619_ _11611_/A _11611_/B _11612_/B wire360/X vssd1 vssd1 vccd1 vccd1 _11619_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_15387_ _15389_/CLK _15387_/D vssd1 vssd1 vccd1 vccd1 _15387_/Q sky130_fd_sc_hd__dfxtp_1
X_12599_ _14485_/Q _14453_/Q _13874_/Q _14227_/Q _12522_/S _12521_/A vssd1 vssd1 vccd1
+ vccd1 _12599_/X sky130_fd_sc_hd__mux4_1
XFILLER_128_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14338_ _14468_/CLK _14338_/D vssd1 vssd1 vccd1 vccd1 _14338_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_768 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14269_ _15181_/CLK _14269_/D vssd1 vssd1 vccd1 vccd1 _14269_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_171_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_598 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_632 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08830_ _13853_/Q _13072_/B2 _08846_/S vssd1 vssd1 vccd1 vccd1 _13853_/D sky130_fd_sc_hd__mux2_1
XFILLER_111_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08761_ _14612_/Q _14611_/Q _08772_/A vssd1 vssd1 vccd1 vccd1 _08778_/D sky130_fd_sc_hd__or3_4
XFILLER_97_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07712_ _13491_/Q _07712_/B vssd1 vssd1 vccd1 vccd1 _07713_/B sky130_fd_sc_hd__xnor2_1
X_08692_ _13453_/Q _08746_/A2 _08750_/A2 _13517_/Q _08691_/X vssd1 vssd1 vccd1 vccd1
+ _08692_/X sky130_fd_sc_hd__a221o_1
XFILLER_38_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07643_ _13473_/Q _07647_/C vssd1 vssd1 vccd1 vccd1 _07644_/B sky130_fd_sc_hd__xnor2_1
XFILLER_80_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07574_ _14743_/Q _07629_/A _07573_/Y _12788_/C1 vssd1 vssd1 vccd1 vccd1 _13454_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_80_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09313_ _08519_/A _09311_/X _09312_/X vssd1 vssd1 vccd1 vccd1 _09317_/B sky130_fd_sc_hd__a21o_1
XFILLER_90_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_654 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_60_clk _15031_/CLK vssd1 vssd1 vccd1 vccd1 _15020_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_142_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_1048 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09244_ _14471_/Q _14439_/Q _13860_/Q _14213_/Q _09557_/S _09550_/A1 vssd1 vssd1
+ vccd1 vccd1 _09244_/X sky130_fd_sc_hd__mux4_1
XFILLER_178_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09175_ _09446_/A1 _09419_/A2 _09174_/X _09450_/B1 vssd1 vssd1 vccd1 vccd1 _09175_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_108_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08126_ _08133_/S _06760_/Y _08093_/B vssd1 vssd1 vccd1 vccd1 _08126_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_147_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08057_ _14750_/Q _13628_/Q _08066_/S vssd1 vssd1 vccd1 vccd1 _13628_/D sky130_fd_sc_hd__mux2_1
XFILLER_122_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07008_ _07007_/X _14735_/Q _07098_/S vssd1 vssd1 vccd1 vccd1 _13581_/D sky130_fd_sc_hd__mux2_1
Xoutput37 _07173_/X vssd1 vssd1 vccd1 vccd1 ext_address[11] sky130_fd_sc_hd__clkbuf_2
XFILLER_122_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_203 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput48 _07184_/X vssd1 vssd1 vccd1 vccd1 ext_address[22] sky130_fd_sc_hd__clkbuf_2
Xoutput59 _07165_/X vssd1 vssd1 vccd1 vccd1 ext_address[3] sky130_fd_sc_hd__clkbuf_2
XFILLER_1_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08959_ _09421_/A1 _08955_/X _08958_/X _08954_/X vssd1 vssd1 vccd1 vccd1 _08959_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_56_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11970_ _14070_/Q _14038_/Q _12079_/S vssd1 vssd1 vccd1 vccd1 _11970_/X sky130_fd_sc_hd__mux2_1
XTAP_3935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10921_ _14943_/Q _10929_/B _10920_/Y _11475_/A vssd1 vssd1 vccd1 vccd1 _14943_/D
+ sky130_fd_sc_hd__o22a_1
XTAP_3968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_1095 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10852_ _14884_/Q _13784_/Q _12929_/S vssd1 vssd1 vccd1 vccd1 _14884_/D sky130_fd_sc_hd__mux2_1
X_13640_ _15398_/CLK _13640_/D vssd1 vssd1 vccd1 vccd1 _13640_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10783_ _14815_/Q hold2/X _12928_/S vssd1 vssd1 vccd1 vccd1 _14815_/D sky130_fd_sc_hd__mux2_1
XPHY_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13571_ _13642_/CLK _13571_/D vssd1 vssd1 vccd1 vccd1 _13571_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_158_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_51_clk clkbuf_5_8_0_clk/X vssd1 vssd1 vccd1 vccd1 _14966_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_9_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15310_ _15507_/CLK _15310_/D vssd1 vssd1 vccd1 vccd1 _15310_/Q sky130_fd_sc_hd__dfxtp_1
X_12522_ _14094_/Q _14062_/Q _12522_/S vssd1 vssd1 vccd1 vccd1 _12522_/X sky130_fd_sc_hd__mux2_1
XPHY_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_859 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15241_ _15273_/CLK _15241_/D vssd1 vssd1 vccd1 vccd1 _15241_/Q sky130_fd_sc_hd__dfxtp_1
X_12453_ _14091_/Q _14059_/Q _12453_/S vssd1 vssd1 vccd1 vccd1 _12453_/X sky130_fd_sc_hd__mux2_1
XFILLER_138_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11404_ _11404_/A _11404_/B vssd1 vssd1 vccd1 vccd1 _11404_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_184_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15172_ _15172_/CLK _15172_/D vssd1 vssd1 vccd1 vccd1 _15172_/Q sky130_fd_sc_hd__dfxtp_1
X_12384_ _14088_/Q _14056_/Q _12614_/S vssd1 vssd1 vccd1 vccd1 _12384_/X sky130_fd_sc_hd__mux2_1
XFILLER_181_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11335_ _15039_/Q _11346_/A2 _11334_/X vssd1 vssd1 vccd1 vccd1 _15039_/D sky130_fd_sc_hd__a21o_1
X_14123_ _15518_/CLK _14123_/D vssd1 vssd1 vccd1 vccd1 _14123_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_768 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_351 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14054_ _14537_/CLK _14054_/D vssd1 vssd1 vccd1 vccd1 _14054_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11266_ _11249_/Y _11265_/X _11318_/S vssd1 vssd1 vccd1 vccd1 _11266_/X sky130_fd_sc_hd__mux2_1
XFILLER_140_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13005_ _10679_/X _14882_/Q _14903_/Q vssd1 vssd1 vccd1 vccd1 _13005_/X sky130_fd_sc_hd__mux2_4
X_10217_ input11/X _12515_/C1 _13282_/S vssd1 vssd1 vccd1 vccd1 _14602_/D sky130_fd_sc_hd__mux2_1
X_11197_ _11199_/A _11197_/B vssd1 vssd1 vccd1 vccd1 _11197_/Y sky130_fd_sc_hd__nor2_1
XFILLER_67_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10148_ _14533_/Q _13082_/B2 _10159_/S vssd1 vssd1 vccd1 vccd1 _14533_/D sky130_fd_sc_hd__mux2_1
X_14956_ _15021_/CLK _14956_/D vssd1 vssd1 vccd1 vccd1 _14956_/Q sky130_fd_sc_hd__dfxtp_1
X_10079_ _14435_/Q _13078_/B2 _10092_/S vssd1 vssd1 vccd1 vccd1 _14435_/D sky130_fd_sc_hd__mux2_1
XFILLER_36_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13907_ _15664_/CLK _13907_/D vssd1 vssd1 vccd1 vccd1 _13907_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_130_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14887_ _15607_/CLK _14887_/D vssd1 vssd1 vccd1 vccd1 _14887_/Q sky130_fd_sc_hd__dfxtp_1
X_13838_ _15544_/CLK _13838_/D vssd1 vssd1 vccd1 vccd1 _13838_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13769_ _14863_/CLK _13769_/D vssd1 vssd1 vccd1 vccd1 _13769_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_94_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_42_clk clkbuf_5_9_0_clk/X vssd1 vssd1 vccd1 vccd1 _15581_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_148_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15508_ _15508_/CLK _15508_/D vssd1 vssd1 vccd1 vccd1 _15508_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07290_ _07339_/S _13919_/Q _07288_/Y vssd1 vssd1 vccd1 vccd1 _07292_/A sky130_fd_sc_hd__o21ai_4
XFILLER_31_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15439_ _15632_/CLK _15439_/D vssd1 vssd1 vccd1 vccd1 _15439_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_307 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_172_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09931_ _13318_/D _09964_/B vssd1 vssd1 vccd1 vccd1 _09931_/Y sky130_fd_sc_hd__nand2b_4
X_09862_ _14226_/Q _11816_/A1 _09863_/S vssd1 vssd1 vccd1 vccd1 _14226_/D sky130_fd_sc_hd__mux2_1
XTAP_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08813_ _11847_/A1 _13839_/Q _08816_/S vssd1 vssd1 vccd1 vccd1 _13839_/D sky130_fd_sc_hd__mux2_1
XFILLER_133_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09793_ _14160_/Q _13348_/A0 _09795_/S vssd1 vssd1 vccd1 vccd1 _14160_/D sky130_fd_sc_hd__mux2_1
XFILLER_100_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08744_ _13478_/Q _08747_/B1 _08741_/X _08742_/X _08743_/X vssd1 vssd1 vccd1 vccd1
+ _08744_/X sky130_fd_sc_hd__a2111o_4
XFILLER_27_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08675_ _13795_/Q _08573_/S _08670_/X _08674_/X vssd1 vssd1 vccd1 vccd1 _13795_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_26_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07626_ _07624_/Y _07655_/A _07629_/A vssd1 vssd1 vccd1 vccd1 _07626_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_26_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07557_ _07560_/B _07556_/Y _07651_/A vssd1 vssd1 vccd1 vccd1 _07557_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_41_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_33_clk clkbuf_5_13_0_clk/X vssd1 vssd1 vccd1 vccd1 _14612_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_167_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07488_ _14762_/Q _07487_/X _07500_/S vssd1 vssd1 vccd1 vccd1 _07488_/X sky130_fd_sc_hd__mux2_8
XFILLER_139_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09227_ _14019_/Q _13987_/Q _09230_/S vssd1 vssd1 vccd1 vccd1 _09227_/X sky130_fd_sc_hd__mux2_1
XFILLER_107_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09158_ _13919_/Q _13081_/A2 _09157_/X vssd1 vssd1 vccd1 vccd1 _13919_/D sky130_fd_sc_hd__a21o_1
XFILLER_181_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08109_ _13653_/Q _10344_/S _08096_/X _08108_/X vssd1 vssd1 vccd1 vccd1 _13653_/D
+ sky130_fd_sc_hd__a22o_1
X_09089_ _13948_/Q _13690_/Q _09407_/S vssd1 vssd1 vccd1 vccd1 _09089_/X sky130_fd_sc_hd__mux2_1
XFILLER_107_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11120_ _11047_/B _11088_/S _11356_/C _13251_/A vssd1 vssd1 vccd1 vccd1 _11371_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_122_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11051_ _11380_/A _11032_/X _11050_/Y _10984_/Y vssd1 vssd1 vccd1 vccd1 _11051_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_77_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10002_ _13323_/A0 _14360_/Q _10028_/S vssd1 vssd1 vccd1 vccd1 _14360_/D sky130_fd_sc_hd__mux2_1
XFILLER_77_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14810_ _15628_/CLK _14810_/D vssd1 vssd1 vccd1 vccd1 _14810_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14741_ _15589_/CLK _14741_/D vssd1 vssd1 vccd1 vccd1 _14741_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_3754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11953_ _15308_/Q _10877_/S _11952_/X vssd1 vssd1 vccd1 vccd1 _15308_/D sky130_fd_sc_hd__a21o_1
XTAP_3765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10904_ _11414_/D _10951_/B vssd1 vssd1 vccd1 vccd1 _10904_/Y sky130_fd_sc_hd__nand2_1
XTAP_3798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14672_ _15452_/CLK _14672_/D vssd1 vssd1 vccd1 vccd1 _14672_/Q sky130_fd_sc_hd__dfxtp_1
X_11884_ _15305_/Q _10344_/S _10564_/A _15208_/Q vssd1 vssd1 vccd1 vccd1 _15305_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_33_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_2_3_0_clk clkbuf_2_3_0_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_2_3_1_clk/A sky130_fd_sc_hd__clkbuf_8
X_13623_ _15375_/CLK _13623_/D vssd1 vssd1 vccd1 vccd1 _13623_/Q sky130_fd_sc_hd__dfxtp_1
X_10835_ _14867_/Q _13801_/Q _12932_/S vssd1 vssd1 vccd1 vccd1 _14867_/D sky130_fd_sc_hd__mux2_1
XFILLER_16_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_24_clk clkbuf_5_3_0_clk/X vssd1 vssd1 vccd1 vccd1 _14405_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_186_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13554_ _13627_/CLK _13554_/D vssd1 vssd1 vccd1 vccd1 _13554_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_73_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10766_ _15430_/Q _14798_/Q _13120_/S vssd1 vssd1 vccd1 vccd1 _14798_/D sky130_fd_sc_hd__mux2_1
XFILLER_160_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12505_ _15332_/Q _13105_/A2 _12504_/X vssd1 vssd1 vccd1 vccd1 _15332_/D sky130_fd_sc_hd__a21o_1
XFILLER_157_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10697_ _15018_/Q _10717_/A2 _10652_/B _15035_/Q _10717_/C1 vssd1 vssd1 vccd1 vccd1
+ _10697_/X sky130_fd_sc_hd__a221o_1
X_13485_ _15393_/CLK _13485_/D vssd1 vssd1 vccd1 vccd1 _13485_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_186_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15224_ _15332_/CLK _15224_/D vssd1 vssd1 vccd1 vccd1 _15224_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_157_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12436_ _15329_/Q _10877_/S _12435_/X vssd1 vssd1 vccd1 vccd1 _15329_/D sky130_fd_sc_hd__a21o_1
XFILLER_172_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15155_ _15332_/CLK _15155_/D vssd1 vssd1 vccd1 vccd1 _15155_/Q sky130_fd_sc_hd__dfxtp_1
X_12367_ _15326_/Q _13149_/S _12366_/X vssd1 vssd1 vccd1 vccd1 _15326_/D sky130_fd_sc_hd__a21o_1
X_14106_ _14525_/CLK _14106_/D vssd1 vssd1 vccd1 vccd1 _14106_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_884 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11318_ _11304_/Y _11330_/B _11318_/S vssd1 vssd1 vccd1 vccd1 _11318_/X sky130_fd_sc_hd__mux2_1
X_12298_ _15323_/Q _13093_/A2 _12297_/X vssd1 vssd1 vccd1 vccd1 _15323_/D sky130_fd_sc_hd__a21o_1
X_15086_ _15133_/CLK _15086_/D vssd1 vssd1 vccd1 vccd1 _15086_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_383 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14037_ _15211_/CLK _14037_/D vssd1 vssd1 vccd1 vccd1 _14037_/Q sky130_fd_sc_hd__dfxtp_1
X_11249_ _11249_/A _11249_/B vssd1 vssd1 vccd1 vccd1 _11249_/Y sky130_fd_sc_hd__nor2_1
XFILLER_141_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_1047 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06790_ _14589_/Q _06791_/B vssd1 vssd1 vccd1 vccd1 _08392_/B sky130_fd_sc_hd__nor2_1
XFILLER_94_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14939_ _15580_/CLK _14939_/D vssd1 vssd1 vccd1 vccd1 _14939_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_1071 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08460_ _13760_/Q _12878_/S _08426_/X _08459_/X vssd1 vssd1 vccd1 vccd1 _13760_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_35_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07411_ _13658_/Q _07483_/A2 _07483_/B1 _14686_/Q _07410_/X vssd1 vssd1 vccd1 vccd1
+ _07411_/X sky130_fd_sc_hd__a221o_1
XFILLER_17_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08391_ _14588_/Q _08391_/B vssd1 vssd1 vccd1 vccd1 _08765_/D sky130_fd_sc_hd__nor2_1
XFILLER_23_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_15_clk clkbuf_5_2_0_clk/X vssd1 vssd1 vccd1 vccd1 _15287_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_52_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07342_ _07337_/A _07337_/B _07339_/X _07341_/Y vssd1 vssd1 vccd1 vccd1 _07360_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_176_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07273_ _07235_/X _07273_/B _07273_/C _07273_/D vssd1 vssd1 vccd1 vccd1 _07273_/X
+ sky130_fd_sc_hd__and4b_1
X_09012_ _15081_/Q _08540_/B _09011_/X _08501_/A vssd1 vssd1 vccd1 vccd1 _09012_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_148_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout602 _14599_/Q vssd1 vssd1 vccd1 vccd1 _12379_/A sky130_fd_sc_hd__clkbuf_16
X_09914_ _13334_/A0 _14275_/Q _09925_/S vssd1 vssd1 vccd1 vccd1 _14275_/D sky130_fd_sc_hd__mux2_1
XFILLER_144_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout613 _08457_/A vssd1 vssd1 vccd1 vccd1 _12499_/S sky130_fd_sc_hd__buf_12
Xfanout624 _08405_/A vssd1 vssd1 vccd1 vccd1 _12522_/S sky130_fd_sc_hd__buf_12
XFILLER_113_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout635 _13739_/Q vssd1 vssd1 vccd1 vccd1 _13229_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_98_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout646 fanout647/X vssd1 vssd1 vccd1 vccd1 _07965_/C1 sky130_fd_sc_hd__buf_8
XTAP_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09845_ _14209_/Q _13078_/B2 _09858_/S vssd1 vssd1 vccd1 vccd1 _14209_/D sky130_fd_sc_hd__mux2_1
XTAP_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_666 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09776_ _14143_/Q _11689_/A0 _09790_/S vssd1 vssd1 vccd1 vccd1 _14143_/D sky130_fd_sc_hd__mux2_1
XFILLER_85_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06988_ _06988_/A _08390_/C vssd1 vssd1 vccd1 vccd1 _08773_/B sky130_fd_sc_hd__or2_4
XTAP_3017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_487 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08727_ _14489_/Q _08537_/Y _08667_/X _13576_/Q _08724_/X vssd1 vssd1 vccd1 vccd1
+ _08727_/X sky130_fd_sc_hd__a221o_1
XTAP_2316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08658_ _15381_/Q _08690_/A2 _08656_/X _08657_/X vssd1 vssd1 vccd1 vccd1 _08659_/C
+ sky130_fd_sc_hd__a211o_1
XTAP_1615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1024 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07609_ _13463_/Q _07610_/C _13464_/Q vssd1 vssd1 vccd1 vccd1 _07609_/Y sky130_fd_sc_hd__a21oi_1
XTAP_1648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08589_ _15391_/Q _08690_/A2 _08690_/B1 _13436_/Q vssd1 vssd1 vccd1 vccd1 _08589_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_53_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_246 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10620_ _14742_/Q _10619_/X _10710_/S vssd1 vssd1 vccd1 vccd1 _14742_/D sky130_fd_sc_hd__mux2_1
XFILLER_179_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10551_ _10551_/A _10551_/B vssd1 vssd1 vccd1 vccd1 _10555_/C sky130_fd_sc_hd__nand2_1
XFILLER_155_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13270_ _15354_/Q _15601_/Q _13309_/A vssd1 vssd1 vccd1 vccd1 _15601_/D sky130_fd_sc_hd__mux2_1
X_10482_ _10507_/A1 _13757_/Q _15415_/Q _10515_/B2 vssd1 vssd1 vccd1 vccd1 _10483_/B
+ sky130_fd_sc_hd__a22o_2
XFILLER_108_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12221_ _14017_/Q _13985_/Q _12476_/S vssd1 vssd1 vccd1 vccd1 _12222_/B sky130_fd_sc_hd__mux2_1
XFILLER_163_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12152_ _14014_/Q _13982_/Q _12269_/S vssd1 vssd1 vccd1 vccd1 _12153_/B sky130_fd_sc_hd__mux2_1
XFILLER_155_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11103_ _11010_/Y _11029_/Y _11115_/S vssd1 vssd1 vccd1 vccd1 _11156_/B sky130_fd_sc_hd__mux2_1
XFILLER_2_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12083_ _14011_/Q _13979_/Q _12269_/S vssd1 vssd1 vccd1 vccd1 _12084_/B sky130_fd_sc_hd__mux2_1
XFILLER_96_408 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11034_ _11034_/A _11034_/B vssd1 vssd1 vccd1 vccd1 _11034_/Y sky130_fd_sc_hd__nor2_1
XFILLER_150_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_64 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12985_ _13078_/B2 _13024_/A2 _12984_/X _13024_/B2 vssd1 vssd1 vccd1 vccd1 _12985_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_3551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14724_ _15548_/CLK _14724_/D vssd1 vssd1 vccd1 vccd1 _14724_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_3584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11936_ _14358_/Q _15174_/Q _13813_/Q _14552_/Q _12543_/S _12544_/A vssd1 vssd1 vccd1
+ vccd1 _11936_/X sky130_fd_sc_hd__mux4_2
XFILLER_73_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14655_ _15626_/CLK _14655_/D vssd1 vssd1 vccd1 vccd1 _14655_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11867_ _15288_/Q _13334_/A0 _11878_/S vssd1 vssd1 vccd1 vccd1 _15288_/D sky130_fd_sc_hd__mux2_1
XTAP_2894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13606_ _15644_/CLK _13606_/D vssd1 vssd1 vccd1 vccd1 _13606_/Q sky130_fd_sc_hd__dfxtp_1
X_10818_ _14850_/Q _07265_/A _10868_/S vssd1 vssd1 vccd1 vccd1 _14850_/D sky130_fd_sc_hd__mux2_1
XFILLER_159_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14586_ _15537_/CLK _14586_/D vssd1 vssd1 vccd1 vccd1 _14586_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_158_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11798_ _15221_/Q _13331_/A0 _11816_/S vssd1 vssd1 vccd1 vccd1 _15221_/D sky130_fd_sc_hd__mux2_1
XFILLER_158_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13537_ _14513_/CLK _13537_/D vssd1 vssd1 vccd1 vccd1 _13537_/Q sky130_fd_sc_hd__dfxtp_1
X_10749_ _15413_/Q _14781_/Q _10759_/S vssd1 vssd1 vccd1 vccd1 _14781_/D sky130_fd_sc_hd__mux2_1
XFILLER_159_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13468_ _14510_/CLK _13468_/D vssd1 vssd1 vccd1 vccd1 _13468_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15207_ _15618_/CLK _15207_/D vssd1 vssd1 vccd1 vccd1 _15207_/Q sky130_fd_sc_hd__dfxtp_1
X_12419_ _14379_/Q _15195_/Q _13834_/Q _14573_/Q _12430_/S _12563_/A vssd1 vssd1 vccd1
+ vccd1 _12419_/X sky130_fd_sc_hd__mux4_1
XFILLER_173_479 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13399_ _15665_/CLK _13399_/D vssd1 vssd1 vccd1 vccd1 _13399_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15138_ _15678_/CLK _15138_/D vssd1 vssd1 vccd1 vccd1 _15138_/Q sky130_fd_sc_hd__dfxtp_1
X_07960_ _14748_/Q _07964_/A _07959_/Y _07965_/C1 vssd1 vssd1 vccd1 vccd1 _13555_/D
+ sky130_fd_sc_hd__o211a_1
X_15069_ _15572_/CLK _15069_/D vssd1 vssd1 vccd1 vccd1 _15069_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_leaf_4_clk clkbuf_5_0_0_clk/X vssd1 vssd1 vccd1 vccd1 _15663_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_141_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06911_ _06717_/Y _13463_/Q _06719_/Y _13462_/Q vssd1 vssd1 vccd1 vccd1 _06911_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_96_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07891_ _14762_/Q _07903_/A _07890_/Y _08016_/C1 vssd1 vssd1 vccd1 vccd1 _13537_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_68_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09630_ _14003_/Q _13319_/A0 _09660_/S vssd1 vssd1 vccd1 vccd1 _14003_/D sky130_fd_sc_hd__mux2_1
X_06842_ _12379_/A _06845_/B _14907_/Q _12559_/A _06841_/X vssd1 vssd1 vccd1 vccd1
+ _06842_/X sky130_fd_sc_hd__o221a_1
XFILLER_55_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09561_ _13938_/Q _09560_/X _12904_/S vssd1 vssd1 vccd1 vccd1 _13938_/D sky130_fd_sc_hd__mux2_1
XFILLER_67_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06773_ _14923_/Q _10561_/B vssd1 vssd1 vccd1 vccd1 _06775_/B sky130_fd_sc_hd__nand2_1
X_08512_ _08519_/B _08512_/B vssd1 vssd1 vccd1 vccd1 _08537_/A sky130_fd_sc_hd__nand2_8
X_09492_ _08510_/B _09488_/X _09489_/X _09491_/X vssd1 vssd1 vccd1 vccd1 _09492_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_130_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08443_ _09435_/A _08390_/C _08425_/X vssd1 vssd1 vccd1 vccd1 _08443_/X sky130_fd_sc_hd__a21o_1
X_08374_ _11037_/A _13199_/B vssd1 vssd1 vccd1 vccd1 _10990_/A sky130_fd_sc_hd__nor2_1
XFILLER_56_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07325_ _07319_/X _07321_/Y _07322_/X _07324_/Y vssd1 vssd1 vccd1 vccd1 _07360_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_177_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07256_ _13923_/Q _15510_/Q _07339_/S vssd1 vssd1 vccd1 vccd1 _07256_/X sky130_fd_sc_hd__mux2_8
XFILLER_136_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_830 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07187_ _15361_/Q _15068_/Q _07188_/S vssd1 vssd1 vccd1 vccd1 _07187_/X sky130_fd_sc_hd__mux2_2
XFILLER_152_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_663 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout410 _11237_/S vssd1 vssd1 vccd1 vccd1 _11232_/S sky130_fd_sc_hd__buf_12
XFILLER_59_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout421 _10573_/X vssd1 vssd1 vccd1 vccd1 _10731_/B sky130_fd_sc_hd__buf_12
XFILLER_63_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout432 _08244_/Y vssd1 vssd1 vccd1 vccd1 _10481_/B sky130_fd_sc_hd__buf_12
Xfanout443 _07499_/A2 vssd1 vssd1 vccd1 vccd1 _07483_/A2 sky130_fd_sc_hd__clkbuf_16
XFILLER_24_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout454 _10343_/S vssd1 vssd1 vccd1 vccd1 _10735_/S sky130_fd_sc_hd__buf_12
XFILLER_87_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout465 _06675_/Y vssd1 vssd1 vccd1 vccd1 _13123_/A sky130_fd_sc_hd__buf_12
XFILLER_24_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout476 _12548_/S vssd1 vssd1 vccd1 vccd1 _12502_/S sky130_fd_sc_hd__buf_12
XFILLER_63_1086 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09828_ _14194_/Q _11883_/A1 _09828_/S vssd1 vssd1 vccd1 vccd1 _14194_/D sky130_fd_sc_hd__mux2_1
Xfanout487 _15527_/Q vssd1 vssd1 vccd1 vccd1 _07334_/S sky130_fd_sc_hd__buf_12
XFILLER_98_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout498 _13038_/S vssd1 vssd1 vccd1 vccd1 _13029_/S sky130_fd_sc_hd__buf_12
XFILLER_171_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09759_ _14127_/Q _13347_/A0 _09762_/S vssd1 vssd1 vccd1 vccd1 _14127_/D sky130_fd_sc_hd__mux2_1
XFILLER_39_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12770_ _12828_/A _12770_/B vssd1 vssd1 vccd1 vccd1 _12770_/X sky130_fd_sc_hd__or2_1
XTAP_1401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11721_ _15150_/Q _13329_/A0 _11741_/S vssd1 vssd1 vccd1 vccd1 _15150_/D sky130_fd_sc_hd__mux2_1
XTAP_2179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14440_ _15301_/CLK _14440_/D vssd1 vssd1 vccd1 vccd1 _14440_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11652_ _13327_/A0 _15084_/Q _11670_/S vssd1 vssd1 vccd1 vccd1 _15084_/D sky130_fd_sc_hd__mux2_1
XTAP_1489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_920 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10603_ _15558_/Q _10731_/B _10733_/A2 _14967_/Q vssd1 vssd1 vccd1 vccd1 _10603_/X
+ sky130_fd_sc_hd__a22o_1
X_14371_ _15664_/CLK _14371_/D vssd1 vssd1 vccd1 vccd1 _14371_/Q sky130_fd_sc_hd__dfxtp_1
X_11583_ _11584_/A _11584_/B vssd1 vssd1 vccd1 vccd1 _11585_/A sky130_fd_sc_hd__and2_1
XFILLER_11_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13322_ _13322_/A0 _15652_/Q _13345_/S vssd1 vssd1 vccd1 vccd1 _15652_/D sky130_fd_sc_hd__mux2_1
X_10534_ _11600_/A _13236_/B _10532_/Y _10533_/X _10462_/A vssd1 vssd1 vccd1 vccd1
+ _10534_/X sky130_fd_sc_hd__o221a_1
XFILLER_182_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10465_ _08244_/A _13749_/Q _15423_/Q _08244_/B vssd1 vssd1 vccd1 vccd1 _10465_/X
+ sky130_fd_sc_hd__a22o_1
X_13253_ _11129_/B _13251_/X _13252_/Y _13252_/B _15584_/Q vssd1 vssd1 vccd1 vccd1
+ _15584_/D sky130_fd_sc_hd__a32o_1
XFILLER_182_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12204_ _12503_/A1 _12203_/X _12202_/X _12503_/C1 vssd1 vssd1 vccd1 vccd1 _12205_/C
+ sky130_fd_sc_hd__a211o_1
X_13184_ _13229_/A _13183_/B _11436_/B _13241_/A2 vssd1 vssd1 vccd1 vccd1 _13184_/X
+ sky130_fd_sc_hd__a211o_1
X_10396_ _08240_/A _13800_/Q _13768_/Q _08237_/A vssd1 vssd1 vccd1 vccd1 _10396_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_124_855 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12135_ _12503_/A1 _12134_/X _12133_/X _12503_/C1 vssd1 vssd1 vccd1 vccd1 _12136_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_111_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12066_ _12273_/A1 _12065_/X _12064_/X _12503_/C1 vssd1 vssd1 vccd1 vccd1 _12067_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_38_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11017_ _13217_/B _13215_/B _11025_/A vssd1 vssd1 vccd1 vccd1 _11017_/X sky130_fd_sc_hd__mux2_1
XFILLER_49_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_360 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12968_ _15469_/Q _13105_/A2 _13025_/B1 _12967_/X vssd1 vssd1 vccd1 vccd1 _15469_/D
+ sky130_fd_sc_hd__a22o_1
XTAP_3381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14707_ _14892_/CLK _14707_/D vssd1 vssd1 vccd1 vccd1 _14707_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_45_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11919_ _12383_/A _11919_/B vssd1 vssd1 vccd1 vccd1 _11919_/X sky130_fd_sc_hd__and2_1
XTAP_2680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12899_ _15427_/Q _15612_/Q _12910_/S vssd1 vssd1 vccd1 vccd1 _15427_/D sky130_fd_sc_hd__mux2_1
XTAP_2691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14638_ _15606_/CLK _14638_/D vssd1 vssd1 vccd1 vccd1 _14638_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14569_ _15292_/CLK _14569_/D vssd1 vssd1 vccd1 vccd1 _14569_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_159_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07110_ _14832_/Q _07115_/B _07163_/A vssd1 vssd1 vccd1 vccd1 _07110_/X sky130_fd_sc_hd__and3_4
XFILLER_146_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08090_ _08083_/A _08089_/Y input35/X vssd1 vssd1 vccd1 vccd1 _08090_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_173_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07041_ _07040_/X _14746_/Q _07077_/S vssd1 vssd1 vccd1 vccd1 _13592_/D sky130_fd_sc_hd__mux2_1
XFILLER_173_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_991 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08992_ _13911_/Q _08991_/X _12481_/A vssd1 vssd1 vccd1 vccd1 _13911_/D sky130_fd_sc_hd__mux2_1
XFILLER_173_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07943_ _13551_/Q _07943_/B vssd1 vssd1 vccd1 vccd1 _07943_/X sky130_fd_sc_hd__xor2_1
XFILLER_68_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07874_ _07874_/A _07874_/B vssd1 vssd1 vccd1 vccd1 _07874_/Y sky130_fd_sc_hd__nand2_1
XFILLER_68_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09613_ _13987_/Q _13335_/A0 _09627_/S vssd1 vssd1 vccd1 vccd1 _13987_/D sky130_fd_sc_hd__mux2_1
XFILLER_55_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06825_ _06819_/X _06825_/B _06825_/C _08085_/S vssd1 vssd1 vccd1 vccd1 _06825_/X
+ sky130_fd_sc_hd__and4b_4
XFILLER_83_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09544_ _13123_/A _09541_/X _09543_/X _09554_/A vssd1 vssd1 vccd1 vccd1 _09544_/X
+ sky130_fd_sc_hd__o211a_1
X_06756_ _13477_/Q vssd1 vssd1 vccd1 vccd1 _06756_/Y sky130_fd_sc_hd__inv_2
XFILLER_110_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_544 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09475_ _14384_/Q _15200_/Q _13839_/Q _14578_/Q _09551_/S _09550_/A1 vssd1 vssd1
+ vccd1 vccd1 _09476_/B sky130_fd_sc_hd__mux4_1
X_06687_ _15399_/Q vssd1 vssd1 vccd1 vccd1 _06687_/Y sky130_fd_sc_hd__inv_2
XFILLER_51_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08426_ _10764_/S _08426_/B vssd1 vssd1 vccd1 vccd1 _08426_/X sky130_fd_sc_hd__or2_4
XFILLER_180_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08357_ _08357_/A vssd1 vssd1 vccd1 vccd1 _08357_/Y sky130_fd_sc_hd__inv_2
XFILLER_138_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07308_ _07301_/Y _07302_/X _07306_/Y _07307_/X vssd1 vssd1 vccd1 vccd1 _07350_/C
+ sky130_fd_sc_hd__o22a_1
XFILLER_137_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08288_ _11041_/B _11044_/A vssd1 vssd1 vccd1 vccd1 _08288_/X sky130_fd_sc_hd__or2_1
XFILLER_152_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07239_ _13927_/Q _15514_/Q _07334_/S vssd1 vssd1 vccd1 vccd1 _07265_/A sky130_fd_sc_hd__mux2_8
XFILLER_180_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10250_ _14635_/Q _14788_/Q _10715_/S vssd1 vssd1 vccd1 vccd1 _14635_/D sky130_fd_sc_hd__mux2_1
XFILLER_180_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10181_ _13334_/A0 _14565_/Q _10192_/S vssd1 vssd1 vccd1 vccd1 _14565_/D sky130_fd_sc_hd__mux2_1
XFILLER_78_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout240 _12936_/X vssd1 vssd1 vccd1 vccd1 _13024_/B2 sky130_fd_sc_hd__buf_12
XFILLER_87_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout251 _08518_/Y vssd1 vssd1 vccd1 vccd1 _08746_/A2 sky130_fd_sc_hd__buf_12
Xfanout262 _06775_/Y vssd1 vssd1 vccd1 vccd1 _07193_/S sky130_fd_sc_hd__buf_12
X_13940_ _15077_/CLK _13940_/D vssd1 vssd1 vccd1 vccd1 _13940_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_93_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout273 _08503_/Y vssd1 vssd1 vccd1 vccd1 _08748_/A2 sky130_fd_sc_hd__buf_12
Xfanout284 _13349_/A0 vssd1 vssd1 vccd1 vccd1 _11816_/A1 sky130_fd_sc_hd__buf_6
XFILLER_75_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout295 _13344_/A0 vssd1 vssd1 vccd1 vccd1 _11877_/A1 sky130_fd_sc_hd__buf_6
X_13871_ _15200_/CLK _13871_/D vssd1 vssd1 vccd1 vccd1 _13871_/Q sky130_fd_sc_hd__dfxtp_1
X_15610_ _15645_/CLK _15610_/D vssd1 vssd1 vccd1 vccd1 _15610_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_28_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12822_ _15072_/Q _12834_/B vssd1 vssd1 vccd1 vccd1 _12822_/X sky130_fd_sc_hd__or2_1
XFILLER_28_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15541_ _15542_/CLK _15541_/D vssd1 vssd1 vccd1 vccd1 _15541_/Q sky130_fd_sc_hd__dfxtp_1
X_12753_ _15356_/Q _12754_/B vssd1 vssd1 vccd1 vccd1 _12767_/C sky130_fd_sc_hd__and2_2
XFILLER_188_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_847 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11704_ _13346_/A0 _15135_/Q _11708_/S vssd1 vssd1 vccd1 vccd1 _15135_/D sky130_fd_sc_hd__mux2_1
XFILLER_187_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15472_ _15520_/CLK _15472_/D vssd1 vssd1 vccd1 vccd1 _15472_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_188_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12684_ _13423_/Q _12683_/X _12728_/S vssd1 vssd1 vccd1 vccd1 _12685_/B sky130_fd_sc_hd__mux2_1
XTAP_1286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14423_ _14606_/CLK _14423_/D vssd1 vssd1 vccd1 vccd1 _14423_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11635_ _11635_/A _11635_/B vssd1 vssd1 vccd1 vccd1 _11635_/X sky130_fd_sc_hd__xor2_1
XFILLER_168_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14354_ _15303_/CLK _14354_/D vssd1 vssd1 vccd1 vccd1 _14354_/Q sky130_fd_sc_hd__dfxtp_1
X_11566_ _11576_/C _11567_/B vssd1 vssd1 vccd1 vccd1 _11566_/X sky130_fd_sc_hd__or2_1
XFILLER_128_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13305_ _15637_/Q _12761_/X _13316_/S vssd1 vssd1 vccd1 vccd1 _15637_/D sky130_fd_sc_hd__mux2_1
XFILLER_6_231 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_788 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10517_ _11536_/C _11521_/A vssd1 vssd1 vccd1 vccd1 _10519_/A sky130_fd_sc_hd__nor2_1
XFILLER_6_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14285_ _15662_/CLK _14285_/D vssd1 vssd1 vccd1 vccd1 _14285_/Q sky130_fd_sc_hd__dfxtp_1
X_11497_ _13236_/A _11537_/A vssd1 vssd1 vccd1 vccd1 _11498_/B sky130_fd_sc_hd__or2_1
XFILLER_157_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13236_ _13236_/A _13236_/B vssd1 vssd1 vccd1 vccd1 _13236_/Y sky130_fd_sc_hd__nor2_1
XFILLER_143_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10448_ _11600_/A _13236_/B vssd1 vssd1 vccd1 vccd1 _10470_/A sky130_fd_sc_hd__xnor2_2
XFILLER_170_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_663 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13167_ _15556_/Q _13252_/B _13165_/Y _13166_/X vssd1 vssd1 vccd1 vccd1 _15556_/D
+ sky130_fd_sc_hd__a22o_1
X_10379_ _11457_/A _11475_/B vssd1 vssd1 vccd1 vccd1 _10379_/Y sky130_fd_sc_hd__nor2_1
XFILLER_152_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12118_ _15118_/Q _15086_/Q _15659_/Q _13393_/Q _12472_/S _12465_/S1 vssd1 vssd1
+ vccd1 vccd1 _12118_/X sky130_fd_sc_hd__mux4_1
X_13098_ _13014_/X _13118_/A2 _13114_/B1 _13098_/B2 vssd1 vssd1 vccd1 vccd1 _13098_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_85_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12049_ _15115_/Q _15083_/Q _15656_/Q _13390_/Q _12246_/S _12452_/A vssd1 vssd1 vccd1
+ vccd1 _12049_/X sky130_fd_sc_hd__mux4_1
XFILLER_133_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07590_ _14747_/Q _07607_/A _07589_/Y _12809_/C1 vssd1 vssd1 vccd1 vccd1 _13458_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_92_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09260_ _14374_/Q _15190_/Q _13829_/Q _14568_/Q _09481_/S _08519_/A vssd1 vssd1 vccd1
+ vccd1 _09261_/B sky130_fd_sc_hd__mux4_1
XFILLER_178_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08211_ _13702_/Q _11873_/A1 _08221_/S vssd1 vssd1 vccd1 vccd1 _13702_/D sky130_fd_sc_hd__mux2_1
X_09191_ _13889_/Q _09231_/A2 _09403_/B1 _14404_/Q _09437_/A1 vssd1 vssd1 vccd1 vccd1
+ _09191_/X sky130_fd_sc_hd__a221o_1
XFILLER_21_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08142_ _08133_/S _06764_/Y _08093_/B vssd1 vssd1 vccd1 vccd1 _08142_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_119_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_563 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08073_ _15648_/Q _13644_/Q _08085_/S vssd1 vssd1 vccd1 vccd1 _08075_/B sky130_fd_sc_hd__mux2_1
XFILLER_162_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07024_ _14620_/Q _14652_/Q _07096_/S vssd1 vssd1 vccd1 vccd1 _07024_/X sky130_fd_sc_hd__mux2_1
XFILLER_143_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_919 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08975_ _09445_/C1 _08972_/X _08974_/X _09130_/A vssd1 vssd1 vccd1 vccd1 _08975_/X
+ sky130_fd_sc_hd__o211a_1
X_07926_ _07935_/D _07925_/Y _08012_/A2 vssd1 vssd1 vccd1 vccd1 _07926_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_152_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07857_ _14753_/Q _07874_/A _07856_/Y vssd1 vssd1 vccd1 vccd1 _13528_/D sky130_fd_sc_hd__o21a_1
XFILLER_29_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06808_ _14588_/Q _14587_/Q _08392_/B vssd1 vssd1 vccd1 vccd1 _06808_/X sky130_fd_sc_hd__and3_2
XFILLER_16_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07788_ _13510_/Q _07779_/X _07802_/C vssd1 vssd1 vccd1 vccd1 _07789_/B sky130_fd_sc_hd__o21bai_1
XFILLER_71_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09527_ _15138_/Q _09558_/A2 _08520_/B _09526_/X vssd1 vssd1 vccd1 vccd1 _09527_/X
+ sky130_fd_sc_hd__a22o_1
X_06739_ _13452_/Q vssd1 vssd1 vccd1 vccd1 _06739_/Y sky130_fd_sc_hd__inv_2
XFILLER_36_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09458_ _14094_/Q _13123_/B _08512_/B _14062_/Q _09466_/A vssd1 vssd1 vccd1 vccd1
+ _09458_/X sky130_fd_sc_hd__a221o_1
XFILLER_80_992 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08409_ _08756_/B _06833_/X _08777_/A _13129_/A _13738_/Q vssd1 vssd1 vccd1 vccd1
+ _13738_/D sky130_fd_sc_hd__a32o_1
XFILLER_169_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09389_ _13930_/Q _09388_/X _10868_/S vssd1 vssd1 vccd1 vccd1 _13930_/D sky130_fd_sc_hd__mux2_1
XFILLER_8_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11420_ _11420_/A _11420_/B vssd1 vssd1 vccd1 vccd1 _11460_/D sky130_fd_sc_hd__and2_1
XFILLER_138_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11351_ _11048_/Y _11325_/X _11348_/Y _11350_/X _11351_/C1 vssd1 vssd1 vccd1 vccd1
+ _11351_/X sky130_fd_sc_hd__o221a_1
XFILLER_126_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10302_ _14687_/Q _14872_/Q _10710_/S vssd1 vssd1 vccd1 vccd1 _14687_/D sky130_fd_sc_hd__mux2_1
X_14070_ _15244_/CLK _14070_/D vssd1 vssd1 vccd1 vccd1 _14070_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_125_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11282_ _11251_/Y _11281_/Y _11297_/S vssd1 vssd1 vccd1 vccd1 _11282_/X sky130_fd_sc_hd__mux2_1
XFILLER_4_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_768 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13021_ _13344_/A0 _13024_/A2 _13020_/X _13024_/B2 vssd1 vssd1 vccd1 vccd1 _13021_/X
+ sky130_fd_sc_hd__a22o_1
X_10233_ _14618_/Q _14771_/Q _10615_/S vssd1 vssd1 vccd1 vccd1 _14618_/D sky130_fd_sc_hd__mux2_1
XFILLER_106_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10164_ _14549_/Q _11883_/A1 _10164_/S vssd1 vssd1 vccd1 vccd1 _14549_/D sky130_fd_sc_hd__mux2_1
XFILLER_117_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_1079 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14972_ _14988_/CLK _14972_/D vssd1 vssd1 vccd1 vccd1 _14972_/Q sky130_fd_sc_hd__dfxtp_1
X_10095_ _14451_/Q _13110_/B2 _10097_/S vssd1 vssd1 vccd1 vccd1 _14451_/D sky130_fd_sc_hd__mux2_1
XFILLER_120_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13923_ _15212_/CLK _13923_/D vssd1 vssd1 vccd1 vccd1 _13923_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_48_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_210_clk clkbuf_5_16_0_clk/X vssd1 vssd1 vccd1 vccd1 _15678_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_90_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13854_ _15663_/CLK _13854_/D vssd1 vssd1 vccd1 vccd1 _13854_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_142_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_5_9_0_clk clkbuf_5_9_0_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_5_9_0_clk/X sky130_fd_sc_hd__clkbuf_8
X_12805_ _12828_/A _12805_/B vssd1 vssd1 vccd1 vccd1 _12805_/X sky130_fd_sc_hd__or2_1
XFILLER_34_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13785_ _14495_/CLK _13785_/D vssd1 vssd1 vccd1 vccd1 _13785_/Q sky130_fd_sc_hd__dfxtp_4
X_10997_ _11088_/S _11349_/B _13159_/B _10403_/A _11362_/B vssd1 vssd1 vccd1 vccd1
+ _10997_/X sky130_fd_sc_hd__a311o_1
X_15524_ _15673_/CLK _15524_/D vssd1 vssd1 vccd1 vccd1 _15524_/Q sky130_fd_sc_hd__dfxtp_1
X_12736_ _13430_/Q _12735_/X _12764_/S vssd1 vssd1 vccd1 vccd1 _12737_/B sky130_fd_sc_hd__mux2_1
XTAP_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15455_ _15641_/CLK _15455_/D vssd1 vssd1 vccd1 vccd1 hold9/A sky130_fd_sc_hd__dfxtp_1
XFILLER_188_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12667_ _12679_/C _12667_/B vssd1 vssd1 vccd1 vccd1 _12667_/Y sky130_fd_sc_hd__nor2_1
XFILLER_169_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14406_ _15665_/CLK _14406_/D vssd1 vssd1 vccd1 vccd1 _14406_/Q sky130_fd_sc_hd__dfxtp_1
X_11618_ _13242_/B _11618_/B vssd1 vssd1 vccd1 vccd1 _11621_/A sky130_fd_sc_hd__xor2_2
X_15386_ _15386_/CLK _15386_/D vssd1 vssd1 vccd1 vccd1 _15386_/Q sky130_fd_sc_hd__dfxtp_1
X_12598_ _14259_/Q _14291_/Q _14323_/Q _14355_/Q _12518_/S _12383_/A vssd1 vssd1 vccd1
+ vccd1 _12598_/X sky130_fd_sc_hd__mux4_1
X_14337_ _15298_/CLK _14337_/D vssd1 vssd1 vccd1 vccd1 _14337_/Q sky130_fd_sc_hd__dfxtp_1
X_11549_ _11576_/A _11549_/B vssd1 vssd1 vccd1 vccd1 _11549_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_143_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14268_ _15279_/CLK _14268_/D vssd1 vssd1 vccd1 vccd1 _14268_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_143_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_1072 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13219_ _15573_/Q _13218_/Y _13219_/S vssd1 vssd1 vccd1 vccd1 _15573_/D sky130_fd_sc_hd__mux2_1
X_14199_ _15244_/CLK _14199_/D vssd1 vssd1 vccd1 vccd1 _14199_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_1078 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_1_1_clk clkbuf_1_1_1_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_2_3_0_clk/A sky130_fd_sc_hd__clkbuf_8
XTAP_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08760_ _14608_/Q _14610_/Q _14609_/Q _14614_/Q vssd1 vssd1 vccd1 vccd1 _08772_/A
+ sky130_fd_sc_hd__or4_1
XFILLER_112_688 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07711_ _14747_/Q _07713_/A _07710_/Y _07949_/C1 vssd1 vssd1 vccd1 vccd1 _13490_/D
+ sky130_fd_sc_hd__o211a_1
X_08691_ _13588_/Q _08691_/A2 _08691_/B1 _13485_/Q _08540_/X vssd1 vssd1 vccd1 vccd1
+ _08691_/X sky130_fd_sc_hd__a221o_1
XFILLER_39_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_201_clk clkbuf_5_17_0_clk/X vssd1 vssd1 vccd1 vccd1 _15278_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_38_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07642_ _14761_/Q _07651_/A _07641_/Y _08012_/C1 vssd1 vssd1 vccd1 vccd1 _13472_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_38_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07573_ _07570_/X _07575_/B _07629_/A vssd1 vssd1 vccd1 vccd1 _07573_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_18_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09312_ _13895_/Q _09522_/A2 _09519_/B1 _14410_/Q _08507_/A vssd1 vssd1 vccd1 vccd1
+ _09312_/X sky130_fd_sc_hd__a221o_1
XFILLER_62_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09243_ _14245_/Q _14277_/Q _14309_/Q _14341_/Q _09557_/S _09550_/A1 vssd1 vssd1
+ vccd1 vccd1 _09243_/X sky130_fd_sc_hd__mux4_1
XFILLER_178_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09174_ _15662_/Q _13396_/Q _09444_/S vssd1 vssd1 vccd1 vccd1 _09174_/X sky130_fd_sc_hd__mux2_1
XFILLER_21_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08125_ input32/X input9/X _08133_/S vssd1 vssd1 vccd1 vccd1 _08125_/X sky130_fd_sc_hd__mux2_1
XFILLER_179_1040 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_162_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08056_ _14749_/Q _13627_/Q _08066_/S vssd1 vssd1 vccd1 vccd1 _13627_/D sky130_fd_sc_hd__mux2_1
XFILLER_162_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07007_ _14646_/Q _13581_/Q _12640_/S vssd1 vssd1 vccd1 vccd1 _07007_/X sky130_fd_sc_hd__mux2_1
XFILLER_103_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput38 _07174_/X vssd1 vssd1 vccd1 vccd1 ext_address[12] sky130_fd_sc_hd__clkbuf_2
Xoutput49 _07185_/X vssd1 vssd1 vccd1 vccd1 ext_address[23] sky130_fd_sc_hd__clkbuf_2
XFILLER_163_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08958_ _14457_/Q _09536_/A2 _08957_/X _06676_/A vssd1 vssd1 vccd1 vccd1 _08958_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_56_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07909_ _14734_/Q _08022_/B _07908_/X _08016_/C1 vssd1 vssd1 vccd1 vccd1 _13541_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_3914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08889_ _09445_/C1 _08888_/X _08887_/X _09130_/A vssd1 vssd1 vccd1 vccd1 _08889_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_57_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_1011 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10920_ _13195_/B _10944_/B vssd1 vssd1 vccd1 vccd1 _10920_/Y sky130_fd_sc_hd__nand2_1
XFILLER_5_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10851_ _14883_/Q _13785_/Q _12933_/S vssd1 vssd1 vccd1 vccd1 _14883_/D sky130_fd_sc_hd__mux2_1
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_96 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13570_ _13642_/CLK _13570_/D vssd1 vssd1 vccd1 vccd1 _13570_/Q sky130_fd_sc_hd__dfxtp_1
X_10782_ _14814_/Q _15446_/Q _12917_/S vssd1 vssd1 vccd1 vccd1 _14814_/D sky130_fd_sc_hd__mux2_1
XFILLER_169_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12521_ _12521_/A _12521_/B vssd1 vssd1 vccd1 vccd1 _12521_/X sky130_fd_sc_hd__and2_1
XPHY_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_636 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15240_ _15304_/CLK _15240_/D vssd1 vssd1 vccd1 vccd1 _15240_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12452_ _12452_/A _12452_/B vssd1 vssd1 vccd1 vccd1 _12452_/X sky130_fd_sc_hd__and2_1
XFILLER_185_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11403_ _11386_/B _11423_/C _11402_/Y vssd1 vssd1 vccd1 vccd1 _11404_/B sky130_fd_sc_hd__a21oi_2
X_15171_ _15304_/CLK _15171_/D vssd1 vssd1 vccd1 vccd1 _15171_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_153_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12383_ _12383_/A _12383_/B vssd1 vssd1 vccd1 vccd1 _12383_/X sky130_fd_sc_hd__and2_1
XFILLER_165_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14122_ _15336_/CLK _14122_/D vssd1 vssd1 vccd1 vccd1 _14122_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_181_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11334_ _08233_/B _08359_/X _11329_/Y _11333_/X wire438/X vssd1 vssd1 vccd1 vccd1
+ _11334_/X sky130_fd_sc_hd__o221a_1
XFILLER_141_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14053_ _14373_/CLK _14053_/D vssd1 vssd1 vccd1 vccd1 _14053_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_125_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11265_ _11037_/A _13215_/B _11020_/A vssd1 vssd1 vccd1 vccd1 _11265_/X sky130_fd_sc_hd__o21ba_1
XFILLER_107_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13004_ _15481_/Q _13093_/A2 _13116_/C _13003_/X vssd1 vssd1 vccd1 vccd1 _15481_/D
+ sky130_fd_sc_hd__a22o_1
X_10216_ input10/X _08451_/A _13284_/S vssd1 vssd1 vccd1 vccd1 _14601_/D sky130_fd_sc_hd__mux2_1
XFILLER_97_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11196_ _14990_/Q _11164_/S _11170_/X _11195_/Y vssd1 vssd1 vccd1 vccd1 _14990_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_39_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10147_ _14532_/Q _13333_/A0 _10159_/S vssd1 vssd1 vccd1 vccd1 _14532_/D sky130_fd_sc_hd__mux2_1
X_14955_ _15021_/CLK _14955_/D vssd1 vssd1 vccd1 vccd1 _14955_/Q sky130_fd_sc_hd__dfxtp_1
X_10078_ _14434_/Q _11689_/A0 _10092_/S vssd1 vssd1 vccd1 vccd1 _14434_/D sky130_fd_sc_hd__mux2_1
X_13906_ _15326_/CLK _13906_/D vssd1 vssd1 vccd1 vccd1 _13906_/Q sky130_fd_sc_hd__dfxtp_1
X_14886_ _15607_/CLK _14886_/D vssd1 vssd1 vccd1 vccd1 _14886_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_130_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_436 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13837_ _15267_/CLK _13837_/D vssd1 vssd1 vccd1 vccd1 _13837_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13768_ _15589_/CLK _13768_/D vssd1 vssd1 vccd1 vccd1 _13768_/Q sky130_fd_sc_hd__dfxtp_1
X_12719_ _13595_/Q _12718_/X _12785_/B vssd1 vssd1 vccd1 vccd1 _12719_/X sky130_fd_sc_hd__mux2_1
X_15507_ _15507_/CLK _15507_/D vssd1 vssd1 vccd1 vccd1 _15507_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0_clk clk vssd1 vssd1 vccd1 vccd1 clkbuf_0_clk/X sky130_fd_sc_hd__clkbuf_16
XFILLER_30_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13699_ _15094_/CLK _13699_/D vssd1 vssd1 vccd1 vccd1 _13699_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_175_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15438_ _15438_/CLK _15438_/D vssd1 vssd1 vccd1 vccd1 _15438_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_164_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15369_ _15372_/CLK _15369_/D vssd1 vssd1 vccd1 vccd1 _15369_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_157_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_511 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09930_ _13350_/A0 _14291_/Q _09930_/S vssd1 vssd1 vccd1 vccd1 _14291_/D sky130_fd_sc_hd__mux2_1
XFILLER_98_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09861_ _14225_/Q _13110_/B2 _09863_/S vssd1 vssd1 vccd1 vccd1 _14225_/D sky130_fd_sc_hd__mux2_1
XFILLER_98_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08812_ _11879_/A1 _13838_/Q _08816_/S vssd1 vssd1 vccd1 vccd1 _13838_/D sky130_fd_sc_hd__mux2_1
XTAP_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09792_ _14159_/Q _13347_/A0 _09795_/S vssd1 vssd1 vccd1 vccd1 _14159_/D sky130_fd_sc_hd__mux2_1
XTAP_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08743_ _13581_/Q _08749_/A2 _08538_/Y _15369_/Q vssd1 vssd1 vccd1 vccd1 _08743_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_39_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08674_ _13575_/Q _08667_/X _08671_/X _08673_/X _08722_/A vssd1 vssd1 vccd1 vccd1
+ _08674_/X sky130_fd_sc_hd__a2111o_1
X_07625_ _13468_/Q _07625_/B vssd1 vssd1 vccd1 vccd1 _07655_/A sky130_fd_sc_hd__and2_2
XTAP_1808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07556_ _13449_/Q _07559_/D _13450_/Q vssd1 vssd1 vccd1 vccd1 _07556_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_167_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07487_ _13677_/Q _07499_/A2 _07499_/B1 _14705_/Q _07486_/X vssd1 vssd1 vccd1 vccd1
+ _07487_/X sky130_fd_sc_hd__a221o_1
XFILLER_158_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09226_ _09449_/A1 _09224_/X _09225_/X _09449_/B2 _09223_/X vssd1 vssd1 vccd1 vccd1
+ _09226_/X sky130_fd_sc_hd__a221o_1
XFILLER_167_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_166_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_628 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09157_ _09155_/X _09156_/X _12596_/A _09146_/X vssd1 vssd1 vccd1 vccd1 _09157_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_107_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08108_ input27/X input4/X input13/X input21/X _08150_/S _08151_/S vssd1 vssd1 vccd1
+ vccd1 _08108_/X sky130_fd_sc_hd__mux4_1
XFILLER_181_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09088_ _09427_/A1 _09086_/X _09087_/X vssd1 vssd1 vccd1 vccd1 _09088_/X sky130_fd_sc_hd__a21o_1
XFILLER_135_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08039_ _13579_/Q _14741_/Q _08039_/S vssd1 vssd1 vccd1 vccd1 _13579_/D sky130_fd_sc_hd__mux2_1
XFILLER_150_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11050_ _11380_/A _11050_/B vssd1 vssd1 vccd1 vccd1 _11050_/Y sky130_fd_sc_hd__nor2_1
XFILLER_115_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10001_ _13322_/A0 _14359_/Q _10028_/S vssd1 vssd1 vccd1 vccd1 _14359_/D sky130_fd_sc_hd__mux2_1
XFILLER_131_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_1087 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14740_ _14892_/CLK _14740_/D vssd1 vssd1 vccd1 vccd1 _14740_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_3744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11952_ _12573_/A _11952_/B _11952_/C vssd1 vssd1 vccd1 vccd1 _11952_/X sky130_fd_sc_hd__and3_2
XFILLER_85_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10903_ _14934_/Q _10951_/B _10902_/Y _13168_/B vssd1 vssd1 vccd1 vccd1 _14934_/D
+ sky130_fd_sc_hd__o22a_1
XTAP_3788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14671_ _15453_/CLK _14671_/D vssd1 vssd1 vccd1 vccd1 _14671_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11883_ _15304_/Q _11883_/A1 _11883_/S vssd1 vssd1 vccd1 vccd1 _15304_/D sky130_fd_sc_hd__mux2_1
X_13622_ _15378_/CLK _13622_/D vssd1 vssd1 vccd1 vccd1 _13622_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_60 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10834_ _13802_/Q _14866_/Q _10834_/S vssd1 vssd1 vccd1 vccd1 _14866_/D sky130_fd_sc_hd__mux2_1
X_13553_ _13627_/CLK _13553_/D vssd1 vssd1 vccd1 vccd1 _13553_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_158_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10765_ _15429_/Q _14797_/Q _10765_/S vssd1 vssd1 vccd1 vccd1 _14797_/D sky130_fd_sc_hd__mux2_1
XFILLER_12_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_956 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12504_ _12504_/A _12504_/B _12504_/C vssd1 vssd1 vccd1 vccd1 _12504_/X sky130_fd_sc_hd__and3_1
XFILLER_160_1047 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13484_ _13798_/CLK _13484_/D vssd1 vssd1 vccd1 vccd1 _13484_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_186_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10696_ _15577_/Q _10731_/B vssd1 vssd1 vccd1 vccd1 _10696_/X sky130_fd_sc_hd__and2_1
XFILLER_173_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15223_ _15287_/CLK _15223_/D vssd1 vssd1 vccd1 vccd1 _15223_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_173_628 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12435_ _12573_/A _12435_/B _12435_/C vssd1 vssd1 vccd1 vccd1 _12435_/X sky130_fd_sc_hd__and3_1
XFILLER_139_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15154_ _15287_/CLK _15154_/D vssd1 vssd1 vccd1 vccd1 _15154_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_126_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12366_ _12573_/A _12366_/B _12366_/C vssd1 vssd1 vccd1 vccd1 _12366_/X sky130_fd_sc_hd__and3_1
XFILLER_5_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14105_ _14462_/CLK _14105_/D vssd1 vssd1 vccd1 vccd1 _14105_/Q sky130_fd_sc_hd__dfxtp_1
X_11317_ _11317_/A _11317_/B vssd1 vssd1 vccd1 vccd1 _11330_/B sky130_fd_sc_hd__nor2_1
XFILLER_153_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15085_ _15658_/CLK _15085_/D vssd1 vssd1 vccd1 vccd1 _15085_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12297_ _12320_/A _12297_/B _12297_/C vssd1 vssd1 vccd1 vccd1 _12297_/X sky130_fd_sc_hd__and3_1
XFILLER_141_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14036_ _15125_/CLK _14036_/D vssd1 vssd1 vccd1 vccd1 _14036_/Q sky130_fd_sc_hd__dfxtp_1
X_11248_ _15027_/Q wire438/A _11246_/X _11247_/X vssd1 vssd1 vccd1 vccd1 _15027_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_80_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11179_ _11199_/A _11179_/B vssd1 vssd1 vccd1 vccd1 _11179_/Y sky130_fd_sc_hd__nor2_1
XFILLER_80_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14938_ _15006_/CLK _14938_/D vssd1 vssd1 vccd1 vccd1 _14938_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_1083 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14869_ _15589_/CLK _14869_/D vssd1 vssd1 vccd1 vccd1 _14869_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07410_ _14654_/Q _07474_/B _07482_/C vssd1 vssd1 vccd1 vccd1 _07410_/X sky130_fd_sc_hd__and3_1
XFILLER_35_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08390_ _08390_/A _08390_/B _08390_/C vssd1 vssd1 vccd1 vccd1 _08390_/X sky130_fd_sc_hd__or3_2
XFILLER_35_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07341_ _07341_/A vssd1 vssd1 vccd1 vccd1 _07341_/Y sky130_fd_sc_hd__inv_2
X_07272_ _07235_/A _07235_/B _07237_/Y _07238_/X _07268_/B vssd1 vssd1 vccd1 vccd1
+ _07273_/D sky130_fd_sc_hd__o221a_1
XFILLER_176_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09011_ _15113_/Q _09558_/A2 _13130_/C1 _09010_/X vssd1 vssd1 vccd1 vccd1 _09011_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_12_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09913_ _13080_/B2 _14274_/Q _09925_/S vssd1 vssd1 vccd1 vccd1 _14274_/D sky130_fd_sc_hd__mux2_1
Xfanout603 _12470_/S vssd1 vssd1 vccd1 vccd1 _12154_/S sky130_fd_sc_hd__buf_12
Xfanout614 _14598_/Q vssd1 vssd1 vccd1 vccd1 _08457_/A sky130_fd_sc_hd__buf_12
Xfanout625 _08405_/A vssd1 vssd1 vccd1 vccd1 _12518_/S sky130_fd_sc_hd__buf_6
Xfanout636 fanout647/X vssd1 vssd1 vccd1 vccd1 _12809_/C1 sky130_fd_sc_hd__clkbuf_16
XFILLER_101_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09844_ _14208_/Q _11689_/A0 _09858_/S vssd1 vssd1 vccd1 vccd1 _14208_/D sky130_fd_sc_hd__mux2_1
Xfanout647 _06684_/Y vssd1 vssd1 vccd1 vccd1 fanout647/X sky130_fd_sc_hd__buf_12
XFILLER_85_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09775_ _14142_/Q _13074_/B2 _09790_/S vssd1 vssd1 vccd1 vccd1 _14142_/D sky130_fd_sc_hd__mux2_1
XFILLER_85_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06987_ _14586_/Q _14589_/Q _14587_/Q _06987_/D vssd1 vssd1 vccd1 vccd1 _08390_/C
+ sky130_fd_sc_hd__and4bb_4
XTAP_3007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08726_ _13615_/Q _08750_/B1 _08535_/X _13416_/Q _08725_/X vssd1 vssd1 vccd1 vccd1
+ _08726_/X sky130_fd_sc_hd__a221o_1
XTAP_3029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08657_ _13490_/Q _08691_/B1 _08693_/B1 _13625_/Q vssd1 vssd1 vccd1 vccd1 _08657_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_1605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1036 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07608_ _14752_/Q _07607_/A _07607_/Y _07987_/C1 vssd1 vssd1 vccd1 vccd1 _13463_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_1638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_36 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08588_ _13532_/Q _08683_/A2 _08693_/B1 _13635_/Q _08587_/X vssd1 vssd1 vccd1 vccd1
+ _08588_/X sky130_fd_sc_hd__a221o_1
XFILLER_41_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07539_ _13445_/Q _07644_/A vssd1 vssd1 vccd1 vccd1 _07539_/Y sky130_fd_sc_hd__nand2_1
XFILLER_23_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10550_ _11362_/B _13162_/B vssd1 vssd1 vccd1 vccd1 _10556_/C sky130_fd_sc_hd__xnor2_1
XFILLER_183_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09209_ _14018_/Q _13986_/Q _09407_/S vssd1 vssd1 vccd1 vccd1 _09209_/X sky130_fd_sc_hd__mux2_1
XFILLER_185_13 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_627 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10481_ _10481_/A _10481_/B vssd1 vssd1 vccd1 vccd1 _10483_/A sky130_fd_sc_hd__and2_2
XFILLER_120_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12220_ _12477_/A1 _12219_/X _12168_/A vssd1 vssd1 vccd1 vccd1 _12220_/X sky130_fd_sc_hd__a21o_1
XFILLER_108_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12151_ _12500_/A1 _12150_/X _12582_/A vssd1 vssd1 vccd1 vccd1 _12151_/X sky130_fd_sc_hd__a21o_1
X_11102_ _14966_/Q _10984_/Y _11101_/X vssd1 vssd1 vccd1 vccd1 _14966_/D sky130_fd_sc_hd__a21bo_1
XFILLER_123_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12082_ _12500_/A1 _12081_/X _12582_/A vssd1 vssd1 vccd1 vccd1 _12082_/X sky130_fd_sc_hd__a21o_1
XFILLER_111_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11033_ _11033_/A _11033_/B vssd1 vssd1 vccd1 vccd1 _11033_/Y sky130_fd_sc_hd__nor2_1
XFILLER_77_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12984_ _10644_/X _14875_/Q _13029_/S vssd1 vssd1 vccd1 vccd1 _12984_/X sky130_fd_sc_hd__mux2_8
XTAP_3530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11935_ _11931_/X _11932_/X _12536_/A vssd1 vssd1 vccd1 vccd1 _11935_/X sky130_fd_sc_hd__mux2_1
X_14723_ _15548_/CLK _14723_/D vssd1 vssd1 vccd1 vccd1 _14723_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_3574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_60 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_715 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14654_ _15626_/CLK _14654_/D vssd1 vssd1 vccd1 vccd1 _14654_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11866_ _15287_/Q _13080_/B2 _11878_/S vssd1 vssd1 vccd1 vccd1 _15287_/D sky130_fd_sc_hd__mux2_1
XTAP_2884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13605_ _15375_/CLK _13605_/D vssd1 vssd1 vccd1 vccd1 _13605_/Q sky130_fd_sc_hd__dfxtp_2
X_10817_ _14849_/Q _07264_/A _10868_/S vssd1 vssd1 vccd1 vccd1 _14849_/D sky130_fd_sc_hd__mux2_1
X_14585_ _15537_/CLK _14585_/D vssd1 vssd1 vccd1 vccd1 _14585_/Q sky130_fd_sc_hd__dfxtp_1
X_11797_ _15220_/Q _13330_/A0 _11816_/S vssd1 vssd1 vccd1 vccd1 _15220_/D sky130_fd_sc_hd__mux2_1
XFILLER_60_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13536_ _14511_/CLK _13536_/D vssd1 vssd1 vccd1 vccd1 _13536_/Q sky130_fd_sc_hd__dfxtp_1
X_10748_ _15412_/Q _14780_/Q _10759_/S vssd1 vssd1 vccd1 vccd1 _14780_/D sky130_fd_sc_hd__mux2_1
XFILLER_158_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13467_ _14510_/CLK _13467_/D vssd1 vssd1 vccd1 vccd1 _13467_/Q sky130_fd_sc_hd__dfxtp_1
X_10679_ _15063_/Q _10714_/A2 _10676_/X _10678_/X vssd1 vssd1 vccd1 vccd1 _10679_/X
+ sky130_fd_sc_hd__o22a_4
XFILLER_173_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15206_ _15208_/CLK _15206_/D vssd1 vssd1 vccd1 vccd1 _15206_/Q sky130_fd_sc_hd__dfxtp_1
X_12418_ _12414_/X _12415_/X _12559_/A vssd1 vssd1 vccd1 vccd1 _12418_/X sky130_fd_sc_hd__mux2_1
X_13398_ _15664_/CLK _13398_/D vssd1 vssd1 vccd1 vccd1 _13398_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_182_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15137_ _15226_/CLK _15137_/D vssd1 vssd1 vccd1 vccd1 _15137_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12349_ _12345_/X _12346_/X _12536_/A vssd1 vssd1 vccd1 vccd1 _12349_/X sky130_fd_sc_hd__mux2_1
XFILLER_99_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15068_ _15572_/CLK _15068_/D vssd1 vssd1 vccd1 vccd1 _15068_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_4_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06910_ _06894_/X _06909_/X _06910_/S vssd1 vssd1 vccd1 vccd1 _06923_/A sky130_fd_sc_hd__mux2_1
X_14019_ _14083_/CLK _14019_/D vssd1 vssd1 vccd1 vccd1 _14019_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07890_ _07903_/A _07890_/B vssd1 vssd1 vccd1 vccd1 _07890_/Y sky130_fd_sc_hd__nand2_1
XFILLER_68_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06841_ _08405_/C _06834_/B _06681_/Y _12515_/C1 vssd1 vssd1 vccd1 vccd1 _06841_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_96_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09560_ _09544_/X _09547_/X _09554_/X _09559_/X vssd1 vssd1 vccd1 vccd1 _09560_/X
+ sky130_fd_sc_hd__o22a_2
X_06772_ _08150_/S _08121_/A _08185_/A _06661_/Y vssd1 vssd1 vccd1 vccd1 _10561_/B
+ sky130_fd_sc_hd__o2bb2a_4
XFILLER_167_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08511_ _08668_/C _13125_/A vssd1 vssd1 vccd1 vccd1 _08511_/Y sky130_fd_sc_hd__nor2_2
X_09491_ _15136_/Q _09558_/A2 _13130_/C1 _09490_/X vssd1 vssd1 vccd1 vccd1 _09491_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_70_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08442_ _13751_/Q _12878_/S _08426_/X _08441_/X vssd1 vssd1 vccd1 vccd1 _13751_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_169_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08373_ _07281_/X _10523_/A2 _08372_/X vssd1 vssd1 vccd1 vccd1 _13199_/B sky130_fd_sc_hd__a21oi_4
XFILLER_51_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07324_ _07324_/A vssd1 vssd1 vccd1 vccd1 _07324_/Y sky130_fd_sc_hd__inv_2
XFILLER_176_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07255_ _10481_/A vssd1 vssd1 vccd1 vccd1 _07261_/B sky130_fd_sc_hd__inv_2
XFILLER_118_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07186_ _15360_/Q _15067_/Q _07188_/S vssd1 vssd1 vccd1 vccd1 _07186_/X sky130_fd_sc_hd__mux2_4
XFILLER_117_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_2_2_0_clk clkbuf_2_3_0_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_2_2_1_clk/A sky130_fd_sc_hd__clkbuf_8
Xfanout400 _12662_/S vssd1 vssd1 vccd1 vccd1 _12640_/S sky130_fd_sc_hd__buf_12
Xfanout411 _11204_/X vssd1 vssd1 vccd1 vccd1 _11237_/S sky130_fd_sc_hd__buf_12
Xfanout422 _10569_/B vssd1 vssd1 vccd1 vccd1 _10717_/A2 sky130_fd_sc_hd__clkbuf_16
Xfanout433 _10457_/A2 vssd1 vssd1 vccd1 vccd1 _10360_/B sky130_fd_sc_hd__buf_12
XFILLER_171_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout444 _07372_/X vssd1 vssd1 vccd1 vccd1 _07499_/A2 sky130_fd_sc_hd__buf_12
XFILLER_150_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout455 _10244_/S vssd1 vssd1 vccd1 vccd1 _10343_/S sky130_fd_sc_hd__buf_12
Xfanout466 _12503_/C1 vssd1 vssd1 vccd1 vccd1 _12618_/C1 sky130_fd_sc_hd__buf_12
XFILLER_58_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09827_ _14193_/Q _11816_/A1 _09828_/S vssd1 vssd1 vccd1 vccd1 _14193_/D sky130_fd_sc_hd__mux2_1
Xfanout477 _12548_/S vssd1 vssd1 vccd1 vccd1 _12594_/S sky130_fd_sc_hd__buf_12
XFILLER_100_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_1098 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout488 _15526_/Q vssd1 vssd1 vccd1 vccd1 _07340_/S sky130_fd_sc_hd__buf_12
XFILLER_46_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout499 _14903_/Q vssd1 vssd1 vccd1 vccd1 _13038_/S sky130_fd_sc_hd__buf_12
XFILLER_58_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09758_ _14126_/Q _13346_/A0 _09762_/S vssd1 vssd1 vccd1 vccd1 _14126_/D sky130_fd_sc_hd__mux2_1
XFILLER_64_13 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_64 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08709_ _08722_/A _08709_/B _08709_/C vssd1 vssd1 vccd1 vccd1 _08709_/X sky130_fd_sc_hd__or3_4
XTAP_2125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09689_ _14060_/Q _13344_/A0 _09690_/S vssd1 vssd1 vccd1 vccd1 _14060_/D sky130_fd_sc_hd__mux2_1
XFILLER_73_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11720_ _15149_/Q _11861_/A1 _11741_/S vssd1 vssd1 vccd1 vccd1 _15149_/D sky130_fd_sc_hd__mux2_1
XFILLER_82_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11651_ _13326_/A0 _15083_/Q _11670_/S vssd1 vssd1 vccd1 vccd1 _15083_/D sky130_fd_sc_hd__mux2_1
XFILLER_42_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10602_ _13718_/Q _10602_/B vssd1 vssd1 vccd1 vccd1 _10602_/X sky130_fd_sc_hd__and2_1
XFILLER_11_932 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14370_ _15287_/CLK _14370_/D vssd1 vssd1 vccd1 vccd1 _14370_/Q sky130_fd_sc_hd__dfxtp_1
X_11582_ _11582_/A _11582_/B vssd1 vssd1 vccd1 vccd1 _11584_/B sky130_fd_sc_hd__xor2_1
XFILLER_80_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_403 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13321_ _13321_/A0 _15651_/Q _13350_/S vssd1 vssd1 vccd1 vccd1 _15651_/D sky130_fd_sc_hd__mux2_1
X_10533_ _11600_/A _13236_/B _10469_/B vssd1 vssd1 vccd1 vccd1 _10533_/X sky130_fd_sc_hd__a21o_1
XFILLER_10_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_745 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13252_ _13252_/A _13252_/B vssd1 vssd1 vccd1 vccd1 _13252_/Y sky130_fd_sc_hd__nor2_1
X_10464_ _07206_/X _10360_/B _10463_/X vssd1 vssd1 vccd1 vccd1 _11598_/A sky130_fd_sc_hd__a21o_4
XFILLER_143_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12203_ _12186_/X _12187_/X _12490_/A vssd1 vssd1 vccd1 vccd1 _12203_/X sky130_fd_sc_hd__mux2_1
XFILLER_108_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13183_ _13229_/A _13183_/B vssd1 vssd1 vccd1 vccd1 _13183_/Y sky130_fd_sc_hd__nor2_1
XFILLER_170_439 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10395_ _10395_/A _10395_/B vssd1 vssd1 vccd1 vccd1 _10399_/A sky130_fd_sc_hd__nand2_1
XFILLER_2_630 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12134_ _12117_/X _12118_/X _12490_/A vssd1 vssd1 vccd1 vccd1 _12134_/X sky130_fd_sc_hd__mux2_1
XFILLER_124_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12065_ _12048_/X _12049_/X _12582_/A vssd1 vssd1 vccd1 vccd1 _12065_/X sky130_fd_sc_hd__mux2_1
XFILLER_42_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11016_ _11010_/Y _11015_/X _11362_/B vssd1 vssd1 vccd1 vccd1 _11016_/X sky130_fd_sc_hd__mux2_1
XFILLER_49_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12967_ _12967_/A1 _13024_/A2 _12966_/X _13024_/B2 vssd1 vssd1 vccd1 vccd1 _12967_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_3371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_372 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11918_ _13940_/Q _13682_/Q _12614_/S vssd1 vssd1 vccd1 vccd1 _11919_/B sky130_fd_sc_hd__mux2_1
X_14706_ _15622_/CLK _14706_/D vssd1 vssd1 vccd1 vccd1 _14706_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12898_ _15426_/Q _15611_/Q _12932_/S vssd1 vssd1 vccd1 vccd1 _15426_/D sky130_fd_sc_hd__mux2_1
XTAP_2681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14637_ _15422_/CLK _14637_/D vssd1 vssd1 vccd1 vccd1 _14637_/Q sky130_fd_sc_hd__dfxtp_1
X_11849_ _15271_/Q _13349_/A0 _11849_/S vssd1 vssd1 vccd1 vccd1 _15271_/D sky130_fd_sc_hd__mux2_1
XFILLER_21_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14568_ _15291_/CLK _14568_/D vssd1 vssd1 vccd1 vccd1 _14568_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_147_915 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13519_ _15378_/CLK _13519_/D vssd1 vssd1 vccd1 vccd1 _13519_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_173_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14499_ _15379_/CLK _14499_/D vssd1 vssd1 vccd1 vccd1 _14499_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_173_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07040_ _07039_/X _13592_/Q _12728_/S vssd1 vssd1 vccd1 vccd1 _07040_/X sky130_fd_sc_hd__mux2_1
XFILLER_174_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08991_ _08975_/X _08978_/X _08985_/X _08990_/X vssd1 vssd1 vccd1 vccd1 _08991_/X
+ sky130_fd_sc_hd__o22a_2
XFILLER_141_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07942_ _14743_/Q _07964_/A _07941_/X _07949_/C1 vssd1 vssd1 vccd1 vccd1 _13550_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_69_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07873_ _13533_/Q _07884_/C vssd1 vssd1 vccd1 vccd1 _07874_/B sky130_fd_sc_hd__xnor2_1
XFILLER_95_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09612_ _13986_/Q _13082_/B2 _09627_/S vssd1 vssd1 vccd1 vccd1 _13986_/D sky130_fd_sc_hd__mux2_1
X_06824_ _14730_/Q _14732_/Q vssd1 vssd1 vccd1 vccd1 _08085_/S sky130_fd_sc_hd__nand2_4
XFILLER_55_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09543_ _09543_/A _09543_/B vssd1 vssd1 vccd1 vccd1 _09543_/X sky130_fd_sc_hd__or2_1
XFILLER_55_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06755_ _13446_/Q vssd1 vssd1 vccd1 vccd1 _06755_/Y sky130_fd_sc_hd__inv_2
XFILLER_52_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09474_ _15301_/Q _15269_/Q _15237_/Q _15168_/Q _09551_/S _09550_/A1 vssd1 vssd1
+ vccd1 vccd1 _09474_/X sky130_fd_sc_hd__mux4_1
X_06686_ _14517_/Q vssd1 vssd1 vccd1 vccd1 _06872_/A sky130_fd_sc_hd__inv_2
XFILLER_169_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08425_ _14586_/Q _14614_/Q _08469_/A vssd1 vssd1 vccd1 vccd1 _08425_/X sky130_fd_sc_hd__and3_4
XFILLER_24_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08356_ _08336_/Y _08355_/Y _11318_/S vssd1 vssd1 vccd1 vccd1 _08357_/A sky130_fd_sc_hd__mux2_1
XFILLER_177_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07307_ _15314_/Q _15470_/Q _07340_/S vssd1 vssd1 vccd1 vccd1 _07307_/X sky130_fd_sc_hd__mux2_8
XFILLER_50_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08287_ _11356_/C _13171_/B vssd1 vssd1 vccd1 vccd1 _11044_/A sky130_fd_sc_hd__and2_1
XFILLER_166_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_918 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07238_ _15328_/Q _15484_/Q _07335_/S vssd1 vssd1 vccd1 vccd1 _07238_/X sky130_fd_sc_hd__mux2_8
XFILLER_146_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07169_ _15343_/Q _15050_/Q _07193_/S vssd1 vssd1 vccd1 vccd1 _07169_/X sky130_fd_sc_hd__mux2_8
XFILLER_3_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10180_ _13080_/B2 _14564_/Q _10192_/S vssd1 vssd1 vccd1 vccd1 _14564_/D sky130_fd_sc_hd__mux2_1
XFILLER_132_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout230 _07736_/A vssd1 vssd1 vccd1 vccd1 _07713_/A sky130_fd_sc_hd__buf_8
XFILLER_121_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout241 _10165_/X vssd1 vssd1 vccd1 vccd1 _10192_/S sky130_fd_sc_hd__buf_12
Xfanout252 _08518_/Y vssd1 vssd1 vccd1 vccd1 _08684_/A2 sky130_fd_sc_hd__clkbuf_16
Xfanout263 _13104_/A2 vssd1 vssd1 vccd1 vccd1 _13118_/A2 sky130_fd_sc_hd__buf_8
Xfanout274 _08503_/Y vssd1 vssd1 vccd1 vccd1 _08690_/A2 sky130_fd_sc_hd__buf_6
XFILLER_87_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout285 _07496_/X vssd1 vssd1 vccd1 vccd1 _13349_/A0 sky130_fd_sc_hd__buf_6
XFILLER_101_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout296 _07476_/X vssd1 vssd1 vccd1 vccd1 _13344_/A0 sky130_fd_sc_hd__buf_8
XFILLER_101_583 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13870_ _15300_/CLK _13870_/D vssd1 vssd1 vccd1 vccd1 _13870_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_46_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12821_ _12828_/A _12821_/B vssd1 vssd1 vccd1 vccd1 _12821_/X sky130_fd_sc_hd__or2_1
XFILLER_34_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12752_ _12743_/A _12750_/X _12751_/X _12788_/C1 vssd1 vssd1 vccd1 vccd1 _15355_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_1210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15540_ _15540_/CLK _15540_/D vssd1 vssd1 vccd1 vccd1 _15540_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_854 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11703_ _13345_/A0 _15134_/Q _11703_/S vssd1 vssd1 vccd1 vccd1 _15134_/D sky130_fd_sc_hd__mux2_1
XTAP_1254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15471_ _15507_/CLK _15471_/D vssd1 vssd1 vccd1 vccd1 _15471_/Q sky130_fd_sc_hd__dfxtp_1
X_12683_ _13590_/Q _12682_/X _12785_/B vssd1 vssd1 vccd1 vccd1 _12683_/X sky130_fd_sc_hd__mux2_1
XTAP_1265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14422_ _15273_/CLK _14422_/D vssd1 vssd1 vccd1 vccd1 _14422_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11634_ _11625_/Y _11629_/B _11627_/B vssd1 vssd1 vccd1 vccd1 _11635_/B sky130_fd_sc_hd__o21ai_2
XFILLER_156_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_740 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14353_ _15526_/CLK _14353_/D vssd1 vssd1 vccd1 vccd1 _14353_/Q sky130_fd_sc_hd__dfxtp_1
X_11565_ _11542_/A _11548_/Y _11556_/A _11554_/X vssd1 vssd1 vccd1 vccd1 _11567_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_128_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13304_ _15636_/Q _12755_/X _13316_/S vssd1 vssd1 vccd1 vccd1 _15636_/D sky130_fd_sc_hd__mux2_1
X_10516_ _07248_/A _10523_/A2 _10515_/X vssd1 vssd1 vccd1 vccd1 _11521_/A sky130_fd_sc_hd__a21o_4
X_14284_ _15518_/CLK _14284_/D vssd1 vssd1 vccd1 vccd1 _14284_/Q sky130_fd_sc_hd__dfxtp_1
X_11496_ _11496_/A _11496_/B _11496_/C vssd1 vssd1 vccd1 vccd1 _11537_/A sky130_fd_sc_hd__and3_2
XFILLER_6_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13235_ _15578_/Q _13219_/S _13234_/X vssd1 vssd1 vccd1 vccd1 _15578_/D sky130_fd_sc_hd__o21a_1
XFILLER_40_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10447_ _07211_/X _10523_/A2 _10446_/X vssd1 vssd1 vccd1 vccd1 _13236_/B sky130_fd_sc_hd__a21o_4
XFILLER_124_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13166_ _13217_/A _13165_/B _13219_/S _11371_/A vssd1 vssd1 vccd1 vccd1 _13166_/X
+ sky130_fd_sc_hd__o211a_1
X_10378_ _11457_/A _11475_/B vssd1 vssd1 vccd1 vccd1 _10381_/A sky130_fd_sc_hd__nand2_1
XFILLER_151_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12117_ _14528_/Q _14141_/Q _14173_/Q _14109_/Q _12472_/S _12465_/S1 vssd1 vssd1
+ vccd1 vccd1 _12117_/X sky130_fd_sc_hd__mux4_1
XFILLER_123_174 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13097_ _15516_/Q _10877_/S _13042_/A _13096_/X vssd1 vssd1 vccd1 vccd1 _15516_/D
+ sky130_fd_sc_hd__a22o_1
X_12048_ _14525_/Q _14138_/Q _14170_/Q _14106_/Q _12246_/S _12268_/A vssd1 vssd1 vccd1
+ vccd1 _12048_/X sky130_fd_sc_hd__mux4_1
XFILLER_66_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13999_ _15677_/CLK _13999_/D vssd1 vssd1 vccd1 vccd1 _13999_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_46_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15669_ _15669_/CLK _15669_/D vssd1 vssd1 vccd1 vccd1 _15669_/Q sky130_fd_sc_hd__dfxtp_1
X_08210_ _13701_/Q _11872_/A1 _08221_/S vssd1 vssd1 vccd1 vccd1 _13701_/D sky130_fd_sc_hd__mux2_1
XFILLER_21_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09190_ _13953_/Q _13695_/Q _09190_/S vssd1 vssd1 vccd1 vccd1 _09190_/X sky130_fd_sc_hd__mux2_1
XFILLER_60_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08141_ input5/X input14/X _08150_/S vssd1 vssd1 vccd1 vccd1 _08141_/X sky130_fd_sc_hd__mux2_1
XFILLER_14_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08072_ _14765_/Q _13643_/Q _08072_/S vssd1 vssd1 vccd1 vccd1 _13643_/D sky130_fd_sc_hd__mux2_1
XFILLER_140_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07023_ _07022_/X _14740_/Q _07098_/S vssd1 vssd1 vccd1 vccd1 _13586_/D sky130_fd_sc_hd__mux2_1
XFILLER_161_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08974_ _09221_/A _08974_/B vssd1 vssd1 vccd1 vccd1 _08974_/X sky130_fd_sc_hd__or2_1
XFILLER_103_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07925_ _13545_/Q _13544_/Q _07924_/D _13546_/Q vssd1 vssd1 vccd1 vccd1 _07925_/Y
+ sky130_fd_sc_hd__a31oi_1
XFILLER_29_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07856_ _07874_/A _07855_/X input35/X vssd1 vssd1 vccd1 vccd1 _07856_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_57_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06807_ _14587_/Q _08392_/B vssd1 vssd1 vccd1 vccd1 _08390_/A sky130_fd_sc_hd__and2_2
XFILLER_16_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07787_ _07787_/A _14730_/Q _12640_/S _07787_/D vssd1 vssd1 vccd1 vccd1 _07802_/C
+ sky130_fd_sc_hd__and4_2
XFILLER_25_810 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09526_ _15679_/Q _13413_/Q _09535_/S vssd1 vssd1 vccd1 vccd1 _09526_/X sky130_fd_sc_hd__mux2_1
XFILLER_37_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06738_ _14493_/Q vssd1 vssd1 vccd1 vccd1 _06738_/Y sky130_fd_sc_hd__inv_2
XPHY_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09457_ _14030_/Q _13998_/Q _09469_/S vssd1 vssd1 vccd1 vccd1 _09457_/X sky130_fd_sc_hd__mux2_1
XPHY_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06669_ _12567_/A vssd1 vssd1 vccd1 vccd1 _06669_/Y sky130_fd_sc_hd__inv_6
XPHY_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08408_ _08756_/B _08777_/A _08407_/Y _13129_/A _13737_/Q vssd1 vssd1 vccd1 vccd1
+ _13737_/D sky130_fd_sc_hd__a32o_1
X_09388_ _09372_/X _09375_/X _09382_/X _09387_/X vssd1 vssd1 vccd1 vccd1 _09388_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_138_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08339_ _11347_/A _08338_/X _08320_/Y _08292_/B vssd1 vssd1 vccd1 vccd1 _08339_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_177_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11350_ _11362_/C _13251_/B _11349_/X _11307_/A vssd1 vssd1 vccd1 vccd1 _11350_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_126_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10301_ _14686_/Q _14871_/Q _10710_/S vssd1 vssd1 vccd1 vccd1 _14686_/D sky130_fd_sc_hd__mux2_1
XFILLER_153_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_992 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11281_ _11330_/A _11265_/X _11280_/Y vssd1 vssd1 vccd1 vccd1 _11281_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_118_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13020_ _10704_/X _14887_/Q _13029_/S vssd1 vssd1 vccd1 vccd1 _13020_/X sky130_fd_sc_hd__mux2_4
X_10232_ _14617_/Q _14770_/Q _10615_/S vssd1 vssd1 vccd1 vccd1 _14617_/D sky130_fd_sc_hd__mux2_1
XFILLER_105_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10163_ _14548_/Q _13349_/A0 _10164_/S vssd1 vssd1 vccd1 vccd1 _14548_/D sky130_fd_sc_hd__mux2_1
XFILLER_133_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14971_ _14988_/CLK _14971_/D vssd1 vssd1 vccd1 vccd1 _14971_/Q sky130_fd_sc_hd__dfxtp_1
X_10094_ _14450_/Q _13347_/A0 _10097_/S vssd1 vssd1 vccd1 vccd1 _14450_/D sky130_fd_sc_hd__mux2_1
XFILLER_59_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13922_ _15664_/CLK _13922_/D vssd1 vssd1 vccd1 vccd1 _13922_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13853_ _14468_/CLK _13853_/D vssd1 vssd1 vccd1 vccd1 _13853_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_28_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12804_ _15363_/Q _12810_/C vssd1 vssd1 vccd1 vccd1 _12805_/B sky130_fd_sc_hd__xor2_1
XFILLER_15_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13784_ _14510_/CLK _13784_/D vssd1 vssd1 vccd1 vccd1 _13784_/Q sky130_fd_sc_hd__dfxtp_4
X_10996_ _11088_/S _10996_/B vssd1 vssd1 vccd1 vccd1 _10996_/Y sky130_fd_sc_hd__nor2_1
XFILLER_37_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15523_ _15523_/CLK _15523_/D vssd1 vssd1 vccd1 vccd1 _15523_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_187_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12735_ _13597_/Q _12734_/X _12785_/B vssd1 vssd1 vccd1 vccd1 _12735_/X sky130_fd_sc_hd__mux2_1
XTAP_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_1034 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15454_ _15606_/CLK _15454_/D vssd1 vssd1 vccd1 vccd1 _15454_/Q sky130_fd_sc_hd__dfxtp_1
X_12666_ _15344_/Q _12666_/B vssd1 vssd1 vccd1 vccd1 _12667_/B sky130_fd_sc_hd__nor2_1
XTAP_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11617_ _11618_/B vssd1 vssd1 vccd1 vccd1 _11617_/Y sky130_fd_sc_hd__inv_2
X_14405_ _14405_/CLK _14405_/D vssd1 vssd1 vccd1 vccd1 _14405_/Q sky130_fd_sc_hd__dfxtp_1
X_15385_ _15385_/CLK _15385_/D vssd1 vssd1 vccd1 vccd1 _15385_/Q sky130_fd_sc_hd__dfxtp_1
X_12597_ _15336_/Q _13139_/S _12596_/X vssd1 vssd1 vccd1 vccd1 _15336_/D sky130_fd_sc_hd__a21o_1
X_11548_ _11576_/A _11549_/B vssd1 vssd1 vccd1 vccd1 _11548_/Y sky130_fd_sc_hd__nand2b_1
X_14336_ _15285_/CLK _14336_/D vssd1 vssd1 vccd1 vccd1 _14336_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_156_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14267_ _15660_/CLK _14267_/D vssd1 vssd1 vccd1 vccd1 _14267_/Q sky130_fd_sc_hd__dfxtp_1
X_11479_ _13199_/B _11480_/B vssd1 vssd1 vccd1 vccd1 _11502_/A sky130_fd_sc_hd__nor2_2
XFILLER_143_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13218_ _13218_/A _13218_/B vssd1 vssd1 vccd1 vccd1 _13218_/Y sky130_fd_sc_hd__nor2_1
X_14198_ _15651_/CLK _14198_/D vssd1 vssd1 vccd1 vccd1 _14198_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13149_ _14609_/Q _15547_/Q _13149_/S vssd1 vssd1 vccd1 vccd1 _15547_/D sky130_fd_sc_hd__mux2_1
XFILLER_32_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07710_ _07708_/Y _07712_/B _07713_/A vssd1 vssd1 vccd1 vccd1 _07710_/Y sky130_fd_sc_hd__o21ai_1
X_08690_ _15376_/Q _08690_/A2 _08690_/B1 _13421_/Q vssd1 vssd1 vccd1 vccd1 _08690_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_66_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07641_ _07638_/Y _07647_/C _07651_/A vssd1 vssd1 vccd1 vccd1 _07641_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_38_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07572_ _13452_/Q _07576_/C _07576_/D vssd1 vssd1 vccd1 vccd1 _07575_/B sky130_fd_sc_hd__and3_1
XFILLER_18_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09311_ _13959_/Q _13701_/Q _09481_/S vssd1 vssd1 vccd1 vccd1 _09311_/X sky130_fd_sc_hd__mux2_1
XFILLER_15_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_179_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09242_ _08507_/A _09239_/X _09241_/X _09524_/A vssd1 vssd1 vccd1 vccd1 _09242_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_22_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09173_ _14531_/Q _14144_/Q _14176_/Q _14112_/Q _09444_/S _09446_/A1 vssd1 vssd1
+ vccd1 vccd1 _09173_/X sky130_fd_sc_hd__mux4_1
XFILLER_159_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08124_ _13657_/Q _10285_/S _08119_/X _08123_/X vssd1 vssd1 vccd1 vccd1 _13657_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_119_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_1052 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08055_ _14748_/Q _13626_/Q _08066_/S vssd1 vssd1 vccd1 vccd1 _13626_/D sky130_fd_sc_hd__mux2_1
X_07006_ _07005_/X _14734_/Q _07098_/S vssd1 vssd1 vccd1 vccd1 _13580_/D sky130_fd_sc_hd__mux2_1
Xoutput39 _07175_/X vssd1 vssd1 vccd1 vccd1 ext_address[13] sky130_fd_sc_hd__clkbuf_2
XFILLER_162_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08957_ _14425_/Q _13130_/B1 _08520_/B _08956_/X vssd1 vssd1 vccd1 vccd1 _08957_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_29_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07908_ _07910_/B _07906_/X _08022_/B vssd1 vssd1 vccd1 vccd1 _07908_/X sky130_fd_sc_hd__a21bo_1
XTAP_3904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08888_ _15273_/Q _15241_/Q _15209_/Q _15140_/Q _09225_/S0 _09225_/S1 vssd1 vssd1
+ vccd1 vccd1 _08888_/X sky130_fd_sc_hd__mux4_1
XFILLER_116_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07839_ _14748_/Q _07830_/A _07838_/Y _12788_/C1 vssd1 vssd1 vccd1 vccd1 _13523_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_3948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_1023 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10850_ _14882_/Q _13786_/Q _12929_/S vssd1 vssd1 vccd1 vccd1 _14882_/D sky130_fd_sc_hd__mux2_1
XFILLER_72_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09509_ _08494_/B _09507_/X _09508_/X vssd1 vssd1 vccd1 vccd1 _09510_/C sky130_fd_sc_hd__a21o_1
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10781_ _14813_/Q _15445_/Q _12917_/S vssd1 vssd1 vccd1 vccd1 _14813_/D sky130_fd_sc_hd__mux2_1
XFILLER_188_13 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12520_ _14030_/Q _13998_/Q _12522_/S vssd1 vssd1 vccd1 vccd1 _12521_/B sky130_fd_sc_hd__mux2_1
XPHY_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12451_ _14027_/Q _13995_/Q _12453_/S vssd1 vssd1 vccd1 vccd1 _12452_/B sky130_fd_sc_hd__mux2_1
XFILLER_166_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11402_ _11382_/Y _11401_/B _11401_/C vssd1 vssd1 vccd1 vccd1 _11402_/Y sky130_fd_sc_hd__a21boi_2
XFILLER_172_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_166_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15170_ _15303_/CLK _15170_/D vssd1 vssd1 vccd1 vccd1 _15170_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_123_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12382_ _14024_/Q _13992_/Q _12518_/S vssd1 vssd1 vccd1 vccd1 _12383_/B sky130_fd_sc_hd__mux2_1
XANTENNA_90 _07265_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_181_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14121_ _15679_/CLK _14121_/D vssd1 vssd1 vccd1 vccd1 _14121_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11333_ _11047_/Y _11307_/B _11332_/X _11344_/A vssd1 vssd1 vccd1 vccd1 _11333_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_125_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14052_ _15651_/CLK _14052_/D vssd1 vssd1 vccd1 vccd1 _14052_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_153_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11264_ _15029_/Q _11302_/A _11262_/Y _11263_/X vssd1 vssd1 vccd1 vccd1 _15029_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_97_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13003_ _07452_/X _13039_/A2 _13002_/X _12944_/A vssd1 vssd1 vccd1 vccd1 _13003_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_180_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10215_ input9/X _08453_/A _13300_/S vssd1 vssd1 vccd1 vccd1 _14600_/D sky130_fd_sc_hd__mux2_1
X_11195_ _11199_/A _11195_/B vssd1 vssd1 vccd1 vccd1 _11195_/Y sky130_fd_sc_hd__nor2_1
X_10146_ _14531_/Q _13332_/A0 _10159_/S vssd1 vssd1 vccd1 vccd1 _14531_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14954_ _14988_/CLK _14954_/D vssd1 vssd1 vccd1 vccd1 _14954_/Q sky130_fd_sc_hd__dfxtp_1
X_10077_ _14433_/Q _13330_/A0 _10092_/S vssd1 vssd1 vccd1 vccd1 _14433_/D sky130_fd_sc_hd__mux2_1
XFILLER_47_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13905_ _14420_/CLK _13905_/D vssd1 vssd1 vccd1 vccd1 _13905_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14885_ _15438_/CLK _14885_/D vssd1 vssd1 vccd1 vccd1 _14885_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_195_clk clkbuf_5_20_0_clk/X vssd1 vssd1 vccd1 vccd1 _15668_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_47_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13836_ _15286_/CLK _13836_/D vssd1 vssd1 vccd1 vccd1 _13836_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10979_ _11259_/S _10979_/B vssd1 vssd1 vccd1 vccd1 _10979_/X sky130_fd_sc_hd__or2_1
X_13767_ _15588_/CLK _13767_/D vssd1 vssd1 vccd1 vccd1 _13767_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15506_ _15519_/CLK _15506_/D vssd1 vssd1 vccd1 vccd1 _15506_/Q sky130_fd_sc_hd__dfxtp_1
X_12718_ _15058_/Q _12717_/X _12792_/B vssd1 vssd1 vccd1 vccd1 _12718_/X sky130_fd_sc_hd__mux2_1
XFILLER_176_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13698_ _14373_/CLK _13698_/D vssd1 vssd1 vccd1 vccd1 _13698_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_188_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15437_ _15623_/CLK _15437_/D vssd1 vssd1 vccd1 vccd1 _15437_/Q sky130_fd_sc_hd__dfxtp_1
X_12649_ _12743_/A _12649_/B vssd1 vssd1 vccd1 vccd1 _12649_/X sky130_fd_sc_hd__or2_1
XFILLER_175_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15368_ _15543_/CLK _15368_/D vssd1 vssd1 vccd1 vccd1 _15368_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14319_ _15199_/CLK _14319_/D vssd1 vssd1 vccd1 vccd1 _14319_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_171_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15299_ _15332_/CLK _15299_/D vssd1 vssd1 vccd1 vccd1 _15299_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_770 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09860_ _14224_/Q _11847_/A1 _09863_/S vssd1 vssd1 vccd1 vccd1 _14224_/D sky130_fd_sc_hd__mux2_1
XTAP_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08811_ _13345_/A0 _13837_/Q _08811_/S vssd1 vssd1 vccd1 vccd1 _13837_/D sky130_fd_sc_hd__mux2_1
X_09791_ _14158_/Q _13346_/A0 _09795_/S vssd1 vssd1 vccd1 vccd1 _14158_/D sky130_fd_sc_hd__mux2_1
XTAP_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08742_ _13446_/Q _08746_/A2 _08750_/A2 _13510_/Q vssd1 vssd1 vccd1 vccd1 _08742_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_38_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08673_ _14497_/Q _08537_/Y _08538_/Y _15379_/Q _08672_/X vssd1 vssd1 vccd1 vccd1
+ _08673_/X sky130_fd_sc_hd__a221o_1
Xclkbuf_leaf_186_clk clkbuf_5_21_0_clk/X vssd1 vssd1 vccd1 vccd1 _15291_/CLK sky130_fd_sc_hd__clkbuf_16
X_07624_ _13468_/Q _07625_/B vssd1 vssd1 vccd1 vccd1 _07624_/Y sky130_fd_sc_hd__nor2_1
XFILLER_54_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07555_ _13450_/Q _13449_/Q _07559_/D vssd1 vssd1 vccd1 vccd1 _07560_/B sky130_fd_sc_hd__and3_1
XFILLER_22_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07486_ _14673_/Q _07490_/B _07498_/C vssd1 vssd1 vccd1 vccd1 _07486_/X sky130_fd_sc_hd__and3_1
X_09225_ _14244_/Q _14276_/Q _14308_/Q _14340_/Q _09225_/S0 _09225_/S1 vssd1 vssd1
+ vccd1 vccd1 _09225_/X sky130_fd_sc_hd__mux4_1
XFILLER_158_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09156_ _09405_/A _09149_/X _09152_/X _09450_/B1 vssd1 vssd1 vccd1 vccd1 _09156_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_147_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_175_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08107_ input13/X input21/X _08133_/S vssd1 vssd1 vccd1 vccd1 _08163_/B sky130_fd_sc_hd__mux2_1
XFILLER_107_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09087_ _14076_/Q _09231_/A2 _09403_/B1 _14044_/Q _09221_/A vssd1 vssd1 vccd1 vccd1
+ _09087_/X sky130_fd_sc_hd__a221o_1
Xclkbuf_leaf_110_clk clkbuf_5_26_0_clk/X vssd1 vssd1 vccd1 vccd1 _15635_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_174_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08038_ _14737_/Q _13577_/Q _08038_/S vssd1 vssd1 vccd1 vccd1 _13577_/D sky130_fd_sc_hd__mux2_1
Xclkbuf_5_8_0_clk clkbuf_5_9_0_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_5_8_0_clk/X sky130_fd_sc_hd__clkbuf_8
XFILLER_123_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10000_ _11854_/A1 _14358_/Q _10029_/S vssd1 vssd1 vccd1 vccd1 _14358_/D sky130_fd_sc_hd__mux2_1
XFILLER_131_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09989_ _11876_/A1 _14348_/Q _09991_/S vssd1 vssd1 vccd1 vccd1 _14348_/D sky130_fd_sc_hd__mux2_1
XFILLER_67_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_1099 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11951_ _12595_/A1 _11950_/X _11949_/X _12618_/C1 vssd1 vssd1 vccd1 vccd1 _11952_/C
+ sky130_fd_sc_hd__a211o_1
Xclkbuf_leaf_177_clk clkbuf_5_23_0_clk/X vssd1 vssd1 vccd1 vccd1 _15680_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_3745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10902_ _11414_/A _10951_/B vssd1 vssd1 vccd1 vccd1 _10902_/Y sky130_fd_sc_hd__nand2_1
XTAP_3778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14670_ _15606_/CLK _14670_/D vssd1 vssd1 vccd1 vccd1 _14670_/Q sky130_fd_sc_hd__dfxtp_1
X_11882_ _15303_/Q _13349_/A0 _11883_/S vssd1 vssd1 vccd1 vccd1 _15303_/D sky130_fd_sc_hd__mux2_1
XTAP_3789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13621_ _15378_/CLK _13621_/D vssd1 vssd1 vccd1 vccd1 _13621_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10833_ _14865_/Q _13803_/Q _12906_/S vssd1 vssd1 vccd1 vccd1 _14865_/D sky130_fd_sc_hd__mux2_1
XFILLER_60_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13552_ _14495_/CLK _13552_/D vssd1 vssd1 vccd1 vccd1 _13552_/Q sky130_fd_sc_hd__dfxtp_1
X_10764_ _15428_/Q _14796_/Q _10764_/S vssd1 vssd1 vccd1 vccd1 _14796_/D sky130_fd_sc_hd__mux2_1
XFILLER_160_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12503_ _12503_/A1 _12502_/X _12501_/X _12503_/C1 vssd1 vssd1 vccd1 vccd1 _12504_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_186_968 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13483_ _15397_/CLK _13483_/D vssd1 vssd1 vccd1 vccd1 _13483_/Q sky130_fd_sc_hd__dfxtp_2
X_10695_ _14757_/Q _10694_/X _10695_/S vssd1 vssd1 vccd1 vccd1 _14757_/D sky130_fd_sc_hd__mux2_1
XFILLER_9_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_0_1_clk clkbuf_1_0_1_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_2_1_0_clk/A sky130_fd_sc_hd__clkbuf_8
XFILLER_9_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12434_ _12618_/A1 _12433_/X _12432_/X _12618_/C1 vssd1 vssd1 vccd1 vccd1 _12435_/C
+ sky130_fd_sc_hd__a211o_1
X_15222_ _15286_/CLK _15222_/D vssd1 vssd1 vccd1 vccd1 _15222_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_166_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12365_ _12595_/A1 _12364_/X _12363_/X _12618_/C1 vssd1 vssd1 vccd1 vccd1 _12366_/C
+ sky130_fd_sc_hd__a211o_1
X_15153_ _15286_/CLK _15153_/D vssd1 vssd1 vccd1 vccd1 _15153_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_101_clk _15447_/CLK vssd1 vssd1 vccd1 vccd1 _15638_/CLK sky130_fd_sc_hd__clkbuf_16
X_11316_ _15036_/Q _11302_/A _08331_/X _11303_/A _11315_/X vssd1 vssd1 vccd1 vccd1
+ _15036_/D sky130_fd_sc_hd__o221a_1
X_14104_ _15081_/CLK _14104_/D vssd1 vssd1 vccd1 vccd1 _14104_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15084_ _15244_/CLK _15084_/D vssd1 vssd1 vccd1 vccd1 _15084_/Q sky130_fd_sc_hd__dfxtp_1
X_12296_ _12595_/A1 _12295_/X _12294_/X _12618_/C1 vssd1 vssd1 vccd1 vccd1 _12297_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_126_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14035_ _14470_/CLK _14035_/D vssd1 vssd1 vccd1 vccd1 _14035_/Q sky130_fd_sc_hd__dfxtp_1
X_11247_ _11380_/A _10895_/B _11437_/A _08232_/A vssd1 vssd1 vccd1 vccd1 _11247_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_141_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11178_ _14981_/Q _11202_/A _11170_/X _11177_/Y vssd1 vssd1 vccd1 vccd1 _14981_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_121_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10129_ _14515_/Q _14763_/Q _10131_/S vssd1 vssd1 vccd1 vccd1 _14515_/D sky130_fd_sc_hd__mux2_1
XFILLER_110_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14937_ _15553_/CLK _14937_/D vssd1 vssd1 vccd1 vccd1 _14937_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_168_clk clkbuf_5_22_0_clk/X vssd1 vssd1 vccd1 vccd1 _15670_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_36_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14868_ _14868_/CLK _14868_/D vssd1 vssd1 vccd1 vccd1 _14868_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_169_1095 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_407 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13819_ _15279_/CLK _13819_/D vssd1 vssd1 vccd1 vccd1 _13819_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14799_ _15534_/CLK _14799_/D vssd1 vssd1 vccd1 vccd1 _14799_/Q sky130_fd_sc_hd__dfxtp_1
X_07340_ _15309_/Q _15465_/Q _07340_/S vssd1 vssd1 vccd1 vccd1 _07341_/A sky130_fd_sc_hd__mux2_4
XFILLER_177_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07271_ _07256_/X _07258_/Y _07264_/X vssd1 vssd1 vccd1 vccd1 _07273_/C sky130_fd_sc_hd__o21a_1
X_09010_ _15654_/Q _13388_/Q _09521_/S vssd1 vssd1 vccd1 vccd1 _09010_/X sky130_fd_sc_hd__mux2_1
XFILLER_136_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_692 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_190 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09912_ _13078_/B2 _14273_/Q _09925_/S vssd1 vssd1 vccd1 vccd1 _14273_/D sky130_fd_sc_hd__mux2_1
XFILLER_144_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout604 _12470_/S vssd1 vssd1 vccd1 vccd1 _11993_/S sky130_fd_sc_hd__clkbuf_16
Xfanout615 _12545_/S vssd1 vssd1 vccd1 vccd1 _12591_/S sky130_fd_sc_hd__buf_12
XFILLER_99_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout626 _14598_/Q vssd1 vssd1 vccd1 vccd1 _08405_/A sky130_fd_sc_hd__buf_12
XFILLER_59_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout637 fanout647/X vssd1 vssd1 vccd1 vccd1 _12788_/C1 sky130_fd_sc_hd__buf_6
XTAP_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09843_ _14207_/Q _13330_/A0 _09858_/S vssd1 vssd1 vccd1 vccd1 _14207_/D sky130_fd_sc_hd__mux2_1
XFILLER_58_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09774_ _14141_/Q _13329_/A0 _09790_/S vssd1 vssd1 vccd1 vccd1 _14141_/D sky130_fd_sc_hd__mux2_1
X_06986_ _14586_/Q _08469_/A vssd1 vssd1 vccd1 vccd1 _06988_/A sky130_fd_sc_hd__and2_1
XFILLER_37_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08725_ _13647_/Q _08523_/Y _08747_/B1 _13480_/Q vssd1 vssd1 vccd1 vccd1 _08725_/X
+ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_159_clk clkbuf_5_19_0_clk/X vssd1 vssd1 vccd1 vccd1 _14606_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_54_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08656_ _13426_/Q _08690_/B1 _08693_/A2 _14499_/Q vssd1 vssd1 vccd1 vccd1 _08656_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_2329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07607_ _07607_/A _07607_/B vssd1 vssd1 vccd1 vccd1 _07607_/Y sky130_fd_sc_hd__nand2_1
XFILLER_53_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_1048 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08587_ _13468_/Q _08684_/A2 _08691_/A2 _13603_/Q vssd1 vssd1 vccd1 vccd1 _08587_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_1639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07538_ _12839_/B _07783_/B vssd1 vssd1 vccd1 vccd1 _07614_/A sky130_fd_sc_hd__or2_4
XFILLER_167_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07469_ _13342_/A0 _13406_/Q _07501_/S vssd1 vssd1 vccd1 vccd1 _13406_/D sky130_fd_sc_hd__mux2_1
XFILLER_10_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09208_ _08487_/A _09206_/X _09207_/X vssd1 vssd1 vccd1 vccd1 _09212_/B sky130_fd_sc_hd__a21o_1
X_10480_ _07261_/A _10360_/B _10479_/X vssd1 vssd1 vccd1 vccd1 _11536_/A sky130_fd_sc_hd__a21oi_4
XFILLER_183_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_25 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09139_ _09221_/A _09139_/B vssd1 vssd1 vccd1 vccd1 _09139_/X sky130_fd_sc_hd__or2_1
XFILLER_5_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12150_ _13886_/Q _14401_/Q _12269_/S vssd1 vssd1 vccd1 vccd1 _12150_/X sky130_fd_sc_hd__mux2_1
XFILLER_136_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11101_ _11344_/A _11179_/B _11099_/Y _11100_/X _10984_/Y vssd1 vssd1 vccd1 vccd1
+ _11101_/X sky130_fd_sc_hd__a221o_1
XFILLER_118_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12081_ _13883_/Q _14398_/Q _12269_/S vssd1 vssd1 vccd1 vccd1 _12081_/X sky130_fd_sc_hd__mux2_1
XFILLER_150_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11032_ _11016_/X _11031_/Y _11129_/A vssd1 vssd1 vccd1 vccd1 _11032_/X sky130_fd_sc_hd__mux2_1
XFILLER_104_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_11 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12983_ _15474_/Q _13105_/A2 _13025_/B1 _12982_/X vssd1 vssd1 vccd1 vccd1 _15474_/D
+ sky130_fd_sc_hd__a22o_1
XTAP_3542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14722_ _15552_/CLK _14722_/D vssd1 vssd1 vccd1 vccd1 _14722_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_3564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11934_ _15110_/Q _15078_/Q _15651_/Q _13385_/Q _12407_/S _12406_/A vssd1 vssd1 vccd1
+ vccd1 _11934_/X sky130_fd_sc_hd__mux4_1
XTAP_3575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_72 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14653_ _14774_/CLK _14653_/D vssd1 vssd1 vccd1 vccd1 _14653_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11865_ _15286_/Q _13332_/A0 _11878_/S vssd1 vssd1 vccd1 vccd1 _15286_/D sky130_fd_sc_hd__mux2_1
XTAP_2874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_790 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13604_ _15624_/CLK _13604_/D vssd1 vssd1 vccd1 vccd1 _13604_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_32_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10816_ _14848_/Q _07260_/A _13138_/S vssd1 vssd1 vccd1 vccd1 _14848_/D sky130_fd_sc_hd__mux2_1
X_11796_ _15219_/Q _13329_/A0 _11816_/S vssd1 vssd1 vccd1 vccd1 _15219_/D sky130_fd_sc_hd__mux2_1
X_14584_ _15530_/CLK _14584_/D vssd1 vssd1 vccd1 vccd1 _14584_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_159_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13535_ _14513_/CLK _13535_/D vssd1 vssd1 vccd1 vccd1 _13535_/Q sky130_fd_sc_hd__dfxtp_1
X_10747_ _15411_/Q _14779_/Q _10759_/S vssd1 vssd1 vccd1 vccd1 _14779_/D sky130_fd_sc_hd__mux2_1
XFILLER_40_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13466_ _15389_/CLK _13466_/D vssd1 vssd1 vccd1 vccd1 _13466_/Q sky130_fd_sc_hd__dfxtp_2
X_10678_ _14982_/Q _10718_/A2 _10722_/B1 _14950_/Q _10677_/X vssd1 vssd1 vccd1 vccd1
+ _10678_/X sky130_fd_sc_hd__a221o_2
XFILLER_127_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15205_ _15615_/CLK _15205_/D vssd1 vssd1 vccd1 vccd1 _15205_/Q sky130_fd_sc_hd__dfxtp_1
X_12417_ _15131_/Q _15099_/Q _15672_/Q _13406_/Q _12430_/S _12563_/A vssd1 vssd1 vccd1
+ vccd1 _12417_/X sky130_fd_sc_hd__mux4_1
X_13397_ _15663_/CLK _13397_/D vssd1 vssd1 vccd1 vccd1 _13397_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_142_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15136_ _15259_/CLK _15136_/D vssd1 vssd1 vccd1 vccd1 _15136_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12348_ _15128_/Q _15096_/Q _15669_/Q _13403_/Q _12541_/S _12540_/A vssd1 vssd1 vccd1
+ vccd1 _12348_/X sky130_fd_sc_hd__mux4_1
XFILLER_141_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_492 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15067_ _15067_/CLK _15067_/D vssd1 vssd1 vccd1 vccd1 _15067_/Q sky130_fd_sc_hd__dfxtp_4
X_12279_ _15125_/Q _15093_/Q _15666_/Q _13400_/Q _12612_/S _12383_/A vssd1 vssd1 vccd1
+ vccd1 _12279_/X sky130_fd_sc_hd__mux4_1
XFILLER_4_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14018_ _15661_/CLK _14018_/D vssd1 vssd1 vccd1 vccd1 _14018_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06840_ _08465_/B _06808_/X _06835_/X _06839_/X _15615_/Q vssd1 vssd1 vccd1 vccd1
+ _06840_/X sky130_fd_sc_hd__o2111a_1
XFILLER_67_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06771_ _08151_/S _14900_/Q _06771_/C vssd1 vssd1 vccd1 vccd1 _08185_/A sky130_fd_sc_hd__and3b_4
XFILLER_83_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08510_ _08724_/C _08510_/B _08512_/B vssd1 vssd1 vccd1 vccd1 _08510_/X sky130_fd_sc_hd__and3_4
X_09490_ _15677_/Q _13411_/Q _09551_/S vssd1 vssd1 vccd1 vccd1 _09490_/X sky130_fd_sc_hd__mux2_1
XFILLER_36_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_159 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08441_ _09405_/A _08390_/C _08425_/X vssd1 vssd1 vccd1 vccd1 _08441_/X sky130_fd_sc_hd__a21o_1
XFILLER_23_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08372_ _08244_/A _13760_/Q _15412_/Q _08244_/B vssd1 vssd1 vccd1 vccd1 _08372_/X
+ sky130_fd_sc_hd__a22o_2
XFILLER_51_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07323_ _15310_/Q _15466_/Q _07340_/S vssd1 vssd1 vccd1 vccd1 _07324_/A sky130_fd_sc_hd__mux2_4
XFILLER_177_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07254_ _15323_/Q _15479_/Q _07335_/S vssd1 vssd1 vccd1 vccd1 _10481_/A sky130_fd_sc_hd__mux2_8
XFILLER_104_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07185_ _15359_/Q _15066_/Q _07193_/S vssd1 vssd1 vccd1 vccd1 _07185_/X sky130_fd_sc_hd__mux2_2
XFILLER_145_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_824 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout401 _06825_/X vssd1 vssd1 vccd1 vccd1 _12662_/S sky130_fd_sc_hd__clkbuf_16
Xfanout412 _10983_/X vssd1 vssd1 vccd1 vccd1 _11202_/A sky130_fd_sc_hd__buf_12
XFILLER_99_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout423 _10567_/Y vssd1 vssd1 vccd1 vccd1 _10569_/B sky130_fd_sc_hd__buf_12
Xfanout434 _08225_/Y vssd1 vssd1 vccd1 vccd1 _10457_/A2 sky130_fd_sc_hd__buf_12
Xfanout445 _12763_/S vssd1 vssd1 vccd1 vccd1 _12785_/B sky130_fd_sc_hd__buf_12
XFILLER_86_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout456 _10244_/S vssd1 vssd1 vccd1 vccd1 _10715_/S sky130_fd_sc_hd__buf_12
Xfanout467 _06672_/Y vssd1 vssd1 vccd1 vccd1 _12503_/C1 sky130_fd_sc_hd__buf_12
X_09826_ _14192_/Q _13348_/A0 _09828_/S vssd1 vssd1 vccd1 vccd1 _14192_/D sky130_fd_sc_hd__mux2_1
XFILLER_59_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout478 _12548_/S vssd1 vssd1 vccd1 vccd1 _12536_/A sky130_fd_sc_hd__buf_12
Xfanout489 _15526_/Q vssd1 vssd1 vccd1 vccd1 _07335_/S sky130_fd_sc_hd__buf_12
XFILLER_100_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09757_ _14125_/Q _13345_/A0 _09757_/S vssd1 vssd1 vccd1 vccd1 _14125_/D sky130_fd_sc_hd__mux2_1
X_06969_ _06969_/A _06977_/A _06976_/B _06969_/D vssd1 vssd1 vccd1 vccd1 _06974_/A
+ sky130_fd_sc_hd__or4_1
XFILLER_73_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08708_ _14492_/Q _08748_/B1 _08706_/X _08707_/X vssd1 vssd1 vccd1 vccd1 _08709_/C
+ sky130_fd_sc_hd__a211o_1
XTAP_2126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09688_ _14059_/Q _13343_/A0 _09690_/S vssd1 vssd1 vccd1 vccd1 _14059_/D sky130_fd_sc_hd__mux2_1
XTAP_2137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08639_ _13790_/Q _08638_/X _12917_/S vssd1 vssd1 vccd1 vccd1 _13790_/D sky130_fd_sc_hd__mux2_1
XTAP_1425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11650_ _13325_/A0 _15082_/Q _11675_/S vssd1 vssd1 vccd1 vccd1 _15082_/D sky130_fd_sc_hd__mux2_1
XTAP_1458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10601_ _14999_/Q _10569_/B _10733_/B1 _14935_/Q _10732_/C1 vssd1 vssd1 vccd1 vccd1
+ _10601_/X sky130_fd_sc_hd__a221o_1
XFILLER_168_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11581_ _11589_/B _11589_/C _13236_/A vssd1 vssd1 vccd1 vccd1 _11582_/B sky130_fd_sc_hd__a21o_1
XFILLER_120_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10532_ _10532_/A _10532_/B vssd1 vssd1 vccd1 vccd1 _10532_/Y sky130_fd_sc_hd__nor2_1
X_13320_ _13320_/A0 _15650_/Q _13350_/S vssd1 vssd1 vccd1 vccd1 _15650_/D sky130_fd_sc_hd__mux2_1
XFILLER_155_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10463_ _10520_/A1 _13781_/Q _13749_/Q _10520_/B2 vssd1 vssd1 vccd1 vccd1 _10463_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_108_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13251_ _13251_/A _13251_/B vssd1 vssd1 vccd1 vccd1 _13251_/X sky130_fd_sc_hd__or2_1
XFILLER_129_62 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12202_ _12195_/X _12197_/X _12199_/X _12201_/X _12501_/C1 vssd1 vssd1 vccd1 vccd1
+ _12202_/X sky130_fd_sc_hd__o221a_1
XFILLER_89_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13182_ _15561_/Q _13241_/A2 _13180_/Y _13181_/Y vssd1 vssd1 vccd1 vccd1 _15561_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_159_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10394_ _13177_/A _13178_/B vssd1 vssd1 vccd1 vccd1 _10395_/B sky130_fd_sc_hd__nand2b_1
X_12133_ _12126_/X _12128_/X _12130_/X _12132_/X _12501_/C1 vssd1 vssd1 vccd1 vccd1
+ _12133_/X sky130_fd_sc_hd__o221a_1
XFILLER_89_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12064_ _12057_/X _12059_/X _12061_/X _12063_/X _12455_/C1 vssd1 vssd1 vccd1 vccd1
+ _12064_/X sky130_fd_sc_hd__o221a_1
XFILLER_150_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11015_ _10350_/Y _11357_/B _11079_/B _11349_/A vssd1 vssd1 vccd1 vccd1 _11015_/X
+ sky130_fd_sc_hd__a2bb2o_1
XTAP_4040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12966_ _10614_/X _14869_/Q _13038_/S vssd1 vssd1 vccd1 vccd1 _12966_/X sky130_fd_sc_hd__mux2_2
XTAP_3361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14705_ _15623_/CLK _14705_/D vssd1 vssd1 vccd1 vccd1 _14705_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11917_ _12618_/A1 _11912_/X _11915_/X _11916_/X _08405_/D vssd1 vssd1 vccd1 vccd1
+ _11929_/B sky130_fd_sc_hd__a221o_1
XFILLER_73_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12897_ _15425_/Q _15610_/Q _12933_/S vssd1 vssd1 vccd1 vccd1 _15425_/D sky130_fd_sc_hd__mux2_1
XTAP_2682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14636_ _15641_/CLK _14636_/D vssd1 vssd1 vccd1 vccd1 _14636_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11848_ _15270_/Q _11881_/A1 _11850_/S vssd1 vssd1 vccd1 vccd1 _15270_/D sky130_fd_sc_hd__mux2_1
XFILLER_33_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14567_ _15666_/CLK _14567_/D vssd1 vssd1 vccd1 vccd1 _14567_/Q sky130_fd_sc_hd__dfxtp_1
X_11779_ _15205_/Q _10344_/S _11777_/B _10563_/B vssd1 vssd1 vccd1 vccd1 _15205_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_13_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13518_ _15378_/CLK _13518_/D vssd1 vssd1 vccd1 vccd1 _13518_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_159_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14498_ _15379_/CLK _14498_/D vssd1 vssd1 vccd1 vccd1 _14498_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_158_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13449_ _15399_/CLK _13449_/D vssd1 vssd1 vccd1 vccd1 _13449_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_155_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15119_ _15253_/CLK _15119_/D vssd1 vssd1 vccd1 vccd1 _15119_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_126_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08990_ _09449_/B2 _08986_/X _08989_/X vssd1 vssd1 vccd1 vccd1 _08990_/X sky130_fd_sc_hd__a21o_1
XFILLER_142_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07941_ _07943_/B _07940_/X _07964_/A vssd1 vssd1 vccd1 vccd1 _07941_/X sky130_fd_sc_hd__a21bo_1
XFILLER_142_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07872_ _14757_/Q _07874_/A _07871_/Y _08002_/C1 vssd1 vssd1 vccd1 vccd1 _13532_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_28_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09611_ _13985_/Q _13333_/A0 _09627_/S vssd1 vssd1 vccd1 vccd1 _13985_/D sky130_fd_sc_hd__mux2_1
XFILLER_84_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06823_ _08086_/A _06825_/C vssd1 vssd1 vccd1 vccd1 _08078_/B sky130_fd_sc_hd__nand2_1
XFILLER_23_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09542_ _14387_/Q _15203_/Q _13842_/Q _14581_/Q _09557_/S _13144_/A0 vssd1 vssd1
+ vccd1 vccd1 _09543_/B sky130_fd_sc_hd__mux4_1
X_06754_ _13478_/Q vssd1 vssd1 vccd1 vccd1 _06754_/Y sky130_fd_sc_hd__inv_2
XFILLER_83_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09473_ _12320_/A _09463_/X _09472_/X _09453_/X vssd1 vssd1 vccd1 vccd1 _13934_/D
+ sky130_fd_sc_hd__a31o_1
X_06685_ _14613_/Q vssd1 vssd1 vccd1 vccd1 _06685_/Y sky130_fd_sc_hd__inv_2
XFILLER_51_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_90_clk clkbuf_5_13_0_clk/X vssd1 vssd1 vccd1 vccd1 _14851_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_145_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08424_ _13743_/Q _13120_/S _08423_/X vssd1 vssd1 vccd1 vccd1 _13743_/D sky130_fd_sc_hd__a21o_1
X_08355_ _08355_/A _10991_/A vssd1 vssd1 vccd1 vccd1 _08355_/Y sky130_fd_sc_hd__nor2_1
X_07306_ _07306_/A vssd1 vssd1 vccd1 vccd1 _07306_/Y sky130_fd_sc_hd__inv_2
XFILLER_133_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08286_ _07321_/A _10481_/B _08285_/X vssd1 vssd1 vccd1 vccd1 _13171_/B sky130_fd_sc_hd__a21o_4
XFILLER_109_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07237_ _07237_/A vssd1 vssd1 vccd1 vccd1 _07237_/Y sky130_fd_sc_hd__inv_2
XFILLER_109_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_166_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07168_ _15342_/Q _15049_/Q _07193_/S vssd1 vssd1 vccd1 vccd1 _07168_/X sky130_fd_sc_hd__mux2_8
XFILLER_180_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07099_ _14924_/Q _14923_/Q _14898_/Q _10561_/B vssd1 vssd1 vccd1 vccd1 _07157_/A
+ sky130_fd_sc_hd__and4b_4
XFILLER_182_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout220 _08784_/X vssd1 vssd1 vccd1 vccd1 _08816_/S sky130_fd_sc_hd__buf_12
Xfanout231 _07614_/A vssd1 vssd1 vccd1 vccd1 _07644_/A sky130_fd_sc_hd__buf_8
XFILLER_132_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout242 _10165_/X vssd1 vssd1 vccd1 vccd1 _10197_/S sky130_fd_sc_hd__buf_12
Xfanout253 _08189_/Y vssd1 vssd1 vccd1 vccd1 _08216_/S sky130_fd_sc_hd__buf_12
Xfanout264 _13044_/X vssd1 vssd1 vccd1 vccd1 _13104_/A2 sky130_fd_sc_hd__buf_12
XFILLER_101_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout275 _07157_/A vssd1 vssd1 vccd1 vccd1 _07163_/A sky130_fd_sc_hd__buf_12
Xfanout286 _13348_/A0 vssd1 vssd1 vccd1 vccd1 _11881_/A1 sky130_fd_sc_hd__buf_6
XFILLER_87_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09809_ _14175_/Q _13331_/A0 _09823_/S vssd1 vssd1 vccd1 vccd1 _14175_/D sky130_fd_sc_hd__mux2_1
Xfanout297 _13343_/A0 vssd1 vssd1 vccd1 vccd1 _11876_/A1 sky130_fd_sc_hd__buf_6
XFILLER_59_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12820_ _12827_/B _12820_/B vssd1 vssd1 vccd1 vccd1 _12821_/B sky130_fd_sc_hd__nor2_1
XFILLER_131_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12751_ _15355_/Q _12765_/B vssd1 vssd1 vccd1 vccd1 _12751_/X sky130_fd_sc_hd__or2_1
XTAP_1211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_81_clk clkbuf_5_15_0_clk/X vssd1 vssd1 vccd1 vccd1 _15607_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_1233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11702_ _13344_/A0 _15133_/Q _11703_/S vssd1 vssd1 vccd1 vccd1 _15133_/D sky130_fd_sc_hd__mux2_1
XFILLER_91_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15470_ _15519_/CLK _15470_/D vssd1 vssd1 vccd1 vccd1 _15470_/Q sky130_fd_sc_hd__dfxtp_1
X_12682_ _15053_/Q _12681_/Y _12792_/B vssd1 vssd1 vccd1 vccd1 _12682_/X sky130_fd_sc_hd__mux2_1
XTAP_1266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14421_ _15324_/CLK _14421_/D vssd1 vssd1 vccd1 vccd1 _14421_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11633_ _11633_/A _11633_/B vssd1 vssd1 vccd1 vccd1 _11635_/A sky130_fd_sc_hd__xnor2_2
XFILLER_24_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_752 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14352_ _15200_/CLK _14352_/D vssd1 vssd1 vccd1 vccd1 _14352_/Q sky130_fd_sc_hd__dfxtp_1
X_11564_ _11564_/A _11564_/B vssd1 vssd1 vccd1 vccd1 _11576_/C sky130_fd_sc_hd__nand2_2
XFILLER_10_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13303_ _15635_/Q _12747_/Y _13316_/S vssd1 vssd1 vccd1 vccd1 _15635_/D sky130_fd_sc_hd__mux2_1
XFILLER_156_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10515_ _14582_/Q _13756_/Q _15416_/Q _10515_/B2 vssd1 vssd1 vccd1 vccd1 _10515_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_10_273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11495_ _15058_/Q _11474_/S _11493_/Y _11494_/X vssd1 vssd1 vccd1 vccd1 _15058_/D
+ sky130_fd_sc_hd__a22o_1
X_14283_ _15527_/CLK _14283_/D vssd1 vssd1 vccd1 vccd1 _14283_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_157_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13234_ _11598_/A _13232_/X _13233_/Y _13214_/B vssd1 vssd1 vccd1 vccd1 _13234_/X
+ sky130_fd_sc_hd__a31o_1
X_10446_ _08244_/A _13748_/Q _15424_/Q _08244_/B vssd1 vssd1 vccd1 vccd1 _10446_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_109_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10377_ _07289_/X _10360_/B _10376_/X vssd1 vssd1 vccd1 vccd1 _11475_/B sky130_fd_sc_hd__a21o_4
X_13165_ _13217_/A _13165_/B vssd1 vssd1 vccd1 vccd1 _13165_/Y sky130_fd_sc_hd__nand2_1
XFILLER_97_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12116_ _14464_/Q _14432_/Q _13853_/Q _14206_/Q _08457_/A _12489_/S1 vssd1 vssd1
+ vccd1 vccd1 _12116_/X sky130_fd_sc_hd__mux4_1
XFILLER_151_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13096_ _13011_/X _13118_/A2 _13114_/B1 _07464_/X vssd1 vssd1 vccd1 vccd1 _13096_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_111_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12047_ _14461_/Q _14429_/Q _13850_/Q _14203_/Q _12154_/S _12253_/S1 vssd1 vssd1
+ vccd1 vccd1 _12047_/X sky130_fd_sc_hd__mux4_1
XFILLER_46_1072 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_1075 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_800 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_351 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13998_ _15334_/CLK _13998_/D vssd1 vssd1 vccd1 vccd1 _13998_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12949_ _07380_/X _13039_/A2 _12948_/X _12944_/A vssd1 vssd1 vccd1 vccd1 _12949_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_3191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_72_clk clkbuf_5_14_0_clk/X vssd1 vssd1 vccd1 vccd1 _15596_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_178_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15668_ _15668_/CLK _15668_/D vssd1 vssd1 vccd1 vccd1 _15668_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_2_1_0_clk clkbuf_2_1_0_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_2_1_1_clk/A sky130_fd_sc_hd__clkbuf_8
XFILLER_92_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14619_ _14892_/CLK _14619_/D vssd1 vssd1 vccd1 vccd1 _14619_/Q sky130_fd_sc_hd__dfxtp_1
X_15599_ _15599_/CLK _15599_/D vssd1 vssd1 vccd1 vccd1 _15599_/Q sky130_fd_sc_hd__dfxtp_1
X_08140_ _13661_/Q _10285_/S _08119_/X _08139_/X vssd1 vssd1 vccd1 vccd1 _13661_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_53_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08071_ _14764_/Q _13642_/Q _08072_/S vssd1 vssd1 vccd1 vccd1 _13642_/D sky130_fd_sc_hd__mux2_1
X_07022_ _07021_/X _13586_/Q _12662_/S vssd1 vssd1 vccd1 vccd1 _07022_/X sky130_fd_sc_hd__mux2_1
XFILLER_134_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_248 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08973_ _14360_/Q _15176_/Q _13815_/Q _14554_/Q _09225_/S0 _09225_/S1 vssd1 vssd1
+ vccd1 vccd1 _08974_/B sky130_fd_sc_hd__mux4_1
XFILLER_114_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07924_ _13546_/Q _13545_/Q _13544_/Q _07924_/D vssd1 vssd1 vccd1 vccd1 _07935_/D
+ sky130_fd_sc_hd__and4_2
XFILLER_152_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1058 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07855_ _13528_/Q _07855_/B vssd1 vssd1 vccd1 vccd1 _07855_/X sky130_fd_sc_hd__xor2_1
XFILLER_28_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06806_ _06806_/A _06806_/B _06806_/C vssd1 vssd1 vccd1 vccd1 _06806_/X sky130_fd_sc_hd__and3_1
XFILLER_25_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07786_ _13510_/Q _13509_/Q vssd1 vssd1 vccd1 vccd1 _07787_/D sky130_fd_sc_hd__and2_1
XFILLER_43_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_822 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09525_ _14548_/Q _14161_/Q _14193_/Q _14129_/Q _09535_/S _08494_/B vssd1 vssd1 vccd1
+ vccd1 _09525_/X sky130_fd_sc_hd__mux4_1
X_06737_ _13453_/Q vssd1 vssd1 vccd1 vccd1 _07571_/B sky130_fd_sc_hd__clkinv_2
XFILLER_71_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_63_clk clkbuf_5_11_0_clk/X vssd1 vssd1 vccd1 vccd1 _15054_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_64_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09456_ _09546_/S1 _09454_/X _09455_/X vssd1 vssd1 vccd1 vccd1 _09456_/X sky130_fd_sc_hd__a21o_1
X_06668_ _14588_/Q vssd1 vssd1 vccd1 vccd1 _08392_/A sky130_fd_sc_hd__inv_2
XFILLER_101_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08407_ _14596_/Q _12946_/B vssd1 vssd1 vccd1 vccd1 _08407_/Y sky130_fd_sc_hd__nand2_1
XFILLER_101_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09387_ _08668_/D _09383_/X _09384_/X _09386_/X vssd1 vssd1 vccd1 vccd1 _09387_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_184_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_509 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08338_ _08298_/B _08337_/X _11297_/S vssd1 vssd1 vccd1 vccd1 _08338_/X sky130_fd_sc_hd__mux2_1
XFILLER_165_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08269_ _11356_/C _13162_/B vssd1 vssd1 vccd1 vccd1 _08273_/A sky130_fd_sc_hd__nor2_1
X_10300_ _14685_/Q _14870_/Q _10710_/S vssd1 vssd1 vccd1 vccd1 _14685_/D sky130_fd_sc_hd__mux2_1
XFILLER_137_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11280_ _11330_/A _11280_/B vssd1 vssd1 vccd1 vccd1 _11280_/Y sky130_fd_sc_hd__nor2_1
XFILLER_3_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10231_ _14616_/Q _14769_/Q _10735_/S vssd1 vssd1 vccd1 vccd1 _14616_/D sky130_fd_sc_hd__mux2_1
XFILLER_152_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10162_ _14547_/Q _11881_/A1 _10164_/S vssd1 vssd1 vccd1 vccd1 _14547_/D sky130_fd_sc_hd__mux2_1
XFILLER_106_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_156_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14970_ _14988_/CLK _14970_/D vssd1 vssd1 vccd1 vccd1 _14970_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10093_ _14449_/Q _11879_/A1 _10097_/S vssd1 vssd1 vccd1 vccd1 _14449_/D sky130_fd_sc_hd__mux2_1
XFILLER_102_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13921_ _15497_/CLK _13921_/D vssd1 vssd1 vccd1 vccd1 _13921_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13852_ _15181_/CLK _13852_/D vssd1 vssd1 vccd1 vccd1 _13852_/Q sky130_fd_sc_hd__dfxtp_1
X_12803_ _15362_/Q _12765_/B _12802_/X _12809_/C1 vssd1 vssd1 vccd1 vccd1 _15362_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_28_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13783_ _14510_/CLK _13783_/D vssd1 vssd1 vccd1 vccd1 _13783_/Q sky130_fd_sc_hd__dfxtp_4
X_10995_ _13162_/B _13165_/B _11349_/B vssd1 vssd1 vccd1 vccd1 _10996_/B sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_54_clk clkbuf_5_8_0_clk/X vssd1 vssd1 vccd1 vccd1 _15000_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15522_ _15527_/CLK _15522_/D vssd1 vssd1 vccd1 vccd1 _15522_/Q sky130_fd_sc_hd__dfxtp_1
X_12734_ _15060_/Q _12733_/Y _12792_/B vssd1 vssd1 vccd1 vccd1 _12734_/X sky130_fd_sc_hd__mux2_1
XFILLER_163_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15453_ _15453_/CLK _15453_/D vssd1 vssd1 vccd1 vccd1 _15453_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_679 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12665_ _15344_/Q _12666_/B vssd1 vssd1 vccd1 vccd1 _12679_/C sky130_fd_sc_hd__and2_2
XTAP_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14404_ _14415_/CLK _14404_/D vssd1 vssd1 vccd1 vccd1 _14404_/Q sky130_fd_sc_hd__dfxtp_1
X_11616_ _11616_/A _11616_/B vssd1 vssd1 vccd1 vccd1 _11618_/B sky130_fd_sc_hd__xor2_4
X_15384_ _15385_/CLK _15384_/D vssd1 vssd1 vccd1 vccd1 _15384_/Q sky130_fd_sc_hd__dfxtp_1
X_12596_ _12596_/A _12596_/B _12596_/C vssd1 vssd1 vccd1 vccd1 _12596_/X sky130_fd_sc_hd__and3_1
XFILLER_184_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14335_ _15181_/CLK _14335_/D vssd1 vssd1 vccd1 vccd1 _14335_/Q sky130_fd_sc_hd__dfxtp_1
X_11547_ _11508_/B _11546_/X _11545_/X vssd1 vssd1 vccd1 vccd1 _11549_/B sky130_fd_sc_hd__a21o_2
XFILLER_171_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14266_ _14462_/CLK _14266_/D vssd1 vssd1 vccd1 vccd1 _14266_/Q sky130_fd_sc_hd__dfxtp_1
X_11478_ _11496_/A _11478_/B vssd1 vssd1 vccd1 vccd1 _11480_/B sky130_fd_sc_hd__xor2_2
XFILLER_109_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13217_ _13217_/A _13217_/B vssd1 vssd1 vccd1 vccd1 _13218_/B sky130_fd_sc_hd__xnor2_1
X_10429_ _10429_/A _10429_/B vssd1 vssd1 vccd1 vccd1 _10430_/B sky130_fd_sc_hd__and2_1
X_14197_ _14197_/CLK _14197_/D vssd1 vssd1 vccd1 vccd1 _14197_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_140_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13148_ _14608_/Q _15546_/Q _13154_/S vssd1 vssd1 vccd1 vccd1 _15546_/D sky130_fd_sc_hd__mux2_1
XTAP_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13079_ _15507_/Q _13105_/A2 _13105_/B1 _13078_/X vssd1 vssd1 vccd1 vccd1 _15507_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_111_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07640_ _07655_/A _07655_/B vssd1 vssd1 vccd1 vccd1 _07647_/C sky130_fd_sc_hd__and2_2
XFILLER_54_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07571_ _07571_/A _07571_/B vssd1 vssd1 vccd1 vccd1 _07576_/D sky130_fd_sc_hd__nor2_1
XFILLER_47_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_45_clk clkbuf_5_9_0_clk/X vssd1 vssd1 vccd1 vccd1 _15046_/CLK sky130_fd_sc_hd__clkbuf_16
X_09310_ _08510_/B _09308_/X _09309_/X _08519_/B _13049_/A1 vssd1 vssd1 vccd1 vccd1
+ _09310_/X sky130_fd_sc_hd__a221o_1
XFILLER_179_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09241_ _09543_/A _09241_/B vssd1 vssd1 vccd1 vccd1 _09241_/X sky130_fd_sc_hd__or2_1
XFILLER_61_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09172_ _09405_/A _09172_/B _09172_/C vssd1 vssd1 vccd1 vccd1 _09172_/X sky130_fd_sc_hd__and3_1
XFILLER_178_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08123_ _08093_/B _08120_/X _08121_/X _08122_/Y vssd1 vssd1 vccd1 vccd1 _08123_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_174_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_418 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08054_ _14747_/Q _13625_/Q _08066_/S vssd1 vssd1 vccd1 vccd1 _13625_/D sky130_fd_sc_hd__mux2_1
XFILLER_147_598 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07005_ _14645_/Q _13580_/Q _12640_/S vssd1 vssd1 vccd1 vccd1 _07005_/X sky130_fd_sc_hd__mux2_1
XFILLER_162_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08956_ _13846_/Q _14199_/Q _09230_/S vssd1 vssd1 vccd1 vccd1 _08956_/X sky130_fd_sc_hd__mux2_1
X_07907_ _07907_/A _08074_/B vssd1 vssd1 vccd1 vccd1 _07907_/Y sky130_fd_sc_hd__nand2_4
XFILLER_29_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08887_ _09221_/A _08887_/B vssd1 vssd1 vccd1 vccd1 _08887_/X sky130_fd_sc_hd__or2_1
XFILLER_84_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07838_ _07847_/D _07837_/Y _07830_/A vssd1 vssd1 vccd1 vccd1 _07838_/Y sky130_fd_sc_hd__o21ai_1
XTAP_3938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07769_ _13506_/Q _07769_/B vssd1 vssd1 vccd1 vccd1 _07776_/C sky130_fd_sc_hd__and2_2
Xclkbuf_leaf_36_clk clkbuf_5_12_0_clk/X vssd1 vssd1 vccd1 vccd1 _15588_/CLK sky130_fd_sc_hd__clkbuf_16
X_09508_ _14096_/Q _09522_/A2 _09519_/B1 _14064_/Q _09532_/A vssd1 vssd1 vccd1 vccd1
+ _09508_/X sky130_fd_sc_hd__a221o_1
XFILLER_25_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10780_ _14812_/Q _15444_/Q _12917_/S vssd1 vssd1 vccd1 vccd1 _14812_/D sky130_fd_sc_hd__mux2_1
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09439_ _14254_/Q _14286_/Q _14318_/Q _14350_/Q _09444_/S _09448_/S1 vssd1 vssd1
+ vccd1 vccd1 _09439_/X sky130_fd_sc_hd__mux4_1
XPHY_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12450_ _12477_/A1 _12449_/X _12502_/S vssd1 vssd1 vccd1 vccd1 _12450_/X sky130_fd_sc_hd__a21o_1
XFILLER_36_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11401_ _11401_/A _11401_/B _11401_/C vssd1 vssd1 vccd1 vccd1 _11423_/C sky130_fd_sc_hd__and3_1
XFILLER_138_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12381_ _12615_/A1 _12380_/X _12617_/S vssd1 vssd1 vccd1 vccd1 _12381_/X sky130_fd_sc_hd__a21o_1
XANTENNA_80 _07110_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_91 _13202_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_1085 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14120_ _15161_/CLK _14120_/D vssd1 vssd1 vccd1 vccd1 _14120_/Q sky130_fd_sc_hd__dfxtp_1
X_11332_ _11330_/A _11331_/Y _11330_/Y _08249_/Y vssd1 vssd1 vccd1 vccd1 _11332_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_67_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14051_ _14083_/CLK _14051_/D vssd1 vssd1 vccd1 vccd1 _14051_/Q sky130_fd_sc_hd__dfxtp_1
X_11263_ _11344_/A _08249_/Y _08292_/B _11346_/A2 vssd1 vssd1 vccd1 vccd1 _11263_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_180_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13002_ _10674_/X _14881_/Q _13029_/S vssd1 vssd1 vccd1 vccd1 _13002_/X sky130_fd_sc_hd__mux2_8
XFILLER_4_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10214_ input8/X _12379_/A _13309_/A vssd1 vssd1 vccd1 vccd1 _14599_/D sky130_fd_sc_hd__mux2_1
XFILLER_79_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11194_ _14989_/Q _11164_/S _11170_/X _11193_/Y vssd1 vssd1 vccd1 vccd1 _14989_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_79_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10145_ _14530_/Q _11689_/A0 _10159_/S vssd1 vssd1 vccd1 vccd1 _14530_/D sky130_fd_sc_hd__mux2_1
XFILLER_97_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10076_ _14432_/Q _13329_/A0 _10092_/S vssd1 vssd1 vccd1 vccd1 _14432_/D sky130_fd_sc_hd__mux2_1
X_14953_ _15581_/CLK _14953_/D vssd1 vssd1 vccd1 vccd1 _14953_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13904_ _15226_/CLK _13904_/D vssd1 vssd1 vccd1 vccd1 _13904_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_78_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14884_ _15624_/CLK _14884_/D vssd1 vssd1 vccd1 vccd1 _14884_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13835_ _15652_/CLK _13835_/D vssd1 vssd1 vccd1 vccd1 _13835_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_27_clk clkbuf_5_6_0_clk/X vssd1 vssd1 vccd1 vccd1 _15508_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_16_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xcore_650 vssd1 vssd1 vccd1 vccd1 ext_valid core_650/LO sky130_fd_sc_hd__conb_1
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13766_ _14888_/CLK _13766_/D vssd1 vssd1 vccd1 vccd1 _13766_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_188_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10978_ _11037_/A _13217_/B _11305_/C vssd1 vssd1 vccd1 vccd1 _10978_/X sky130_fd_sc_hd__o21a_1
XFILLER_43_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15505_ _15508_/CLK _15505_/D vssd1 vssd1 vccd1 vccd1 _15505_/Q sky130_fd_sc_hd__dfxtp_1
X_12717_ _15351_/Q _12723_/C vssd1 vssd1 vccd1 vccd1 _12717_/X sky130_fd_sc_hd__xor2_1
X_13697_ _15657_/CLK _13697_/D vssd1 vssd1 vccd1 vccd1 _13697_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15436_ _15622_/CLK _15436_/D vssd1 vssd1 vccd1 vccd1 _15436_/Q sky130_fd_sc_hd__dfxtp_1
X_12648_ _13418_/Q _12640_/S _06863_/B _12646_/X _12647_/X vssd1 vssd1 vccd1 vccd1
+ _12649_/B sky130_fd_sc_hd__o221a_1
XFILLER_129_510 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15367_ _15461_/CLK _15367_/D vssd1 vssd1 vccd1 vccd1 _15367_/Q sky130_fd_sc_hd__dfxtp_2
X_12579_ _12575_/X _12576_/X _12594_/S vssd1 vssd1 vccd1 vccd1 _12579_/X sky130_fd_sc_hd__mux2_1
XFILLER_156_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14318_ _15235_/CLK _14318_/D vssd1 vssd1 vccd1 vccd1 _14318_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15298_ _15298_/CLK _15298_/D vssd1 vssd1 vccd1 vccd1 _15298_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_171_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14249_ _15300_/CLK _14249_/D vssd1 vssd1 vccd1 vccd1 _14249_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_125_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08810_ _11877_/A1 _13836_/Q _08811_/S vssd1 vssd1 vccd1 vccd1 _13836_/D sky130_fd_sc_hd__mux2_1
XTAP_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09790_ _14157_/Q _13345_/A0 _09790_/S vssd1 vssd1 vccd1 vccd1 _14157_/D sky130_fd_sc_hd__mux2_1
XFILLER_85_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08741_ _13645_/Q _08523_/Y _08747_/A2 _13542_/Q _08740_/X vssd1 vssd1 vccd1 vccd1
+ _08741_/X sky130_fd_sc_hd__a221o_1
XTAP_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08672_ _13591_/Q _08749_/A2 _08668_/X input34/X vssd1 vssd1 vccd1 vccd1 _08672_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_26_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07623_ _14756_/Q _07629_/A _07622_/Y _08002_/C1 vssd1 vssd1 vccd1 vccd1 _13467_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_93_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_18_clk clkbuf_5_2_0_clk/X vssd1 vssd1 vccd1 vccd1 _15675_/CLK sky130_fd_sc_hd__clkbuf_16
X_07554_ _14738_/Q _07644_/A _07553_/Y _08084_/C1 vssd1 vssd1 vccd1 vccd1 _13449_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_34_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07485_ _13346_/A0 _13410_/Q _07501_/S vssd1 vssd1 vccd1 vccd1 _13410_/D sky130_fd_sc_hd__mux2_1
XFILLER_179_476 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09224_ _14470_/Q _14438_/Q _13859_/Q _14212_/Q _09225_/S0 _09225_/S1 vssd1 vssd1
+ vccd1 vccd1 _09224_/X sky130_fd_sc_hd__mux4_1
XFILLER_148_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09155_ _09419_/A2 _09153_/X _09154_/X _09421_/A1 vssd1 vssd1 vccd1 vccd1 _09155_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_163_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08106_ _13652_/Q _10344_/S _08096_/X _08105_/X vssd1 vssd1 vccd1 vccd1 _13652_/D
+ sky130_fd_sc_hd__a22o_1
X_09086_ _14012_/Q _13980_/Q _09190_/S vssd1 vssd1 vccd1 vccd1 _09086_/X sky130_fd_sc_hd__mux2_1
XFILLER_174_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08037_ _14717_/Q _14718_/Q _08037_/C _08037_/D vssd1 vssd1 vccd1 vccd1 _08038_/S
+ sky130_fd_sc_hd__or4_2
XFILLER_162_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_579 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09988_ _13098_/B2 _14347_/Q _09996_/S vssd1 vssd1 vccd1 vccd1 _14347_/D sky130_fd_sc_hd__mux2_1
XFILLER_131_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08939_ _08519_/A _08937_/X _08938_/X vssd1 vssd1 vccd1 vccd1 _08943_/B sky130_fd_sc_hd__a21o_1
XTAP_3702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11950_ _11933_/X _11934_/X _12594_/S vssd1 vssd1 vccd1 vccd1 _11950_/X sky130_fd_sc_hd__mux2_1
XTAP_3735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_177_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_427 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10901_ _14933_/Q _10951_/B _10900_/Y _11371_/A vssd1 vssd1 vccd1 vccd1 _14933_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_123_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11881_ _15302_/Q _11881_/A1 _11883_/S vssd1 vssd1 vccd1 vccd1 _15302_/D sky130_fd_sc_hd__mux2_1
XFILLER_72_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13620_ _15377_/CLK _13620_/D vssd1 vssd1 vccd1 vccd1 _13620_/Q sky130_fd_sc_hd__dfxtp_1
X_10832_ _14864_/Q _13804_/Q _12932_/S vssd1 vssd1 vccd1 vccd1 _14864_/D sky130_fd_sc_hd__mux2_1
X_13551_ _14495_/CLK _13551_/D vssd1 vssd1 vccd1 vccd1 _13551_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_186_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_644 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10763_ _15427_/Q hold6/A _10764_/S vssd1 vssd1 vccd1 vccd1 _14795_/D sky130_fd_sc_hd__mux2_1
XFILLER_186_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_964 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12502_ _12485_/X _12486_/X _12502_/S vssd1 vssd1 vccd1 vccd1 _12502_/X sky130_fd_sc_hd__mux2_1
XFILLER_185_435 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13482_ _15399_/CLK _13482_/D vssd1 vssd1 vccd1 vccd1 _13482_/Q sky130_fd_sc_hd__dfxtp_2
X_10694_ _15066_/Q _10714_/A2 _10691_/X _10693_/X vssd1 vssd1 vccd1 vccd1 _10694_/X
+ sky130_fd_sc_hd__o22a_2
XFILLER_139_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15221_ _15253_/CLK _15221_/D vssd1 vssd1 vccd1 vccd1 _15221_/Q sky130_fd_sc_hd__dfxtp_1
X_12433_ _12416_/X _12417_/X _12594_/S vssd1 vssd1 vccd1 vccd1 _12433_/X sky130_fd_sc_hd__mux2_1
XFILLER_154_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_72 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15152_ _15253_/CLK _15152_/D vssd1 vssd1 vccd1 vccd1 _15152_/Q sky130_fd_sc_hd__dfxtp_1
X_12364_ _12347_/X _12348_/X _12536_/A vssd1 vssd1 vccd1 vccd1 _12364_/X sky130_fd_sc_hd__mux2_1
XFILLER_165_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14103_ _15273_/CLK _14103_/D vssd1 vssd1 vccd1 vccd1 _14103_/Q sky130_fd_sc_hd__dfxtp_1
X_11315_ _11327_/A _11315_/B vssd1 vssd1 vccd1 vccd1 _11315_/X sky130_fd_sc_hd__or2_1
XFILLER_141_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15083_ _15656_/CLK _15083_/D vssd1 vssd1 vccd1 vccd1 _15083_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12295_ _12278_/X _12279_/X _12617_/S vssd1 vssd1 vccd1 vccd1 _12295_/X sky130_fd_sc_hd__mux2_1
XFILLER_113_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14034_ _15324_/CLK _14034_/D vssd1 vssd1 vccd1 vccd1 _14034_/Q sky130_fd_sc_hd__dfxtp_1
X_11246_ _11283_/A _08319_/X _11245_/Y _08233_/B vssd1 vssd1 vccd1 vccd1 _11246_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_180_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11177_ _11380_/A _11177_/B vssd1 vssd1 vccd1 vccd1 _11177_/Y sky130_fd_sc_hd__nor2_1
XFILLER_110_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10128_ _14514_/Q _14762_/Q _10131_/S vssd1 vssd1 vccd1 vccd1 _14514_/D sky130_fd_sc_hd__mux2_1
XFILLER_48_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10059_ _14416_/Q _13104_/B2 _10059_/S vssd1 vssd1 vccd1 vccd1 _14416_/D sky130_fd_sc_hd__mux2_1
X_14936_ _15000_/CLK _14936_/D vssd1 vssd1 vccd1 vccd1 _14936_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_235 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14867_ _15620_/CLK _14867_/D vssd1 vssd1 vccd1 vccd1 _14867_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13818_ _15220_/CLK _13818_/D vssd1 vssd1 vccd1 vccd1 _13818_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14798_ _14861_/CLK _14798_/D vssd1 vssd1 vccd1 vccd1 _14798_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13749_ _14868_/CLK _13749_/D vssd1 vssd1 vccd1 vccd1 _13749_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_188_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07270_ _07270_/A _07270_/B _07270_/C vssd1 vssd1 vccd1 vccd1 _07274_/C sky130_fd_sc_hd__or3_1
X_15419_ _15638_/CLK _15419_/D vssd1 vssd1 vccd1 vccd1 _15419_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_117_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_176_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_7_clk clkbuf_5_1_0_clk/X vssd1 vssd1 vccd1 vccd1 _14415_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_172_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09911_ _13331_/A0 _14272_/Q _09925_/S vssd1 vssd1 vccd1 vccd1 _14272_/D sky130_fd_sc_hd__mux2_1
XFILLER_176_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_171_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout605 _12472_/S vssd1 vssd1 vccd1 vccd1 _12476_/S sky130_fd_sc_hd__buf_12
Xfanout616 _12545_/S vssd1 vssd1 vccd1 vccd1 _12407_/S sky130_fd_sc_hd__buf_12
XTAP_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09842_ _14206_/Q _13329_/A0 _09858_/S vssd1 vssd1 vccd1 vccd1 _14206_/D sky130_fd_sc_hd__mux2_1
XFILLER_112_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout627 _10507_/A1 vssd1 vssd1 vccd1 vccd1 _08244_/A sky130_fd_sc_hd__buf_8
XTAP_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout638 fanout647/X vssd1 vssd1 vccd1 vccd1 _12832_/C1 sky130_fd_sc_hd__buf_12
XFILLER_98_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09773_ _14140_/Q _13328_/A0 _09790_/S vssd1 vssd1 vccd1 vccd1 _14140_/D sky130_fd_sc_hd__mux2_1
XTAP_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06985_ _14586_/Q _06987_/D vssd1 vssd1 vccd1 vccd1 _08753_/D sky130_fd_sc_hd__nand2_1
XTAP_3009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08724_ _13574_/Q _08724_/B _08724_/C vssd1 vssd1 vccd1 vccd1 _08724_/X sky130_fd_sc_hd__and3_1
XFILLER_160_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08655_ _13593_/Q _08691_/A2 _08685_/A2 _13554_/Q _08654_/X vssd1 vssd1 vccd1 vccd1
+ _08659_/B sky130_fd_sc_hd__a221o_1
XFILLER_26_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07606_ _13463_/Q _07610_/C vssd1 vssd1 vccd1 vccd1 _07607_/B sky130_fd_sc_hd__xnor2_1
XFILLER_54_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08586_ _13782_/Q _08585_/X _08626_/S vssd1 vssd1 vccd1 vccd1 _13782_/D sky130_fd_sc_hd__mux2_1
XFILLER_41_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07537_ _07504_/C _07658_/B vssd1 vssd1 vccd1 vccd1 _07783_/B sky130_fd_sc_hd__nand2b_1
XFILLER_23_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07468_ _14757_/Q _07467_/X _07500_/S vssd1 vssd1 vccd1 vccd1 _07468_/X sky130_fd_sc_hd__mux2_8
XFILLER_22_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09207_ _13890_/Q _09445_/A2 _09522_/B1 _14405_/Q _09437_/A1 vssd1 vssd1 vccd1 vccd1
+ _09207_/X sky130_fd_sc_hd__a221o_1
XFILLER_33_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07399_ _13655_/Q _07499_/A2 _07499_/B1 _14683_/Q _07398_/X vssd1 vssd1 vccd1 vccd1
+ _07399_/X sky130_fd_sc_hd__a221o_1
XFILLER_148_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_37 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09138_ _14368_/Q _15184_/Q _13823_/Q _14562_/Q _09425_/S _09427_/A1 vssd1 vssd1
+ vccd1 vccd1 _09139_/B sky130_fd_sc_hd__mux4_1
XFILLER_5_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09069_ _14364_/Q _15180_/Q _13819_/Q _14558_/Q _09073_/S _09234_/S1 vssd1 vssd1
+ vccd1 vccd1 _09070_/B sky130_fd_sc_hd__mux4_1
XFILLER_123_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11100_ _11347_/A _11098_/X _11000_/X _11307_/A vssd1 vssd1 vccd1 vccd1 _11100_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_162_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12080_ _12080_/A _12080_/B vssd1 vssd1 vccd1 vccd1 _12080_/X sky130_fd_sc_hd__and2_1
XFILLER_118_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11031_ _11031_/A vssd1 vssd1 vccd1 vccd1 _11031_/Y sky130_fd_sc_hd__inv_2
XFILLER_77_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12982_ _07424_/X _13024_/A2 _12981_/X _13024_/B2 vssd1 vssd1 vccd1 vccd1 _12982_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_3521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14721_ _15670_/CLK _14721_/D vssd1 vssd1 vccd1 vccd1 _14721_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_3554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11933_ _14520_/Q _14133_/Q _14165_/Q _14101_/Q _12407_/S _12406_/A vssd1 vssd1 vccd1
+ vccd1 _11933_/X sky130_fd_sc_hd__mux4_1
XFILLER_57_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14652_ _15623_/CLK _14652_/D vssd1 vssd1 vccd1 vccd1 _14652_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11864_ _15285_/Q _13331_/A0 _11878_/S vssd1 vssd1 vccd1 vccd1 _15285_/D sky130_fd_sc_hd__mux2_1
XFILLER_73_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13603_ _15378_/CLK _13603_/D vssd1 vssd1 vccd1 vccd1 _13603_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_2886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10815_ _14847_/Q _07261_/A _10868_/S vssd1 vssd1 vccd1 vccd1 _14847_/D sky130_fd_sc_hd__mux2_1
XTAP_2897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14583_ _15616_/CLK _14583_/D vssd1 vssd1 vccd1 vccd1 _14583_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11795_ _15218_/Q _11861_/A1 _11816_/S vssd1 vssd1 vccd1 vccd1 _15218_/D sky130_fd_sc_hd__mux2_1
XFILLER_129_1091 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13534_ _14511_/CLK _13534_/D vssd1 vssd1 vccd1 vccd1 _13534_/Q sky130_fd_sc_hd__dfxtp_1
X_10746_ _15410_/Q _14778_/Q _10759_/S vssd1 vssd1 vccd1 vccd1 _14778_/D sky130_fd_sc_hd__mux2_1
XFILLER_41_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13465_ _15385_/CLK _13465_/D vssd1 vssd1 vccd1 vccd1 _13465_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_186_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10677_ _15014_/Q _10717_/A2 _10652_/B _15031_/Q _10717_/C1 vssd1 vssd1 vccd1 vccd1
+ _10677_/X sky130_fd_sc_hd__a221o_1
XFILLER_139_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15204_ _15615_/CLK _15204_/D vssd1 vssd1 vccd1 vccd1 _15204_/Q sky130_fd_sc_hd__dfxtp_1
X_12416_ _14541_/Q _14154_/Q _14186_/Q _14122_/Q _12430_/S _12563_/A vssd1 vssd1 vccd1
+ vccd1 _12416_/X sky130_fd_sc_hd__mux4_1
XFILLER_173_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13396_ _15659_/CLK _13396_/D vssd1 vssd1 vccd1 vccd1 _13396_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_126_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15135_ _15670_/CLK _15135_/D vssd1 vssd1 vccd1 vccd1 _15135_/Q sky130_fd_sc_hd__dfxtp_1
X_12347_ _14538_/Q _14151_/Q _14183_/Q _14119_/Q _12541_/S _12540_/A vssd1 vssd1 vccd1
+ vccd1 _12347_/X sky130_fd_sc_hd__mux4_1
XFILLER_5_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_684 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15066_ _15422_/CLK _15066_/D vssd1 vssd1 vccd1 vccd1 _15066_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_142_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12278_ _14535_/Q _14148_/Q _14180_/Q _14116_/Q _12614_/S _12383_/A vssd1 vssd1 vccd1
+ vccd1 _12278_/X sky130_fd_sc_hd__mux4_1
XFILLER_4_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14017_ _15658_/CLK _14017_/D vssd1 vssd1 vccd1 vccd1 _14017_/Q sky130_fd_sc_hd__dfxtp_1
X_11229_ _10527_/A _15017_/Q _11237_/S vssd1 vssd1 vccd1 vccd1 _15017_/D sky130_fd_sc_hd__mux2_1
XFILLER_150_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06770_ _14900_/Q _14899_/Q vssd1 vssd1 vccd1 vccd1 _08121_/A sky130_fd_sc_hd__or2_2
XFILLER_49_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14919_ _15552_/CLK _14919_/D vssd1 vssd1 vccd1 vccd1 _14919_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08440_ _13750_/Q _12878_/S _08426_/B _08439_/X vssd1 vssd1 vccd1 vccd1 _13750_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_63_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_5_7_0_clk clkbuf_5_7_0_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_5_7_0_clk/X sky130_fd_sc_hd__clkbuf_8
XFILLER_23_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08371_ _11025_/A _13195_/B vssd1 vssd1 vccd1 vccd1 _10991_/B sky130_fd_sc_hd__nor2_1
XFILLER_149_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07322_ _13911_/Q _15498_/Q _07339_/S vssd1 vssd1 vccd1 vccd1 _07322_/X sky130_fd_sc_hd__mux2_8
XFILLER_182_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07253_ _13924_/Q _15511_/Q _07334_/S vssd1 vssd1 vccd1 vccd1 _07261_/A sky130_fd_sc_hd__mux2_8
XFILLER_104_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07184_ _15358_/Q _15065_/Q _07188_/S vssd1 vssd1 vccd1 vccd1 _07184_/X sky130_fd_sc_hd__mux2_8
XFILLER_118_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout402 _12764_/S vssd1 vssd1 vccd1 vccd1 _12728_/S sky130_fd_sc_hd__buf_12
Xfanout413 _10983_/X vssd1 vssd1 vccd1 vccd1 _11164_/S sky130_fd_sc_hd__buf_6
Xfanout424 _09445_/A2 vssd1 vssd1 vccd1 vccd1 _09231_/A2 sky130_fd_sc_hd__buf_12
XFILLER_48_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_271 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout435 _08223_/X vssd1 vssd1 vccd1 vccd1 _08232_/A sky130_fd_sc_hd__clkbuf_16
Xfanout446 _10615_/S vssd1 vssd1 vccd1 vccd1 _10730_/S sky130_fd_sc_hd__buf_12
Xfanout457 _10244_/S vssd1 vssd1 vccd1 vccd1 _10665_/S sky130_fd_sc_hd__buf_6
X_09825_ _14191_/Q _13347_/A0 _09828_/S vssd1 vssd1 vccd1 vccd1 _14191_/D sky130_fd_sc_hd__mux2_1
XFILLER_86_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout468 _12503_/A1 vssd1 vssd1 vccd1 vccd1 _12273_/A1 sky130_fd_sc_hd__buf_12
XFILLER_171_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout479 _12559_/A vssd1 vssd1 vccd1 vccd1 _12617_/S sky130_fd_sc_hd__buf_12
XFILLER_86_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09756_ _14124_/Q _11877_/A1 _09757_/S vssd1 vssd1 vccd1 vccd1 _14124_/D sky130_fd_sc_hd__mux2_1
X_06968_ _06716_/Y _13495_/Q _06718_/Y _13494_/Q vssd1 vssd1 vccd1 vccd1 _06969_/D
+ sky130_fd_sc_hd__o22ai_2
X_08707_ _13483_/Q _08747_/B1 _08750_/B1 _13618_/Q vssd1 vssd1 vccd1 vccd1 _08707_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_39_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09687_ _14058_/Q _13342_/A0 _09695_/S vssd1 vssd1 vccd1 vccd1 _14058_/D sky130_fd_sc_hd__mux2_1
XFILLER_66_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06899_ _15373_/Q _06744_/Y _15372_/Q _06747_/Y _06898_/X vssd1 vssd1 vccd1 vccd1
+ _06899_/X sky130_fd_sc_hd__o221a_1
XTAP_2138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08638_ _14502_/Q _08693_/A2 _08635_/X _08636_/X _08637_/X vssd1 vssd1 vccd1 vccd1
+ _08638_/X sky130_fd_sc_hd__a2111o_4
XTAP_1415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08569_ _13535_/Q _08750_/A2 _08747_/B1 _13503_/Q _08568_/X vssd1 vssd1 vccd1 vccd1
+ _08569_/X sky130_fd_sc_hd__a221o_1
X_10600_ _14738_/Q _10599_/X _10615_/S vssd1 vssd1 vccd1 vccd1 _14738_/D sky130_fd_sc_hd__mux2_1
XFILLER_168_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11580_ _11549_/B _11576_/Y _11578_/X _11579_/Y vssd1 vssd1 vccd1 vccd1 _11586_/A
+ sky130_fd_sc_hd__a211o_2
XFILLER_70_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10531_ _11584_/A _11582_/A vssd1 vssd1 vccd1 vccd1 _10532_/B sky130_fd_sc_hd__and2b_1
XFILLER_183_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13250_ _15583_/Q _13252_/B _13248_/Y _13249_/X vssd1 vssd1 vccd1 vccd1 _15583_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_155_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10462_ _10462_/A _10462_/B vssd1 vssd1 vccd1 vccd1 _10470_/C sky130_fd_sc_hd__nand2_1
XFILLER_6_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12201_ _12477_/A1 _12200_/X _12500_/B1 vssd1 vssd1 vccd1 vccd1 _12201_/X sky130_fd_sc_hd__a21o_1
XFILLER_108_343 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13181_ _13217_/A _11419_/A _13241_/A2 vssd1 vssd1 vccd1 vccd1 _13181_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_108_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10393_ _13178_/B _13177_/A vssd1 vssd1 vccd1 vccd1 _10395_/A sky130_fd_sc_hd__nand2b_1
XFILLER_123_313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_1084 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12132_ _12477_/A1 _12131_/X _12500_/B1 vssd1 vssd1 vccd1 vccd1 _12132_/X sky130_fd_sc_hd__a21o_1
XFILLER_124_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12063_ _12500_/A1 _12062_/X _12468_/A1 vssd1 vssd1 vccd1 vccd1 _12063_/X sky130_fd_sc_hd__a21o_1
XFILLER_49_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11014_ _11023_/A _11633_/A _11013_/X vssd1 vssd1 vccd1 vccd1 _11079_/B sky130_fd_sc_hd__o21ai_1
XFILLER_77_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_240_clk clkbuf_5_5_0_clk/X vssd1 vssd1 vccd1 vccd1 _15279_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_65_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12965_ _15468_/Q _13139_/S _13025_/B1 _12964_/X vssd1 vssd1 vccd1 vccd1 _15468_/D
+ sky130_fd_sc_hd__a22o_1
XTAP_4096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_875 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14704_ _15644_/CLK _14704_/D vssd1 vssd1 vccd1 vccd1 _14704_/Q sky130_fd_sc_hd__dfxtp_1
X_11916_ _08405_/B _11913_/X _08405_/C vssd1 vssd1 vccd1 vccd1 _11916_/X sky130_fd_sc_hd__o21a_1
XTAP_3384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12896_ _15424_/Q _15609_/Q _12929_/S vssd1 vssd1 vccd1 vccd1 _15424_/D sky130_fd_sc_hd__mux2_1
XTAP_2650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14635_ _15638_/CLK _14635_/D vssd1 vssd1 vccd1 vccd1 _14635_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11847_ _15269_/Q _11847_/A1 _11850_/S vssd1 vssd1 vccd1 vccd1 _15269_/D sky130_fd_sc_hd__mux2_1
XTAP_2694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14566_ _15289_/CLK _14566_/D vssd1 vssd1 vccd1 vccd1 _14566_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11778_ _10563_/B _11776_/X _11777_/Y _10344_/S _15204_/Q vssd1 vssd1 vccd1 vccd1
+ _15204_/D sky130_fd_sc_hd__a32o_1
X_13517_ _13798_/CLK _13517_/D vssd1 vssd1 vccd1 vccd1 _13517_/Q sky130_fd_sc_hd__dfxtp_1
X_10729_ _15073_/Q _10734_/A2 _10726_/X _10728_/X vssd1 vssd1 vccd1 vccd1 _10729_/X
+ sky130_fd_sc_hd__o22a_2
X_14497_ _15374_/CLK _14497_/D vssd1 vssd1 vccd1 vccd1 _14497_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_173_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13448_ _15372_/CLK _13448_/D vssd1 vssd1 vccd1 vccd1 _13448_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_174_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13379_ _14482_/Q vssd1 vssd1 vccd1 vccd1 _14482_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_55_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_791 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15118_ _15133_/CLK _15118_/D vssd1 vssd1 vccd1 vccd1 _15118_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07940_ _13550_/Q _07946_/D vssd1 vssd1 vccd1 vccd1 _07940_/X sky130_fd_sc_hd__or2_1
X_15049_ _15613_/CLK _15049_/D vssd1 vssd1 vccd1 vccd1 _15049_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_130_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07871_ _07884_/C _07870_/Y _07874_/A vssd1 vssd1 vccd1 vccd1 _07871_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_68_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_231_clk clkbuf_5_4_0_clk/X vssd1 vssd1 vccd1 vccd1 _14530_/CLK sky130_fd_sc_hd__clkbuf_16
X_09610_ _13984_/Q _13078_/B2 _09627_/S vssd1 vssd1 vccd1 vccd1 _13984_/D sky130_fd_sc_hd__mux2_1
XFILLER_96_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06822_ _13574_/Q _13575_/Q input34/X vssd1 vssd1 vccd1 vccd1 _06825_/C sky130_fd_sc_hd__nand3_4
XFILLER_3_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_138 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09541_ _15304_/Q _15272_/Q _15240_/Q _15171_/Q _09469_/S _09546_/S1 vssd1 vssd1
+ vccd1 vccd1 _09541_/X sky130_fd_sc_hd__mux4_1
X_06753_ _14487_/Q vssd1 vssd1 vccd1 vccd1 _06753_/Y sky130_fd_sc_hd__inv_2
XFILLER_24_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09472_ _08510_/B _09468_/X _09471_/X _09467_/X vssd1 vssd1 vccd1 vccd1 _09472_/X
+ sky130_fd_sc_hd__a211o_1
X_06684_ input35/X vssd1 vssd1 vccd1 vccd1 _06684_/Y sky130_fd_sc_hd__inv_2
XFILLER_64_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08423_ _08465_/B _08773_/B _08421_/Y _12906_/S _14614_/Q vssd1 vssd1 vccd1 vccd1
+ _08423_/X sky130_fd_sc_hd__o311a_1
XFILLER_180_1019 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08354_ _11037_/A _08361_/B vssd1 vssd1 vccd1 vccd1 _10991_/A sky130_fd_sc_hd__nor2_1
XFILLER_149_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07305_ _13915_/Q _15502_/Q _07334_/S vssd1 vssd1 vccd1 vccd1 _07306_/A sky130_fd_sc_hd__mux2_8
X_08285_ _10507_/A1 _13769_/Q _15403_/Q _10515_/B2 vssd1 vssd1 vccd1 vccd1 _08285_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_137_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07236_ _13929_/Q _15516_/Q _07334_/S vssd1 vssd1 vccd1 vccd1 _07237_/A sky130_fd_sc_hd__mux2_8
XFILLER_117_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07167_ _15341_/Q _15048_/Q _07193_/S vssd1 vssd1 vccd1 vccd1 _07167_/X sky130_fd_sc_hd__mux2_8
XFILLER_161_920 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_471 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07098_ _07097_/X _14765_/Q _07098_/S vssd1 vssd1 vccd1 vccd1 _13611_/D sky130_fd_sc_hd__mux2_1
XFILLER_161_975 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout210 _09629_/Y vssd1 vssd1 vccd1 vccd1 _09661_/S sky130_fd_sc_hd__buf_12
XFILLER_132_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_496 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout221 _08040_/X vssd1 vssd1 vccd1 vccd1 _08072_/S sky130_fd_sc_hd__buf_12
XFILLER_114_891 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout232 _07614_/A vssd1 vssd1 vccd1 vccd1 _07651_/A sky130_fd_sc_hd__buf_4
Xfanout243 _09831_/Y vssd1 vssd1 vccd1 vccd1 _09858_/S sky130_fd_sc_hd__buf_12
Xfanout254 _08189_/Y vssd1 vssd1 vccd1 vccd1 _08221_/S sky130_fd_sc_hd__buf_12
XFILLER_113_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout265 _08532_/Y vssd1 vssd1 vccd1 vccd1 _08750_/B1 sky130_fd_sc_hd__buf_12
XFILLER_115_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout276 _13130_/B1 vssd1 vssd1 vccd1 vccd1 _08540_/B sky130_fd_sc_hd__buf_12
X_09808_ _14174_/Q _13074_/B2 _09823_/S vssd1 vssd1 vccd1 vccd1 _14174_/D sky130_fd_sc_hd__mux2_1
XFILLER_47_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout287 _13110_/B2 vssd1 vssd1 vccd1 vccd1 _13348_/A0 sky130_fd_sc_hd__clkbuf_4
Xclkbuf_leaf_222_clk clkbuf_opt_1_0_clk/X vssd1 vssd1 vccd1 vccd1 _15530_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_115_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout298 _07472_/X vssd1 vssd1 vccd1 vccd1 _13343_/A0 sky130_fd_sc_hd__buf_6
XFILLER_28_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09739_ _14107_/Q _13327_/A0 _09757_/S vssd1 vssd1 vccd1 vccd1 _14107_/D sky130_fd_sc_hd__mux2_1
XFILLER_55_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12750_ _13432_/Q _12749_/X _12764_/S vssd1 vssd1 vccd1 vccd1 _12750_/X sky130_fd_sc_hd__mux2_1
XTAP_1201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11701_ _13343_/A0 _15132_/Q _11703_/S vssd1 vssd1 vccd1 vccd1 _15132_/D sky130_fd_sc_hd__mux2_1
XFILLER_187_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12681_ _12688_/B _12681_/B vssd1 vssd1 vccd1 vccd1 _12681_/Y sky130_fd_sc_hd__nor2_1
XFILLER_15_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14420_ _14420_/CLK _14420_/D vssd1 vssd1 vccd1 vccd1 _14420_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11632_ _11632_/A _11632_/B vssd1 vssd1 vccd1 vccd1 _11633_/B sky130_fd_sc_hd__xnor2_2
XFILLER_168_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14351_ _15199_/CLK _14351_/D vssd1 vssd1 vccd1 vccd1 _14351_/Q sky130_fd_sc_hd__dfxtp_1
X_11563_ _11563_/A _11563_/B vssd1 vssd1 vccd1 vccd1 _11564_/B sky130_fd_sc_hd__or2_1
XFILLER_11_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13302_ _12739_/X _15634_/Q _13309_/A vssd1 vssd1 vccd1 vccd1 _15634_/D sky130_fd_sc_hd__mux2_1
XFILLER_6_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10514_ _07260_/A _10360_/B _10513_/X vssd1 vssd1 vccd1 vccd1 _11536_/C sky130_fd_sc_hd__a21oi_4
X_14282_ _15295_/CLK _14282_/D vssd1 vssd1 vccd1 vccd1 _14282_/Q sky130_fd_sc_hd__dfxtp_1
X_11494_ _11493_/A _11505_/D _11474_/S vssd1 vssd1 vccd1 vccd1 _11494_/X sky130_fd_sc_hd__o21ba_1
XFILLER_10_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13233_ _13233_/A _13233_/B vssd1 vssd1 vccd1 vccd1 _13233_/Y sky130_fd_sc_hd__nand2_1
XFILLER_170_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_61 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10445_ _07210_/A _10360_/B _10444_/X vssd1 vssd1 vccd1 vccd1 _11600_/A sky130_fd_sc_hd__a21oi_4
XFILLER_170_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13164_ _15555_/Q _13252_/B _13162_/Y _13163_/X vssd1 vssd1 vccd1 vccd1 _15555_/D
+ sky130_fd_sc_hd__a22o_1
X_10376_ _14767_/Q _13794_/Q _13762_/Q _14766_/Q vssd1 vssd1 vccd1 vccd1 _10376_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_123_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12115_ _14238_/Q _14270_/Q _14302_/Q _14334_/Q _12489_/S0 _12489_/S1 vssd1 vssd1
+ vccd1 vccd1 _12115_/X sky130_fd_sc_hd__mux4_1
X_13095_ _15515_/Q _13129_/A _13042_/A _13094_/X vssd1 vssd1 vccd1 vccd1 _15515_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_124_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12046_ _14235_/Q _14267_/Q _14299_/Q _14331_/Q _12154_/S _12253_/S1 vssd1 vssd1
+ vccd1 vccd1 _12046_/X sky130_fd_sc_hd__mux4_1
XFILLER_46_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_775 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_213_clk clkbuf_5_19_0_clk/X vssd1 vssd1 vccd1 vccd1 _15666_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_133_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_1087 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13997_ _15088_/CLK _13997_/D vssd1 vssd1 vccd1 vccd1 _13997_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12948_ _10584_/X _14863_/Q _13038_/S vssd1 vssd1 vccd1 vccd1 _12948_/X sky130_fd_sc_hd__mux2_2
XTAP_3181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12879_ _15407_/Q _15592_/Q _12917_/S vssd1 vssd1 vccd1 vccd1 _15407_/D sky130_fd_sc_hd__mux2_1
X_15667_ _15667_/CLK _15667_/D vssd1 vssd1 vccd1 vccd1 _15667_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14618_ _14861_/CLK _14618_/D vssd1 vssd1 vccd1 vccd1 _14618_/Q sky130_fd_sc_hd__dfxtp_1
X_15598_ _15599_/CLK _15598_/D vssd1 vssd1 vccd1 vccd1 _15598_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_883 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14549_ _15680_/CLK _14549_/D vssd1 vssd1 vccd1 vccd1 _14549_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_174_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08070_ _14763_/Q _13641_/Q _08072_/S vssd1 vssd1 vccd1 vccd1 _13641_/D sky130_fd_sc_hd__mux2_1
XFILLER_101_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07021_ _14619_/Q _14651_/Q _07096_/S vssd1 vssd1 vccd1 vccd1 _07021_/X sky130_fd_sc_hd__mux2_1
XFILLER_143_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08972_ _15277_/Q _15245_/Q _15213_/Q _15144_/Q _09225_/S0 _09225_/S1 vssd1 vssd1
+ vccd1 vccd1 _08972_/X sky130_fd_sc_hd__mux4_1
X_07923_ _14738_/Q _08012_/A2 _07922_/Y vssd1 vssd1 vccd1 vccd1 _13545_/D sky130_fd_sc_hd__o21a_1
Xclkbuf_leaf_204_clk clkbuf_5_16_0_clk/X vssd1 vssd1 vccd1 vccd1 _14572_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_84_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07854_ _14752_/Q _07874_/A _07853_/X _07987_/C1 vssd1 vssd1 vccd1 vccd1 _13527_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_111_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06805_ _13732_/Q _06669_/Y _08405_/C _06664_/Y _06804_/X vssd1 vssd1 vccd1 vccd1
+ _06806_/C sky130_fd_sc_hd__a221oi_1
XFILLER_56_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07785_ _14734_/Q _07816_/A _07784_/Y _12832_/C1 vssd1 vssd1 vccd1 vccd1 _13509_/D
+ sky130_fd_sc_hd__o211a_1
X_09524_ _09524_/A _09524_/B _09524_/C vssd1 vssd1 vccd1 vccd1 _09524_/X sky130_fd_sc_hd__and3_1
X_06736_ _14494_/Q vssd1 vssd1 vccd1 vccd1 _06736_/Y sky130_fd_sc_hd__inv_2
XFILLER_25_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09455_ _13902_/Q _13123_/B _08512_/B _14417_/Q _13123_/A vssd1 vssd1 vccd1 vccd1
+ _09455_/X sky130_fd_sc_hd__a221o_1
X_06667_ _14596_/Q vssd1 vssd1 vccd1 vccd1 _08765_/A sky130_fd_sc_hd__inv_2
XPHY_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08406_ _12379_/A _08406_/B vssd1 vssd1 vccd1 vccd1 _12946_/B sky130_fd_sc_hd__nor2_2
XFILLER_169_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09386_ _15131_/Q _09558_/A2 _08520_/B _09385_/X vssd1 vssd1 vccd1 vccd1 _09386_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_51_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_16 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08337_ _08316_/Y _08336_/Y _11318_/S vssd1 vssd1 vccd1 vccd1 _08337_/X sky130_fd_sc_hd__mux2_1
XFILLER_177_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08268_ _11351_/C1 _08249_/Y _08292_/B _08232_/A _13715_/Q vssd1 vssd1 vccd1 vccd1
+ _13715_/D sky130_fd_sc_hd__a32o_1
XFILLER_153_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07219_ _13931_/Q _15518_/Q _07339_/S vssd1 vssd1 vccd1 vccd1 _07219_/X sky130_fd_sc_hd__mux2_8
X_08199_ _13690_/Q _13328_/A0 _08216_/S vssd1 vssd1 vccd1 vccd1 _13690_/D sky130_fd_sc_hd__mux2_1
XFILLER_152_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10230_ _14615_/Q _14768_/Q _10735_/S vssd1 vssd1 vccd1 vccd1 _14615_/D sky130_fd_sc_hd__mux2_1
XFILLER_105_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10161_ _14546_/Q _13347_/A0 _10164_/S vssd1 vssd1 vccd1 vccd1 _14546_/D sky130_fd_sc_hd__mux2_1
XFILLER_126_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_966 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10092_ _14448_/Q _13345_/A0 _10092_/S vssd1 vssd1 vccd1 vccd1 _14448_/D sky130_fd_sc_hd__mux2_1
XFILLER_87_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13920_ _15332_/CLK _13920_/D vssd1 vssd1 vccd1 vccd1 _13920_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13851_ _15657_/CLK _13851_/D vssd1 vssd1 vccd1 vccd1 _13851_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_74_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12802_ _06861_/Y _12799_/X _12800_/X _12801_/X vssd1 vssd1 vccd1 vccd1 _12802_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_56_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13782_ _15393_/CLK _13782_/D vssd1 vssd1 vccd1 vccd1 _13782_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_16_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10994_ _10988_/Y _10993_/Y _11252_/A vssd1 vssd1 vccd1 vccd1 _10994_/X sky130_fd_sc_hd__mux2_2
XFILLER_43_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12733_ _12745_/C _12733_/B vssd1 vssd1 vccd1 vccd1 _12733_/Y sky130_fd_sc_hd__nor2_1
XTAP_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15521_ _15525_/CLK _15521_/D vssd1 vssd1 vccd1 vccd1 _15521_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15452_ _15452_/CLK _15452_/D vssd1 vssd1 vccd1 vccd1 _15452_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12664_ _15343_/Q _12759_/B _12663_/X _12832_/C1 vssd1 vssd1 vccd1 vccd1 _15343_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_188_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14403_ _15331_/CLK _14403_/D vssd1 vssd1 vccd1 vccd1 _14403_/Q sky130_fd_sc_hd__dfxtp_1
X_11615_ _13217_/A _11610_/A _11610_/B vssd1 vssd1 vccd1 vccd1 _11616_/B sky130_fd_sc_hd__a21boi_4
XFILLER_89_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15383_ _15383_/CLK _15383_/D vssd1 vssd1 vccd1 vccd1 _15383_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_156_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12595_ _12595_/A1 _12594_/X _12593_/X _12618_/C1 vssd1 vssd1 vccd1 vccd1 _12596_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_11_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14334_ _15235_/CLK _14334_/D vssd1 vssd1 vccd1 vccd1 _14334_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_184_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11546_ _11546_/A _11546_/B _11546_/C vssd1 vssd1 vccd1 vccd1 _11546_/X sky130_fd_sc_hd__and3_1
XFILLER_128_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14265_ _15278_/CLK _14265_/D vssd1 vssd1 vccd1 vccd1 _14265_/Q sky130_fd_sc_hd__dfxtp_1
X_11477_ _13233_/A _11496_/C vssd1 vssd1 vccd1 vccd1 _11478_/B sky130_fd_sc_hd__or2_2
XFILLER_171_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13216_ _15572_/Q _13241_/A2 _13214_/Y _13215_/Y vssd1 vssd1 vccd1 vccd1 _15572_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_125_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10428_ _11349_/C _11632_/A vssd1 vssd1 vccd1 vccd1 _10429_/B sky130_fd_sc_hd__nand2_1
X_14196_ _15273_/CLK _14196_/D vssd1 vssd1 vccd1 vccd1 _14196_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13147_ _13125_/B _15545_/Q _13154_/S vssd1 vssd1 vccd1 vccd1 _15545_/D sky130_fd_sc_hd__mux2_1
X_10359_ _13195_/B _11475_/A vssd1 vssd1 vccd1 vccd1 _10366_/B sky130_fd_sc_hd__nor2_1
XTAP_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13078_ _12984_/X _13104_/A2 _13104_/B1 _13078_/B2 vssd1 vssd1 vccd1 vccd1 _13078_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_97_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12029_ _15279_/Q _15247_/Q _15215_/Q _15146_/Q _12079_/S _12080_/A vssd1 vssd1 vccd1
+ vccd1 _12030_/B sky130_fd_sc_hd__mux4_1
XFILLER_18_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07570_ _07571_/B _07567_/B _07571_/A vssd1 vssd1 vccd1 vccd1 _07570_/X sky130_fd_sc_hd__o21a_1
X_09240_ _14373_/Q _15189_/Q _13828_/Q _14567_/Q _09535_/S _08494_/B vssd1 vssd1 vccd1
+ vccd1 _09241_/B sky130_fd_sc_hd__mux4_1
XFILLER_167_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09171_ _09448_/S1 _09169_/X _09170_/X vssd1 vssd1 vccd1 vccd1 _09172_/C sky130_fd_sc_hd__a21o_1
XFILLER_159_371 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08122_ _08133_/S _06759_/Y _08093_/B vssd1 vssd1 vccd1 vccd1 _08122_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_30_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08053_ _14746_/Q _13624_/Q _08066_/S vssd1 vssd1 vccd1 vccd1 _13624_/D sky130_fd_sc_hd__mux2_1
XFILLER_179_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07004_ _14717_/Q _08074_/A _10099_/B vssd1 vssd1 vccd1 vccd1 _07004_/X sky130_fd_sc_hd__and3_4
XFILLER_150_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_923 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08955_ _14231_/Q _14263_/Q _14295_/Q _14327_/Q _09230_/S _09234_/S1 vssd1 vssd1
+ vccd1 vccd1 _08955_/X sky130_fd_sc_hd__mux4_1
XFILLER_5_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07906_ _13541_/Q _07913_/D vssd1 vssd1 vccd1 vccd1 _07906_/X sky130_fd_sc_hd__or2_1
XFILLER_57_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08886_ _14356_/Q _15172_/Q _13811_/Q _14550_/Q _09225_/S0 _09225_/S1 vssd1 vssd1
+ vccd1 vccd1 _08887_/B sky130_fd_sc_hd__mux4_1
XFILLER_56_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07837_ _13523_/Q _07837_/B vssd1 vssd1 vccd1 vccd1 _07837_/Y sky130_fd_sc_hd__nor2_1
XTAP_3928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07768_ _13506_/Q _07769_/B vssd1 vssd1 vccd1 vccd1 _07768_/Y sky130_fd_sc_hd__nor2_1
XFILLER_147_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09507_ _14032_/Q _14000_/Q _09535_/S vssd1 vssd1 vccd1 vccd1 _09507_/X sky130_fd_sc_hd__mux2_1
XFILLER_53_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06719_ _15385_/Q vssd1 vssd1 vccd1 vccd1 _06719_/Y sky130_fd_sc_hd__inv_2
XFILLER_112_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07699_ _14744_/Q _07713_/A _07698_/Y _07949_/C1 vssd1 vssd1 vccd1 vccd1 _13487_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_24_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09438_ _14480_/Q _14448_/Q _13869_/Q _14222_/Q _09438_/S0 _09448_/S1 vssd1 vssd1
+ vccd1 vccd1 _09438_/X sky130_fd_sc_hd__mux4_1
XPHY_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09369_ _15296_/Q _15264_/Q _15232_/Q _15163_/Q _09535_/S _08494_/B vssd1 vssd1 vccd1
+ vccd1 _09369_/X sky130_fd_sc_hd__mux4_1
XFILLER_36_1072 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11400_ _11421_/A _11400_/B vssd1 vssd1 vccd1 vccd1 _11404_/A sky130_fd_sc_hd__nor2_2
XFILLER_162_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12380_ _13896_/Q _14411_/Q _12518_/S vssd1 vssd1 vccd1 vccd1 _12380_/X sky130_fd_sc_hd__mux2_1
XANTENNA_70 _07139_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_81 _07114_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11331_ _11023_/A wire360/X _10963_/B vssd1 vssd1 vccd1 vccd1 _11331_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_21_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_92 _08507_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_180_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_1097 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_536 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14050_ _15088_/CLK _14050_/D vssd1 vssd1 vccd1 vccd1 _14050_/Q sky130_fd_sc_hd__dfxtp_1
X_11262_ _11344_/A _11262_/B vssd1 vssd1 vccd1 vccd1 _11262_/Y sky130_fd_sc_hd__nor2_1
XFILLER_106_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13001_ _15480_/Q _10892_/B _13116_/C _13000_/X vssd1 vssd1 vccd1 vccd1 _15480_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_107_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10213_ input7/X _08457_/A _13282_/S vssd1 vssd1 vccd1 vccd1 _14598_/D sky130_fd_sc_hd__mux2_1
X_11193_ _11199_/A _11193_/B vssd1 vssd1 vccd1 vccd1 _11193_/Y sky130_fd_sc_hd__nor2_1
XFILLER_161_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10144_ _14529_/Q _13074_/B2 _10159_/S vssd1 vssd1 vccd1 vccd1 _14529_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_2_0_0_clk clkbuf_2_1_0_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_2_0_1_clk/A sky130_fd_sc_hd__clkbuf_8
XFILLER_121_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14952_ _15579_/CLK _14952_/D vssd1 vssd1 vccd1 vccd1 _14952_/Q sky130_fd_sc_hd__dfxtp_1
X_10075_ _14431_/Q _11861_/A1 _10092_/S vssd1 vssd1 vccd1 vccd1 _14431_/D sky130_fd_sc_hd__mux2_1
XFILLER_43_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13903_ _15677_/CLK _13903_/D vssd1 vssd1 vccd1 vccd1 _13903_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14883_ _15624_/CLK _14883_/D vssd1 vssd1 vccd1 vccd1 _14883_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_970 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_789 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13834_ _15673_/CLK _13834_/D vssd1 vssd1 vccd1 vccd1 _13834_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13765_ _14649_/CLK _13765_/D vssd1 vssd1 vccd1 vccd1 _13765_/Q sky130_fd_sc_hd__dfxtp_1
X_10977_ _11037_/A _13217_/B vssd1 vssd1 vccd1 vccd1 _11272_/B sky130_fd_sc_hd__nor2_1
XFILLER_90_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15504_ _15507_/CLK _15504_/D vssd1 vssd1 vccd1 vccd1 _15504_/Q sky130_fd_sc_hd__dfxtp_1
X_12716_ _15350_/Q _12765_/B _12715_/X _12809_/C1 vssd1 vssd1 vccd1 vccd1 _15350_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_16_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13696_ _15497_/CLK _13696_/D vssd1 vssd1 vccd1 vccd1 _13696_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_188_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15435_ _15646_/CLK _15435_/D vssd1 vssd1 vccd1 vccd1 _15435_/Q sky130_fd_sc_hd__dfxtp_1
X_12647_ _13585_/Q _12647_/B _12785_/B vssd1 vssd1 vccd1 vccd1 _12647_/X sky130_fd_sc_hd__or3_1
XFILLER_129_522 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15366_ _15646_/CLK _15366_/D vssd1 vssd1 vccd1 vccd1 _15366_/Q sky130_fd_sc_hd__dfxtp_4
X_12578_ _15138_/Q _15106_/Q _15679_/Q _13413_/Q _12430_/S _12563_/A vssd1 vssd1 vccd1
+ vccd1 _12578_/X sky130_fd_sc_hd__mux4_1
XFILLER_172_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11529_ _13214_/A _11529_/B vssd1 vssd1 vccd1 vccd1 _11532_/B sky130_fd_sc_hd__xor2_1
XFILLER_157_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14317_ _15286_/CLK _14317_/D vssd1 vssd1 vccd1 vccd1 _14317_/Q sky130_fd_sc_hd__dfxtp_1
X_15297_ _15652_/CLK _15297_/D vssd1 vssd1 vccd1 vccd1 _15297_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_171_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14248_ _15192_/CLK _14248_/D vssd1 vssd1 vccd1 vccd1 _14248_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_171_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14179_ _15665_/CLK _14179_/D vssd1 vssd1 vccd1 vccd1 _14179_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_271 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_775 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08740_ _13613_/Q _08750_/B1 _08537_/Y _14487_/Q vssd1 vssd1 vccd1 vccd1 _08740_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_112_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08671_ _13623_/Q _08750_/B1 _08535_/X _13424_/Q vssd1 vssd1 vccd1 vccd1 _08671_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_66_575 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07622_ _07620_/X _07625_/B _07629_/A vssd1 vssd1 vccd1 vccd1 _07622_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_53_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07553_ _07644_/A _07553_/B vssd1 vssd1 vccd1 vccd1 _07553_/Y sky130_fd_sc_hd__nand2_1
X_07484_ _14761_/Q _07483_/X _07500_/S vssd1 vssd1 vccd1 vccd1 _07484_/X sky130_fd_sc_hd__mux2_8
XFILLER_21_100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09223_ _09445_/C1 _09222_/X _09221_/X _09130_/A vssd1 vssd1 vccd1 vccd1 _09223_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_42_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_488 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09154_ _14530_/Q _14143_/Q _14175_/Q _14111_/Q _09407_/S _09406_/S1 vssd1 vssd1
+ vccd1 vccd1 _09154_/X sky130_fd_sc_hd__mux4_1
XFILLER_159_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08105_ input26/X input3/X input11/X input20/X _08150_/S _08151_/S vssd1 vssd1 vccd1
+ vccd1 _08105_/X sky130_fd_sc_hd__mux4_1
XFILLER_135_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09085_ _09449_/A1 _09083_/X _09084_/X _09449_/B2 _09082_/X vssd1 vssd1 vccd1 vccd1
+ _09085_/X sky130_fd_sc_hd__a221o_2
XFILLER_174_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08036_ _08036_/A _08074_/A vssd1 vssd1 vccd1 vccd1 _08037_/D sky130_fd_sc_hd__nand2_1
XFILLER_107_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09987_ _11874_/A1 _14346_/Q _09996_/S vssd1 vssd1 vccd1 vccd1 _14346_/D sky130_fd_sc_hd__mux2_1
XFILLER_130_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08938_ _13877_/Q _13123_/B _09519_/B1 _14392_/Q _08507_/A vssd1 vssd1 vccd1 vccd1
+ _08938_/X sky130_fd_sc_hd__a221o_1
XFILLER_188_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08869_ _13890_/Q _13082_/B2 _08880_/S vssd1 vssd1 vccd1 vccd1 _13890_/D sky130_fd_sc_hd__mux2_1
XTAP_3725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10900_ _13165_/B _10951_/B vssd1 vssd1 vccd1 vccd1 _10900_/Y sky130_fd_sc_hd__nand2_1
XTAP_3758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11880_ _15301_/Q _13347_/A0 _11883_/S vssd1 vssd1 vccd1 vccd1 _15301_/D sky130_fd_sc_hd__mux2_1
XTAP_3769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10831_ _14863_/Q _13805_/Q _12900_/S vssd1 vssd1 vccd1 vccd1 _14863_/D sky130_fd_sc_hd__mux2_1
XFILLER_25_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13550_ _14495_/CLK _13550_/D vssd1 vssd1 vccd1 vccd1 _13550_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_932 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10762_ _15426_/Q _14794_/Q _10765_/S vssd1 vssd1 vccd1 vccd1 _14794_/D sky130_fd_sc_hd__mux2_1
XFILLER_25_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_656 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12501_ _12494_/X _12496_/X _12498_/X _12500_/X _12501_/C1 vssd1 vssd1 vccd1 vccd1
+ _12501_/X sky130_fd_sc_hd__o221a_1
XFILLER_157_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13481_ _15399_/CLK _13481_/D vssd1 vssd1 vccd1 vccd1 _13481_/Q sky130_fd_sc_hd__dfxtp_2
X_10693_ _15034_/Q _10602_/B _10692_/X vssd1 vssd1 vccd1 vccd1 _10693_/X sky130_fd_sc_hd__a21o_1
XFILLER_139_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15220_ _15220_/CLK _15220_/D vssd1 vssd1 vccd1 vccd1 _15220_/Q sky130_fd_sc_hd__dfxtp_1
X_12432_ _12425_/X _12427_/X _12429_/X _12431_/X _06671_/A vssd1 vssd1 vccd1 vccd1
+ _12432_/X sky130_fd_sc_hd__o221a_1
XFILLER_172_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15151_ _15220_/CLK _15151_/D vssd1 vssd1 vccd1 vccd1 _15151_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_153_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12363_ _12356_/X _12358_/X _12360_/X _12362_/X _12616_/C1 vssd1 vssd1 vccd1 vccd1
+ _12363_/X sky130_fd_sc_hd__o221a_1
X_14102_ _15276_/CLK _14102_/D vssd1 vssd1 vccd1 vccd1 _14102_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_165_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11314_ _11048_/Y _11281_/Y _11313_/X _11307_/A _11311_/Y vssd1 vssd1 vccd1 vccd1
+ _11315_/B sky130_fd_sc_hd__o221a_1
X_15082_ _15679_/CLK _15082_/D vssd1 vssd1 vccd1 vccd1 _15082_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_180_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12294_ _12287_/X _12289_/X _12291_/X _12293_/X _06671_/A vssd1 vssd1 vccd1 vccd1
+ _12294_/X sky130_fd_sc_hd__o221a_1
XFILLER_107_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14033_ _14420_/CLK _14033_/D vssd1 vssd1 vccd1 vccd1 _14033_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11245_ _11283_/A _11245_/B vssd1 vssd1 vccd1 vccd1 _11245_/Y sky130_fd_sc_hd__nand2_1
X_11176_ _14980_/Q _11164_/S _11170_/X _11175_/Y vssd1 vssd1 vccd1 vccd1 _14980_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_79_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10127_ _14513_/Q _14761_/Q _10131_/S vssd1 vssd1 vccd1 vccd1 _14513_/D sky130_fd_sc_hd__mux2_1
XFILLER_121_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10058_ _14415_/Q _13344_/A0 _10059_/S vssd1 vssd1 vccd1 vccd1 _14415_/D sky130_fd_sc_hd__mux2_1
XFILLER_82_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14935_ _15558_/CLK _14935_/D vssd1 vssd1 vccd1 vccd1 _14935_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14866_ _15587_/CLK _14866_/D vssd1 vssd1 vccd1 vccd1 _14866_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13817_ _15279_/CLK _13817_/D vssd1 vssd1 vccd1 vccd1 _13817_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14797_ _15429_/CLK _14797_/D vssd1 vssd1 vccd1 vccd1 _14797_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13748_ _14868_/CLK _13748_/D vssd1 vssd1 vccd1 vccd1 _13748_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_628 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13679_ _15622_/CLK _13679_/D vssd1 vssd1 vccd1 vccd1 _13679_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_148_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15418_ _15637_/CLK _15418_/D vssd1 vssd1 vccd1 vccd1 _15418_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_163_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15349_ _15634_/CLK _15349_/D vssd1 vssd1 vccd1 vccd1 _15349_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_89_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_1087 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_1057 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09910_ _13330_/A0 _14271_/Q _09925_/S vssd1 vssd1 vccd1 vccd1 _14271_/D sky130_fd_sc_hd__mux2_1
XFILLER_99_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout606 _12470_/S vssd1 vssd1 vccd1 vccd1 _12472_/S sky130_fd_sc_hd__buf_12
X_09841_ _14205_/Q _11861_/A1 _09858_/S vssd1 vssd1 vccd1 vccd1 _14205_/D sky130_fd_sc_hd__mux2_1
XFILLER_59_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout617 _12545_/S vssd1 vssd1 vccd1 vccd1 _12430_/S sky130_fd_sc_hd__buf_12
XTAP_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout628 _14582_/Q vssd1 vssd1 vccd1 vccd1 _10507_/A1 sky130_fd_sc_hd__buf_12
XFILLER_98_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout639 fanout647/X vssd1 vssd1 vccd1 vccd1 _08084_/C1 sky130_fd_sc_hd__buf_8
XTAP_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09772_ _14139_/Q _13327_/A0 _09790_/S vssd1 vssd1 vccd1 vccd1 _14139_/D sky130_fd_sc_hd__mux2_1
XTAP_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06984_ _08237_/A _13120_/S _06983_/X vssd1 vssd1 vccd1 vccd1 _14766_/D sky130_fd_sc_hd__a21bo_1
XTAP_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08723_ _13802_/Q _12900_/S _08722_/X vssd1 vssd1 vccd1 vccd1 _13802_/D sky130_fd_sc_hd__o21a_1
XFILLER_26_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08654_ _13458_/Q _08684_/A2 _08683_/A2 _13522_/Q vssd1 vssd1 vccd1 vccd1 _08654_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_26_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07605_ _14751_/Q _07607_/A _07604_/Y _07949_/C1 vssd1 vssd1 vccd1 vccd1 _13462_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_57_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08585_ _14510_/Q _08693_/A2 _08582_/X _08583_/X _08584_/X vssd1 vssd1 vccd1 vccd1
+ _08585_/X sky130_fd_sc_hd__a2111o_1
XTAP_1619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07536_ _14727_/Q _14728_/Q _14726_/Q _14725_/Q vssd1 vssd1 vccd1 vccd1 _07658_/B
+ sky130_fd_sc_hd__and4b_1
XFILLER_169_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07467_ _13672_/Q _07499_/A2 _07499_/B1 _14700_/Q _07466_/X vssd1 vssd1 vccd1 vccd1
+ _07467_/X sky130_fd_sc_hd__a221o_1
XFILLER_22_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09206_ _13954_/Q _13696_/Q _09407_/S vssd1 vssd1 vccd1 vccd1 _09206_/X sky130_fd_sc_hd__mux2_1
XFILLER_10_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_929 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07398_ _14651_/Q _07498_/B _07498_/C vssd1 vssd1 vccd1 vccd1 _07398_/X sky130_fd_sc_hd__and3_1
XFILLER_176_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09137_ _13918_/Q _09136_/X _12481_/A vssd1 vssd1 vccd1 vccd1 _13918_/D sky130_fd_sc_hd__mux2_1
XFILLER_185_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_856 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09068_ _15281_/Q _15249_/Q _15217_/Q _15148_/Q _09073_/S _09234_/S1 vssd1 vssd1
+ vccd1 vccd1 _09068_/X sky130_fd_sc_hd__mux4_1
XFILLER_162_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08019_ _14764_/Q _08022_/B vssd1 vssd1 vccd1 vccd1 _08019_/Y sky130_fd_sc_hd__nor2_1
XFILLER_1_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11030_ _11021_/X _11029_/A _11362_/B vssd1 vssd1 vccd1 vccd1 _11031_/A sky130_fd_sc_hd__mux2_1
XFILLER_89_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12981_ _10639_/X _14874_/Q _13029_/S vssd1 vssd1 vccd1 vccd1 _12981_/X sky130_fd_sc_hd__mux2_8
XTAP_3500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1024 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14720_ _15543_/CLK _14720_/D vssd1 vssd1 vccd1 vccd1 _14720_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11932_ _14456_/Q _14424_/Q _13845_/Q _14198_/Q _12543_/S _12544_/A vssd1 vssd1 vccd1
+ vccd1 _11932_/X sky130_fd_sc_hd__mux4_1
XFILLER_17_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11863_ _15284_/Q _13330_/A0 _11878_/S vssd1 vssd1 vccd1 vccd1 _15284_/D sky130_fd_sc_hd__mux2_1
X_14651_ _15612_/CLK _14651_/D vssd1 vssd1 vccd1 vccd1 _14651_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13602_ _15378_/CLK _13602_/D vssd1 vssd1 vccd1 vccd1 _13602_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_32_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10814_ _14846_/Q _07256_/X _10868_/S vssd1 vssd1 vccd1 vccd1 _14846_/D sky130_fd_sc_hd__mux2_1
XTAP_2887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11794_ _15217_/Q _13327_/A0 _11816_/S vssd1 vssd1 vccd1 vccd1 _15217_/D sky130_fd_sc_hd__mux2_1
X_14582_ _14861_/CLK _14582_/D vssd1 vssd1 vccd1 vccd1 _14582_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_186_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_712 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10745_ _15409_/Q _14777_/Q _10759_/S vssd1 vssd1 vccd1 vccd1 _14777_/D sky130_fd_sc_hd__mux2_1
X_13533_ _14511_/CLK _13533_/D vssd1 vssd1 vccd1 vccd1 _13533_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_475 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13464_ _15385_/CLK _13464_/D vssd1 vssd1 vccd1 vccd1 _13464_/Q sky130_fd_sc_hd__dfxtp_1
X_10676_ _15573_/Q _10706_/B vssd1 vssd1 vccd1 vccd1 _10676_/X sky130_fd_sc_hd__and2_1
X_15203_ _15203_/CLK _15203_/D vssd1 vssd1 vccd1 vccd1 _15203_/Q sky130_fd_sc_hd__dfxtp_1
X_12415_ _14477_/Q _14445_/Q _13866_/Q _14219_/Q _12430_/S _12563_/A vssd1 vssd1 vccd1
+ vccd1 _12415_/X sky130_fd_sc_hd__mux4_1
XFILLER_126_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13395_ _15088_/CLK _13395_/D vssd1 vssd1 vccd1 vccd1 _13395_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_138_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12346_ _14474_/Q _14442_/Q _13863_/Q _14216_/Q _12541_/S _12540_/A vssd1 vssd1 vccd1
+ vccd1 _12346_/X sky130_fd_sc_hd__mux4_1
X_15134_ _15315_/CLK _15134_/D vssd1 vssd1 vccd1 vccd1 _15134_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_126_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15065_ _15422_/CLK _15065_/D vssd1 vssd1 vccd1 vccd1 _15065_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_5_696 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12277_ _14471_/Q _14439_/Q _13860_/Q _14213_/Q _12614_/S _12383_/A vssd1 vssd1 vccd1
+ vccd1 _12277_/X sky130_fd_sc_hd__mux4_1
XFILLER_175_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14016_ _15133_/CLK _14016_/D vssd1 vssd1 vccd1 vccd1 _14016_/Q sky130_fd_sc_hd__dfxtp_1
X_11228_ _10527_/B _15016_/Q _11237_/S vssd1 vssd1 vccd1 vccd1 _15016_/D sky130_fd_sc_hd__mux2_1
XFILLER_122_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11159_ _14975_/Q _11158_/Y _11164_/S vssd1 vssd1 vccd1 vccd1 _14975_/D sky130_fd_sc_hd__mux2_1
XFILLER_67_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14918_ _15676_/CLK _14918_/D vssd1 vssd1 vccd1 vccd1 _14918_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14849_ _15519_/CLK _14849_/D vssd1 vssd1 vccd1 vccd1 _14849_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08370_ _13726_/Q _11346_/A2 _11351_/C1 _08369_/X vssd1 vssd1 vccd1 vccd1 _13726_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_56_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07321_ _07321_/A vssd1 vssd1 vccd1 vccd1 _07321_/Y sky130_fd_sc_hd__inv_2
XFILLER_149_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07252_ _07260_/A _07260_/B _07264_/A _07264_/B vssd1 vssd1 vccd1 vccd1 _07274_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_158_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07183_ _15357_/Q _15064_/Q _07193_/S vssd1 vssd1 vccd1 vccd1 _07183_/X sky130_fd_sc_hd__mux2_8
XFILLER_145_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_173_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout403 _06825_/X vssd1 vssd1 vccd1 vccd1 _12764_/S sky130_fd_sc_hd__buf_12
XFILLER_98_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout414 _10894_/X vssd1 vssd1 vccd1 vccd1 _10951_/B sky130_fd_sc_hd__clkbuf_16
Xfanout425 _08494_/Y vssd1 vssd1 vccd1 vccd1 _09445_/A2 sky130_fd_sc_hd__buf_12
XFILLER_59_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout436 _08223_/X vssd1 vssd1 vccd1 vccd1 _11346_/A2 sky130_fd_sc_hd__buf_6
XFILLER_113_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09824_ _14190_/Q _13346_/A0 _09828_/S vssd1 vssd1 vccd1 vccd1 _14190_/D sky130_fd_sc_hd__mux2_1
XFILLER_98_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout447 _10615_/S vssd1 vssd1 vccd1 vccd1 _10610_/S sky130_fd_sc_hd__clkbuf_8
Xfanout458 _10566_/B vssd1 vssd1 vccd1 vccd1 _10344_/S sky130_fd_sc_hd__buf_12
Xfanout469 _06671_/Y vssd1 vssd1 vccd1 vccd1 _12503_/A1 sky130_fd_sc_hd__buf_12
XFILLER_150_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06967_ _06718_/Y _13494_/Q _06720_/Y _13493_/Q vssd1 vssd1 vccd1 vccd1 _06976_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_46_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09755_ _14123_/Q _11876_/A1 _09757_/S vssd1 vssd1 vccd1 vccd1 _14123_/D sky130_fd_sc_hd__mux2_1
XFILLER_67_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08706_ _15374_/Q _08748_/A2 _08736_/A2 _13419_/Q vssd1 vssd1 vccd1 vccd1 _08706_/X
+ sky130_fd_sc_hd__a22o_1
X_09686_ _14057_/Q _13341_/A0 _09695_/S vssd1 vssd1 vccd1 vccd1 _14057_/D sky130_fd_sc_hd__mux2_1
XTAP_2106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06898_ _15372_/Q _06747_/Y _15371_/Q _06749_/Y _06897_/X vssd1 vssd1 vccd1 vccd1
+ _06898_/X sky130_fd_sc_hd__a221o_1
XTAP_2128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08637_ _15384_/Q _08690_/A2 _08690_/B1 _13429_/Q vssd1 vssd1 vccd1 vccd1 _08637_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_55_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08568_ _13471_/Q _08746_/A2 _08747_/A2 _13567_/Q vssd1 vssd1 vccd1 vccd1 _08568_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_1449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07519_ _14749_/Q _13428_/Q _07529_/S vssd1 vssd1 vccd1 vccd1 _13428_/D sky130_fd_sc_hd__mux2_1
XFILLER_120_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08499_ _13131_/C _14613_/Q _14614_/Q vssd1 vssd1 vccd1 vccd1 _08536_/A sky130_fd_sc_hd__or3b_4
XFILLER_167_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10530_ _11349_/C _10530_/B _10420_/B vssd1 vssd1 vccd1 vccd1 _10548_/A sky130_fd_sc_hd__or3b_1
XFILLER_183_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10461_ _11610_/A wire360/X vssd1 vssd1 vccd1 vccd1 _10462_/B sky130_fd_sc_hd__or2_1
X_12200_ _14080_/Q _14048_/Q _12499_/S vssd1 vssd1 vccd1 vccd1 _12200_/X sky130_fd_sc_hd__mux2_1
X_13180_ _13229_/A _08313_/Y _11436_/A vssd1 vssd1 vccd1 vccd1 _13180_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_108_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10392_ _07352_/A _10457_/A2 _10391_/X vssd1 vssd1 vccd1 vccd1 _13177_/A sky130_fd_sc_hd__a21oi_4
XFILLER_163_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12131_ _14077_/Q _14045_/Q _12476_/S vssd1 vssd1 vccd1 vccd1 _12131_/X sky130_fd_sc_hd__mux2_1
XFILLER_136_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_159_1096 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12062_ _14074_/Q _14042_/Q _12453_/S vssd1 vssd1 vccd1 vccd1 _12062_/X sky130_fd_sc_hd__mux2_1
XFILLER_89_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11013_ _11013_/A _11626_/A vssd1 vssd1 vccd1 vccd1 _11013_/X sky130_fd_sc_hd__or2_1
XFILLER_2_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_467 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_426 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12964_ _07400_/X _13024_/A2 _12963_/X _12944_/A vssd1 vssd1 vccd1 vccd1 _12964_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_79_1042 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14703_ _14703_/CLK _14703_/D vssd1 vssd1 vccd1 vccd1 _14703_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11915_ _12559_/A _11915_/B vssd1 vssd1 vccd1 vccd1 _11915_/X sky130_fd_sc_hd__or2_1
XTAP_3385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12895_ _15423_/Q _15608_/Q _12927_/S vssd1 vssd1 vccd1 vccd1 _15423_/D sky130_fd_sc_hd__mux2_1
XTAP_3396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14634_ _15638_/CLK _14634_/D vssd1 vssd1 vccd1 vccd1 _14634_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11846_ _15268_/Q _11879_/A1 _11850_/S vssd1 vssd1 vccd1 vccd1 _15268_/D sky130_fd_sc_hd__mux2_1
XTAP_2684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_250 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14565_ _15664_/CLK _14565_/D vssd1 vssd1 vccd1 vccd1 _14565_/Q sky130_fd_sc_hd__dfxtp_1
X_11777_ _14897_/Q _11777_/B vssd1 vssd1 vccd1 vccd1 _11777_/Y sky130_fd_sc_hd__nand2_1
XTAP_1994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10728_ _14992_/Q _10733_/A2 _10733_/B1 _14960_/Q _10727_/X vssd1 vssd1 vccd1 vccd1
+ _10728_/X sky130_fd_sc_hd__a221o_1
X_13516_ _15374_/CLK _13516_/D vssd1 vssd1 vccd1 vccd1 _13516_/Q sky130_fd_sc_hd__dfxtp_1
X_14496_ _15378_/CLK _14496_/D vssd1 vssd1 vccd1 vccd1 _14496_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_173_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10659_ _15059_/Q _10734_/A2 _10656_/X _10658_/X vssd1 vssd1 vccd1 vccd1 _10659_/X
+ sky130_fd_sc_hd__o22a_2
XFILLER_139_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13447_ _15372_/CLK _13447_/D vssd1 vssd1 vccd1 vccd1 _13447_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_139_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13378_ _14481_/Q vssd1 vssd1 vccd1 vccd1 _14481_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_126_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_612 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15117_ _15184_/CLK _15117_/D vssd1 vssd1 vccd1 vccd1 _15117_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12329_ _12536_/A _12329_/B vssd1 vssd1 vccd1 vccd1 _12329_/X sky130_fd_sc_hd__or2_1
XFILLER_142_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15048_ _15553_/CLK _15048_/D vssd1 vssd1 vccd1 vccd1 _15048_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_141_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07870_ _13531_/Q _13530_/Q _07869_/D _13532_/Q vssd1 vssd1 vccd1 vccd1 _07870_/Y
+ sky130_fd_sc_hd__a31oi_1
XFILLER_96_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06821_ _06819_/X _06825_/B vssd1 vssd1 vccd1 vccd1 _08086_/A sky130_fd_sc_hd__and2b_1
XFILLER_28_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09540_ _13937_/Q _13139_/S _09539_/X vssd1 vssd1 vccd1 vccd1 _13937_/D sky130_fd_sc_hd__a21o_1
X_06752_ _13447_/Q vssd1 vssd1 vccd1 vccd1 _06752_/Y sky130_fd_sc_hd__inv_2
XFILLER_36_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09471_ _14481_/Q _09536_/A2 _09470_/X _13049_/A1 vssd1 vssd1 vccd1 vccd1 _09471_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_52_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06683_ _13737_/Q vssd1 vssd1 vccd1 vccd1 _06683_/Y sky130_fd_sc_hd__inv_2
XFILLER_93_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08422_ _08465_/B _08421_/Y _14614_/Q vssd1 vssd1 vccd1 vccd1 _08426_/B sky130_fd_sc_hd__o21a_4
XFILLER_51_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08353_ _07292_/B _10523_/A2 _08352_/X vssd1 vssd1 vccd1 vccd1 _08361_/B sky130_fd_sc_hd__a21oi_4
XFILLER_177_542 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07304_ _07292_/A _07292_/B _07297_/Y _07298_/X vssd1 vssd1 vccd1 vccd1 _07351_/B
+ sky130_fd_sc_hd__a22o_1
X_08284_ _11356_/C _11383_/A vssd1 vssd1 vccd1 vccd1 _11041_/B sky130_fd_sc_hd__nor2_1
XFILLER_20_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07235_ _07235_/A _07235_/B vssd1 vssd1 vccd1 vccd1 _07235_/X sky130_fd_sc_hd__and2_1
XFILLER_166_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07166_ _15340_/Q _15047_/Q _07193_/S vssd1 vssd1 vccd1 vccd1 _07166_/X sky130_fd_sc_hd__mux2_4
XFILLER_161_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07097_ _07096_/X _13611_/Q _12640_/S vssd1 vssd1 vccd1 vccd1 _07097_/X sky130_fd_sc_hd__mux2_1
XFILLER_161_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout200 _09796_/Y vssd1 vssd1 vccd1 vccd1 _09828_/S sky130_fd_sc_hd__buf_12
Xfanout211 _09596_/Y vssd1 vssd1 vccd1 vccd1 _09627_/S sky130_fd_sc_hd__buf_12
Xfanout222 _08040_/X vssd1 vssd1 vccd1 vccd1 _08066_/S sky130_fd_sc_hd__buf_12
XFILLER_8_1024 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout233 _07629_/A vssd1 vssd1 vccd1 vccd1 _07607_/A sky130_fd_sc_hd__buf_6
Xfanout244 _09831_/Y vssd1 vssd1 vccd1 vccd1 _09863_/S sky130_fd_sc_hd__buf_12
Xfanout255 _07903_/A vssd1 vssd1 vccd1 vccd1 _07816_/A sky130_fd_sc_hd__buf_6
Xfanout266 _08532_/Y vssd1 vssd1 vccd1 vccd1 _08693_/B1 sky130_fd_sc_hd__buf_12
X_09807_ _14173_/Q _13329_/A0 _09823_/S vssd1 vssd1 vccd1 vccd1 _14173_/D sky130_fd_sc_hd__mux2_1
XFILLER_75_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout277 _08511_/Y vssd1 vssd1 vccd1 vccd1 _13130_/B1 sky130_fd_sc_hd__buf_12
Xfanout288 _07492_/X vssd1 vssd1 vccd1 vccd1 _13110_/B2 sky130_fd_sc_hd__buf_4
X_07999_ _13566_/Q _08006_/D vssd1 vssd1 vccd1 vccd1 _08003_/B sky130_fd_sc_hd__nand2_1
XFILLER_46_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout299 _13098_/B2 vssd1 vssd1 vccd1 vccd1 _13342_/A0 sky130_fd_sc_hd__buf_6
XFILLER_86_286 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09738_ _14106_/Q _13326_/A0 _09757_/S vssd1 vssd1 vccd1 vccd1 _14106_/D sky130_fd_sc_hd__mux2_1
XFILLER_39_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09669_ _14040_/Q _11857_/A1 _09695_/S vssd1 vssd1 vccd1 vccd1 _14040_/D sky130_fd_sc_hd__mux2_1
XTAP_1202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11700_ _13342_/A0 _15131_/Q _11708_/S vssd1 vssd1 vccd1 vccd1 _15131_/D sky130_fd_sc_hd__mux2_1
XFILLER_131_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12680_ _15345_/Q _12679_/C _15346_/Q vssd1 vssd1 vccd1 vccd1 _12681_/B sky130_fd_sc_hd__a21oi_1
XTAP_1235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11631_ _13217_/A _11624_/A _11624_/B vssd1 vssd1 vccd1 vccd1 _11632_/B sky130_fd_sc_hd__a21boi_4
XFILLER_24_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11562_ _11563_/A _11563_/B vssd1 vssd1 vccd1 vccd1 _11564_/A sky130_fd_sc_hd__nand2_2
XFILLER_24_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14350_ _15267_/CLK _14350_/D vssd1 vssd1 vccd1 vccd1 _14350_/Q sky130_fd_sc_hd__dfxtp_1
X_13301_ _12733_/Y _15633_/Q _13309_/A vssd1 vssd1 vccd1 vccd1 _15633_/D sky130_fd_sc_hd__mux2_1
X_10513_ _10520_/A1 _13788_/Q _13756_/Q _10520_/B2 vssd1 vssd1 vccd1 vccd1 _10513_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_10_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14281_ _15300_/CLK _14281_/D vssd1 vssd1 vccd1 vccd1 _14281_/Q sky130_fd_sc_hd__dfxtp_1
X_11493_ _11493_/A _11505_/D vssd1 vssd1 vccd1 vccd1 _11493_/Y sky130_fd_sc_hd__nand2_1
X_13232_ _13233_/A _13233_/B vssd1 vssd1 vccd1 vccd1 _13232_/X sky130_fd_sc_hd__or2_1
XFILLER_137_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10444_ _08240_/A _13780_/Q _13748_/Q _08237_/A vssd1 vssd1 vccd1 vccd1 _10444_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_171_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13163_ _13217_/A _13162_/B _13219_/S _11362_/B vssd1 vssd1 vccd1 vccd1 _13163_/X
+ sky130_fd_sc_hd__o211a_1
X_10375_ _11449_/A _11476_/A vssd1 vssd1 vccd1 vccd1 _10382_/C sky130_fd_sc_hd__xor2_1
XFILLER_151_420 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12114_ _15315_/Q _13081_/A2 _12113_/X vssd1 vssd1 vccd1 vccd1 _15315_/D sky130_fd_sc_hd__a21o_1
XFILLER_2_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_5_6_0_clk clkbuf_5_7_0_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_5_6_0_clk/X sky130_fd_sc_hd__clkbuf_8
X_13094_ _13008_/X _13118_/A2 _13114_/B1 _07460_/X vssd1 vssd1 vccd1 vccd1 _13094_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_123_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12045_ _15312_/Q _13139_/S _12044_/X vssd1 vssd1 vccd1 vccd1 _15312_/D sky130_fd_sc_hd__a21o_1
XFILLER_133_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_1099 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_908 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13996_ _14405_/CLK _13996_/D vssd1 vssd1 vccd1 vccd1 _13996_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12947_ _15462_/Q _13105_/A2 _12945_/X _13025_/B1 vssd1 vssd1 vccd1 vccd1 _15462_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_34_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_492 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15666_ _15666_/CLK _15666_/D vssd1 vssd1 vccd1 vccd1 _15666_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12878_ _15406_/Q _15591_/Q _12878_/S vssd1 vssd1 vccd1 vccd1 _15406_/D sky130_fd_sc_hd__mux2_1
XTAP_2481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14617_ _15589_/CLK _14617_/D vssd1 vssd1 vccd1 vccd1 _14617_/Q sky130_fd_sc_hd__dfxtp_1
X_11829_ _15251_/Q _13072_/B2 _11849_/S vssd1 vssd1 vccd1 vccd1 _15251_/D sky130_fd_sc_hd__mux2_1
X_15597_ _15632_/CLK _15597_/D vssd1 vssd1 vccd1 vccd1 _15597_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14548_ _15672_/CLK _14548_/D vssd1 vssd1 vccd1 vccd1 _14548_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_147_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14479_ _15675_/CLK _14479_/D vssd1 vssd1 vccd1 vccd1 _14479_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_162_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07020_ _07019_/X _14739_/Q _07098_/S vssd1 vssd1 vccd1 vccd1 _13585_/D sky130_fd_sc_hd__mux2_1
XFILLER_174_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_987 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08971_ _13910_/Q _08970_/X _10868_/S vssd1 vssd1 vccd1 vccd1 _13910_/D sky130_fd_sc_hd__mux2_1
XFILLER_102_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07922_ _08012_/A2 _07921_/X input35/X vssd1 vssd1 vccd1 vccd1 _07922_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_130_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07853_ _07855_/B _07852_/X _07874_/A vssd1 vssd1 vccd1 vccd1 _07853_/X sky130_fd_sc_hd__a21bo_1
XFILLER_68_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06804_ _13730_/Q _12618_/A1 _12515_/C1 _06666_/Y _06801_/X vssd1 vssd1 vccd1 vccd1
+ _06804_/X sky130_fd_sc_hd__a221o_1
XFILLER_84_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07784_ _07779_/X _07780_/Y _07816_/A vssd1 vssd1 vccd1 vccd1 _07784_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_84_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06735_ _13454_/Q vssd1 vssd1 vccd1 vccd1 _07571_/A sky130_fd_sc_hd__inv_2
X_09523_ _09523_/A1 _09521_/X _09522_/X vssd1 vssd1 vccd1 vccd1 _09524_/C sky130_fd_sc_hd__a21o_1
XFILLER_37_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09454_ _13966_/Q _13708_/Q _09469_/S vssd1 vssd1 vccd1 vccd1 _09454_/X sky130_fd_sc_hd__mux2_1
XFILLER_80_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_857 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06666_ _13729_/Q vssd1 vssd1 vccd1 vccd1 _06666_/Y sky130_fd_sc_hd__inv_2
XPHY_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08405_ _08405_/A _08405_/B _08405_/C _08405_/D vssd1 vssd1 vccd1 vccd1 _08406_/B
+ sky130_fd_sc_hd__or4_2
XFILLER_12_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09385_ _15672_/Q _13406_/Q _09535_/S vssd1 vssd1 vccd1 vccd1 _09385_/X sky130_fd_sc_hd__mux2_1
XFILLER_101_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_28 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08336_ _11025_/A _11440_/A _10986_/B vssd1 vssd1 vccd1 vccd1 _08336_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_184_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_28 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08267_ _11088_/S _08266_/A _08261_/X vssd1 vssd1 vccd1 vccd1 _08292_/B sky130_fd_sc_hd__a21oi_4
XFILLER_137_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_140_clk clkbuf_5_29_0_clk/X vssd1 vssd1 vccd1 vccd1 _15543_/CLK sky130_fd_sc_hd__clkbuf_16
X_07218_ _07356_/B vssd1 vssd1 vccd1 vccd1 _07218_/Y sky130_fd_sc_hd__inv_2
XFILLER_137_258 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08198_ _13689_/Q _11860_/A1 _08216_/S vssd1 vssd1 vccd1 vccd1 _13689_/D sky130_fd_sc_hd__mux2_1
XFILLER_3_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07149_ _07163_/A _07149_/B vssd1 vssd1 vccd1 vccd1 _07149_/X sky130_fd_sc_hd__and2_4
XFILLER_106_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10160_ _14545_/Q _13346_/A0 _10164_/S vssd1 vssd1 vccd1 vccd1 _14545_/D sky130_fd_sc_hd__mux2_1
XFILLER_106_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10091_ _14447_/Q _11877_/A1 _10092_/S vssd1 vssd1 vccd1 vccd1 _14447_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13850_ _15284_/CLK _13850_/D vssd1 vssd1 vccd1 vccd1 _13850_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12801_ _13439_/Q _12647_/B _08030_/Y _13606_/Q _12743_/A vssd1 vssd1 vccd1 vccd1
+ _12801_/X sky130_fd_sc_hd__a221o_2
XFILLER_142_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13781_ _15393_/CLK _13781_/D vssd1 vssd1 vccd1 vccd1 _13781_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_62_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_1012 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10993_ _11330_/A _10991_/Y _10992_/X vssd1 vssd1 vccd1 vccd1 _10993_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_43_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15520_ _15520_/CLK _15520_/D vssd1 vssd1 vccd1 vccd1 _15520_/Q sky130_fd_sc_hd__dfxtp_1
X_12732_ _15353_/Q _12732_/B vssd1 vssd1 vccd1 vccd1 _12733_/B sky130_fd_sc_hd__nor2_1
XTAP_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15451_ _15637_/CLK _15451_/D vssd1 vssd1 vccd1 vccd1 _15451_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12663_ _12743_/A _12663_/B vssd1 vssd1 vccd1 vccd1 _12663_/X sky130_fd_sc_hd__or2_1
XTAP_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14402_ _15233_/CLK _14402_/D vssd1 vssd1 vccd1 vccd1 _14402_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_187_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11614_ _11613_/Y _15070_/Q _11614_/S vssd1 vssd1 vccd1 vccd1 _15070_/D sky130_fd_sc_hd__mux2_1
X_15382_ _15383_/CLK _15382_/D vssd1 vssd1 vccd1 vccd1 _15382_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_184_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12594_ _12577_/X _12578_/X _12594_/S vssd1 vssd1 vccd1 vccd1 _12594_/X sky130_fd_sc_hd__mux2_1
XFILLER_129_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14333_ _15181_/CLK _14333_/D vssd1 vssd1 vccd1 vccd1 _14333_/Q sky130_fd_sc_hd__dfxtp_1
X_11545_ _11523_/Y _11546_/C _11543_/Y vssd1 vssd1 vccd1 vccd1 _11545_/X sky130_fd_sc_hd__a21o_1
XFILLER_11_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_522 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_131_clk clkbuf_5_28_0_clk/X vssd1 vssd1 vccd1 vccd1 _13798_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_184_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_183_364 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11476_ _11476_/A _11476_/B _11476_/C _11476_/D vssd1 vssd1 vccd1 vccd1 _11496_/C
+ sky130_fd_sc_hd__and4_1
XFILLER_156_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14264_ _15273_/CLK _14264_/D vssd1 vssd1 vccd1 vccd1 _14264_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_143_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13215_ _13233_/A _13215_/B vssd1 vssd1 vccd1 vccd1 _13215_/Y sky130_fd_sc_hd__xnor2_1
X_10427_ _11349_/C _11632_/A vssd1 vssd1 vccd1 vccd1 _10429_/A sky130_fd_sc_hd__or2_1
X_14195_ _14861_/CLK _14195_/D vssd1 vssd1 vccd1 vccd1 _14195_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_140_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10358_ _07284_/A _10360_/B _10357_/X vssd1 vssd1 vccd1 vccd1 _11475_/A sky130_fd_sc_hd__a21o_4
XFILLER_83_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13146_ _09382_/A _15544_/Q _13154_/S vssd1 vssd1 vccd1 vccd1 _15544_/D sky130_fd_sc_hd__mux2_1
XFILLER_151_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13077_ _15506_/Q _13081_/A2 _13105_/B1 _13076_/X vssd1 vssd1 vccd1 vccd1 _15506_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_183_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10289_ _14674_/Q _14827_/Q _10695_/S vssd1 vssd1 vccd1 vccd1 _14674_/D sky130_fd_sc_hd__mux2_1
XFILLER_39_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12028_ _14362_/Q _15178_/Q _13817_/Q _14556_/Q _12591_/S _12590_/A vssd1 vssd1 vccd1
+ vccd1 _12028_/X sky130_fd_sc_hd__mux4_1
XFILLER_38_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_198_clk clkbuf_5_17_0_clk/X vssd1 vssd1 vccd1 vccd1 _15654_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_66_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13979_ _14083_/CLK _13979_/D vssd1 vssd1 vccd1 vccd1 _13979_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_687 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15649_ _15649_/CLK _15649_/D vssd1 vssd1 vccd1 vccd1 _15649_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09170_ _14080_/Q _09445_/A2 _09522_/B1 _14048_/Q _09435_/A vssd1 vssd1 vccd1 vccd1
+ _09170_/X sky130_fd_sc_hd__a221o_1
XFILLER_187_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08121_ _08121_/A _08121_/B vssd1 vssd1 vccd1 vccd1 _08121_/X sky130_fd_sc_hd__and2_4
XFILLER_159_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_122_clk clkbuf_5_30_0_clk/X vssd1 vssd1 vccd1 vccd1 _13627_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_147_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08052_ _14745_/Q _13623_/Q _08072_/S vssd1 vssd1 vccd1 vccd1 _13623_/D sky130_fd_sc_hd__mux2_1
XFILLER_162_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07003_ _14718_/Q _07783_/A _08027_/A vssd1 vssd1 vccd1 vccd1 _12839_/B sky130_fd_sc_hd__or3_2
XFILLER_115_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_935 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08954_ _09445_/C1 _08953_/X _08952_/X _09130_/A vssd1 vssd1 vccd1 vccd1 _08954_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_57_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07905_ _13541_/Q _07913_/D vssd1 vssd1 vccd1 vccd1 _07910_/B sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_189_clk clkbuf_5_21_0_clk/X vssd1 vssd1 vccd1 vccd1 _15293_/CLK sky130_fd_sc_hd__clkbuf_16
X_08885_ _13906_/Q _13350_/A0 _08885_/S vssd1 vssd1 vccd1 vccd1 _13906_/D sky130_fd_sc_hd__mux2_1
XFILLER_111_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07836_ _13523_/Q _13522_/Q _13521_/Q _07836_/D vssd1 vssd1 vccd1 vccd1 _07847_/D
+ sky130_fd_sc_hd__and4_2
XTAP_3918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07767_ _14762_/Q _07777_/A _07766_/Y _08012_/C1 vssd1 vssd1 vccd1 vccd1 _13505_/D
+ sky130_fd_sc_hd__o211a_1
X_09506_ _08494_/B _09504_/X _09505_/X vssd1 vssd1 vccd1 vccd1 _09510_/B sky130_fd_sc_hd__a21o_1
X_06718_ _14503_/Q vssd1 vssd1 vccd1 vccd1 _06718_/Y sky130_fd_sc_hd__inv_2
X_07698_ _07713_/A _07698_/B vssd1 vssd1 vccd1 vccd1 _07698_/Y sky130_fd_sc_hd__nand2_1
XFILLER_72_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09437_ _09437_/A1 _09436_/X _09435_/X _14606_/Q vssd1 vssd1 vccd1 vccd1 _09437_/X
+ sky130_fd_sc_hd__o211a_1
XPHY_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_668 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09368_ _13929_/Q _13093_/A2 _09367_/X vssd1 vssd1 vccd1 vccd1 _13929_/D sky130_fd_sc_hd__a21o_1
XFILLER_36_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08319_ _08281_/X _08318_/X _11047_/B vssd1 vssd1 vccd1 vccd1 _08319_/X sky130_fd_sc_hd__mux2_2
Xclkbuf_leaf_113_clk _15447_/CLK vssd1 vssd1 vccd1 vccd1 _15381_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_166_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09299_ _14537_/Q _14150_/Q _14182_/Q _14118_/Q _09484_/S _08519_/A vssd1 vssd1 vccd1
+ vccd1 _09299_/X sky130_fd_sc_hd__mux4_1
XFILLER_123_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_60 _07169_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_71 _07145_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_82 _07119_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11330_ _11330_/A _11330_/B vssd1 vssd1 vccd1 vccd1 _11330_/Y sky130_fd_sc_hd__nand2_1
XANTENNA_93 _08507_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11261_ _08338_/X _11260_/X _11329_/A vssd1 vssd1 vccd1 vccd1 _11262_/B sky130_fd_sc_hd__mux2_1
XFILLER_21_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13000_ _07448_/X _13039_/A2 _12999_/X _12944_/A vssd1 vssd1 vccd1 vccd1 _13000_/X
+ sky130_fd_sc_hd__a22o_1
X_10212_ input6/X _14597_/Q _13284_/S vssd1 vssd1 vccd1 vccd1 _14597_/D sky130_fd_sc_hd__mux2_1
X_11192_ _14988_/Q _11164_/S _11170_/X _11191_/Y vssd1 vssd1 vccd1 vccd1 _14988_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_137_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_795 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10143_ _14528_/Q _13329_/A0 _10159_/S vssd1 vssd1 vccd1 vccd1 _14528_/D sky130_fd_sc_hd__mux2_1
XFILLER_122_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10074_ _14430_/Q _11860_/A1 _10092_/S vssd1 vssd1 vccd1 vccd1 _14430_/D sky130_fd_sc_hd__mux2_1
XFILLER_94_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14951_ _15581_/CLK _14951_/D vssd1 vssd1 vccd1 vccd1 _14951_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13902_ _15161_/CLK _13902_/D vssd1 vssd1 vccd1 vccd1 _13902_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_532 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1088 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14882_ _15624_/CLK _14882_/D vssd1 vssd1 vccd1 vccd1 _14882_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13833_ _14572_/CLK _13833_/D vssd1 vssd1 vccd1 vccd1 _13833_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_226 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13764_ _14888_/CLK _13764_/D vssd1 vssd1 vccd1 vccd1 _13764_/Q sky130_fd_sc_hd__dfxtp_1
X_10976_ _11037_/A _13220_/B vssd1 vssd1 vccd1 vccd1 _11305_/C sky130_fd_sc_hd__nand2_1
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15503_ _15508_/CLK _15503_/D vssd1 vssd1 vccd1 vccd1 _15503_/Q sky130_fd_sc_hd__dfxtp_1
X_12715_ _12737_/A _12715_/B vssd1 vssd1 vccd1 vccd1 _12715_/X sky130_fd_sc_hd__or2_1
XFILLER_188_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13695_ _15658_/CLK _13695_/D vssd1 vssd1 vccd1 vccd1 _13695_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15434_ _15434_/CLK _15434_/D vssd1 vssd1 vccd1 vccd1 _15434_/Q sky130_fd_sc_hd__dfxtp_1
X_12646_ _15048_/Q _12645_/Y _12834_/B vssd1 vssd1 vccd1 vccd1 _12646_/X sky130_fd_sc_hd__mux2_1
XFILLER_15_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_104_clk clkbuf_5_26_0_clk/X vssd1 vssd1 vccd1 vccd1 _15438_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_12_882 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15365_ _15645_/CLK _15365_/D vssd1 vssd1 vccd1 vccd1 _15365_/Q sky130_fd_sc_hd__dfxtp_2
X_12577_ _14548_/Q _14161_/Q _14193_/Q _14129_/Q _12430_/S _12563_/A vssd1 vssd1 vccd1
+ vccd1 _12577_/X sky130_fd_sc_hd__mux4_1
XFILLER_50_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14316_ _15510_/CLK _14316_/D vssd1 vssd1 vccd1 vccd1 _14316_/Q sky130_fd_sc_hd__dfxtp_1
X_11528_ _11536_/A _11536_/B _11536_/C _11537_/A _13236_/A vssd1 vssd1 vccd1 vccd1
+ _11529_/B sky130_fd_sc_hd__a41o_1
XFILLER_117_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15296_ _15328_/CLK _15296_/D vssd1 vssd1 vccd1 vccd1 _15296_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_156_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14247_ _15292_/CLK _14247_/D vssd1 vssd1 vccd1 vccd1 _14247_/Q sky130_fd_sc_hd__dfxtp_1
X_11459_ _11440_/Y _11459_/B vssd1 vssd1 vccd1 vccd1 _11460_/C sky130_fd_sc_hd__and2b_1
XFILLER_171_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_378 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14178_ _15315_/CLK _14178_/D vssd1 vssd1 vccd1 vccd1 _14178_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_140_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_283 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13129_ _13129_/A _13129_/B vssd1 vssd1 vccd1 vccd1 _13129_/Y sky130_fd_sc_hd__nor2_1
XFILLER_30_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_990 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08670_ _13520_/Q _08683_/A2 _08691_/B1 _13488_/Q _08669_/X vssd1 vssd1 vccd1 vccd1
+ _08670_/X sky130_fd_sc_hd__a221o_2
XFILLER_66_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07621_ _07621_/A _07621_/B vssd1 vssd1 vccd1 vccd1 _07625_/B sky130_fd_sc_hd__nor2_1
XFILLER_66_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07552_ _13449_/Q _07559_/D vssd1 vssd1 vccd1 vccd1 _07553_/B sky130_fd_sc_hd__xnor2_1
XFILLER_179_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07483_ _13676_/Q _07483_/A2 _07483_/B1 _14704_/Q _07482_/X vssd1 vssd1 vccd1 vccd1
+ _07483_/X sky130_fd_sc_hd__a221o_1
XFILLER_179_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09222_ _15289_/Q _15257_/Q _15225_/Q _15156_/Q _09225_/S0 _09225_/S1 vssd1 vssd1
+ vccd1 vccd1 _09222_/X sky130_fd_sc_hd__mux4_1
XFILLER_22_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09153_ _15120_/Q _15088_/Q _15661_/Q _13395_/Q _09407_/S _09406_/S1 vssd1 vssd1
+ vccd1 vccd1 _09153_/X sky130_fd_sc_hd__mux4_1
XFILLER_148_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08104_ input11/X input20/X _08145_/S vssd1 vssd1 vccd1 vccd1 _08161_/B sky130_fd_sc_hd__mux2_1
XFILLER_148_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09084_ _14237_/Q _14269_/Q _14301_/Q _14333_/Q _09190_/S _09429_/S1 vssd1 vssd1
+ vccd1 vccd1 _09084_/X sky130_fd_sc_hd__mux4_1
XFILLER_135_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08035_ _13576_/Q _14737_/Q _08039_/S vssd1 vssd1 vccd1 vccd1 _13576_/D sky130_fd_sc_hd__mux2_1
XFILLER_162_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09986_ _11873_/A1 _14345_/Q _09996_/S vssd1 vssd1 vccd1 vccd1 _14345_/D sky130_fd_sc_hd__mux2_1
XFILLER_104_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08937_ _13941_/Q _13683_/Q _09484_/S vssd1 vssd1 vccd1 vccd1 _08937_/X sky130_fd_sc_hd__mux2_1
XFILLER_130_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08868_ _13889_/Q _13333_/A0 _08880_/S vssd1 vssd1 vccd1 vccd1 _13889_/D sky130_fd_sc_hd__mux2_1
XTAP_3726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07819_ _07830_/A _07819_/B vssd1 vssd1 vccd1 vccd1 _07819_/Y sky130_fd_sc_hd__nand2_1
XTAP_3759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08799_ _13333_/A0 _13825_/Q _08811_/S vssd1 vssd1 vccd1 vccd1 _13825_/D sky130_fd_sc_hd__mux2_1
X_10830_ _13806_/Q _14862_/Q _10834_/S vssd1 vssd1 vccd1 vccd1 _14862_/D sky130_fd_sc_hd__mux2_1
XFILLER_53_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10761_ _15425_/Q _14793_/Q _10765_/S vssd1 vssd1 vccd1 vccd1 _14793_/D sky130_fd_sc_hd__mux2_1
XFILLER_41_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12500_ _12500_/A1 _12499_/X _12500_/B1 vssd1 vssd1 vccd1 vccd1 _12500_/X sky130_fd_sc_hd__a21o_1
XFILLER_13_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13480_ _15543_/CLK _13480_/D vssd1 vssd1 vccd1 vccd1 _13480_/Q sky130_fd_sc_hd__dfxtp_2
X_10692_ _15576_/Q _10731_/B _10733_/B1 _14953_/Q vssd1 vssd1 vccd1 vccd1 _10692_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_41_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12431_ _12615_/A1 _12430_/X _06670_/A vssd1 vssd1 vccd1 vccd1 _12431_/X sky130_fd_sc_hd__a21o_1
XFILLER_8_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15150_ _15662_/CLK _15150_/D vssd1 vssd1 vccd1 vccd1 _15150_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_148_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12362_ _12592_/A1 _12361_/X _12615_/B1 vssd1 vssd1 vccd1 vccd1 _12362_/X sky130_fd_sc_hd__a21o_1
XFILLER_166_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14101_ _15651_/CLK _14101_/D vssd1 vssd1 vccd1 vccd1 _14101_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_148_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11313_ _11294_/Y _11312_/Y _11349_/A vssd1 vssd1 vccd1 vccd1 _11313_/X sky130_fd_sc_hd__mux2_1
XFILLER_153_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15081_ _15081_/CLK _15081_/D vssd1 vssd1 vccd1 vccd1 _15081_/Q sky130_fd_sc_hd__dfxtp_1
X_12293_ _12592_/A1 _12292_/X _06670_/A vssd1 vssd1 vccd1 vccd1 _12293_/X sky130_fd_sc_hd__a21o_1
XFILLER_180_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11244_ _08357_/A _11243_/X _11297_/S vssd1 vssd1 vccd1 vccd1 _11245_/B sky130_fd_sc_hd__mux2_1
X_14032_ _15226_/CLK _14032_/D vssd1 vssd1 vccd1 vccd1 _14032_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_106_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11175_ _11199_/A _11175_/B vssd1 vssd1 vccd1 vccd1 _11175_/Y sky130_fd_sc_hd__nor2_1
XFILLER_121_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10126_ _14512_/Q _14760_/Q _10131_/S vssd1 vssd1 vccd1 vccd1 _14512_/D sky130_fd_sc_hd__mux2_1
XFILLER_132_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10057_ _14414_/Q _13343_/A0 _10059_/S vssd1 vssd1 vccd1 vccd1 _14414_/D sky130_fd_sc_hd__mux2_1
X_14934_ _15558_/CLK _14934_/D vssd1 vssd1 vccd1 vccd1 _14934_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14865_ _15588_/CLK _14865_/D vssd1 vssd1 vccd1 vccd1 _14865_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_169_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13816_ _15142_/CLK _13816_/D vssd1 vssd1 vccd1 vccd1 _13816_/Q sky130_fd_sc_hd__dfxtp_1
X_14796_ _14868_/CLK _14796_/D vssd1 vssd1 vccd1 vccd1 _14796_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_451 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_996 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13747_ _14649_/CLK _13747_/D vssd1 vssd1 vccd1 vccd1 _13747_/Q sky130_fd_sc_hd__dfxtp_1
X_10959_ _11259_/S _10958_/Y _10955_/Y vssd1 vssd1 vccd1 vccd1 _10959_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_43_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13678_ _14892_/CLK _13678_/D vssd1 vssd1 vccd1 vccd1 _13678_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_148_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15417_ _15453_/CLK _15417_/D vssd1 vssd1 vccd1 vccd1 _15417_/Q sky130_fd_sc_hd__dfxtp_2
X_12629_ _15339_/Q _15338_/Q vssd1 vssd1 vccd1 vccd1 _12629_/X sky130_fd_sc_hd__xor2_1
XFILLER_157_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_1060 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15348_ _15630_/CLK _15348_/D vssd1 vssd1 vccd1 vccd1 _15348_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_106_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15279_ _15279_/CLK _15279_/D vssd1 vssd1 vccd1 vccd1 _15279_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_171_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_1099 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_1069 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout607 _12079_/S vssd1 vssd1 vccd1 vccd1 _12269_/S sky130_fd_sc_hd__buf_12
X_09840_ _14204_/Q _11860_/A1 _09858_/S vssd1 vssd1 vccd1 vccd1 _14204_/D sky130_fd_sc_hd__mux2_1
XTAP_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout618 _12545_/S vssd1 vssd1 vccd1 vccd1 _12568_/S sky130_fd_sc_hd__buf_6
XFILLER_140_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout629 _10515_/B2 vssd1 vssd1 vccd1 vccd1 _08244_/B sky130_fd_sc_hd__buf_8
XFILLER_99_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09771_ _14138_/Q _13326_/A0 _09790_/S vssd1 vssd1 vccd1 vccd1 _14138_/D sky130_fd_sc_hd__mux2_1
XTAP_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06983_ _14596_/Q _08477_/C _06808_/X _13120_/S vssd1 vssd1 vccd1 vccd1 _06983_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_101_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08722_ _08722_/A _08722_/B _08722_/C vssd1 vssd1 vccd1 vccd1 _08722_/X sky130_fd_sc_hd__or3_4
XFILLER_113_1031 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_1075 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08653_ _13792_/Q _12917_/S _08652_/X vssd1 vssd1 vccd1 vccd1 _13792_/D sky130_fd_sc_hd__o21a_1
XFILLER_39_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07604_ _07602_/Y _07610_/C _07607_/A vssd1 vssd1 vccd1 vccd1 _07604_/Y sky130_fd_sc_hd__o21ai_1
XTAP_1609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08584_ _13604_/Q _08691_/A2 _08747_/A2 _13565_/Q vssd1 vssd1 vccd1 vccd1 _08584_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_42_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07535_ _14765_/Q _13444_/Q _07535_/S vssd1 vssd1 vccd1 vccd1 _13444_/D sky130_fd_sc_hd__mux2_1
XFILLER_22_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07466_ _14668_/Q _07474_/B _07482_/C vssd1 vssd1 vccd1 vccd1 _07466_/X sky130_fd_sc_hd__and3_1
XFILLER_179_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09205_ _09421_/A1 _09203_/X _09204_/X _09419_/A2 _14607_/Q vssd1 vssd1 vccd1 vccd1
+ _09205_/X sky130_fd_sc_hd__a221o_1
XFILLER_50_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07397_ _13324_/A0 _13388_/Q _07501_/S vssd1 vssd1 vccd1 vccd1 _13388_/D sky130_fd_sc_hd__mux2_1
XFILLER_10_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09136_ _09120_/X _09123_/X _09130_/X _09135_/X vssd1 vssd1 vccd1 vccd1 _09136_/X
+ sky130_fd_sc_hd__o22a_2
XFILLER_33_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_1024 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09067_ _09421_/A1 _09063_/X _09066_/X _09062_/X vssd1 vssd1 vccd1 vccd1 _09077_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_123_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08018_ _13571_/Q _08018_/B vssd1 vssd1 vccd1 vccd1 _08018_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_151_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09969_ _11681_/A0 _14328_/Q _09991_/S vssd1 vssd1 vccd1 vccd1 _14328_/D sky130_fd_sc_hd__mux2_1
XFILLER_134_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12980_ _15473_/Q _13081_/A2 _13025_/B1 _12979_/X vssd1 vssd1 vccd1 vccd1 _15473_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_182_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11931_ _14230_/Q _14262_/Q _14294_/Q _14326_/Q _12543_/S _12544_/A vssd1 vssd1 vccd1
+ vccd1 _11931_/X sky130_fd_sc_hd__mux4_1
XTAP_3545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14650_ _15620_/CLK _14650_/D vssd1 vssd1 vccd1 vccd1 _14650_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11862_ _15283_/Q _13329_/A0 _11878_/S vssd1 vssd1 vccd1 vccd1 _15283_/D sky130_fd_sc_hd__mux2_1
XTAP_2844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13601_ _15637_/CLK _13601_/D vssd1 vssd1 vccd1 vccd1 _13601_/Q sky130_fd_sc_hd__dfxtp_2
X_10813_ _14845_/Q _10360_/A _12900_/S vssd1 vssd1 vccd1 vccd1 _14845_/D sky130_fd_sc_hd__mux2_1
XTAP_2877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14581_ _15680_/CLK _14581_/D vssd1 vssd1 vccd1 vccd1 _14581_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11793_ _15216_/Q _12967_/A1 _11816_/S vssd1 vssd1 vccd1 vccd1 _15216_/D sky130_fd_sc_hd__mux2_1
XTAP_2899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13532_ _13565_/CLK _13532_/D vssd1 vssd1 vccd1 vccd1 _13532_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_186_724 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10744_ _15408_/Q _14776_/Q _10759_/S vssd1 vssd1 vccd1 vccd1 _14776_/D sky130_fd_sc_hd__mux2_1
XFILLER_9_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_487 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13463_ _15385_/CLK _13463_/D vssd1 vssd1 vccd1 vccd1 _13463_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_9_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_95 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10675_ _14753_/Q _10674_/X _10715_/S vssd1 vssd1 vccd1 vccd1 _14753_/D sky130_fd_sc_hd__mux2_1
X_15202_ _15202_/CLK _15202_/D vssd1 vssd1 vccd1 vccd1 _15202_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_982 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12414_ _14251_/Q _14283_/Q _14315_/Q _14347_/Q _12430_/S _12563_/A vssd1 vssd1 vccd1
+ vccd1 _12414_/X sky130_fd_sc_hd__mux4_1
X_13394_ _15660_/CLK _13394_/D vssd1 vssd1 vccd1 vccd1 _13394_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_138_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15133_ _15133_/CLK _15133_/D vssd1 vssd1 vccd1 vccd1 _15133_/Q sky130_fd_sc_hd__dfxtp_1
X_12345_ _14248_/Q _14280_/Q _14312_/Q _14344_/Q _12541_/S _12540_/A vssd1 vssd1 vccd1
+ vccd1 _12345_/X sky130_fd_sc_hd__mux4_1
XFILLER_153_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15064_ _15422_/CLK _15064_/D vssd1 vssd1 vccd1 vccd1 _15064_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_142_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12276_ _14245_/Q _14277_/Q _14309_/Q _14341_/Q _12614_/S _12383_/A vssd1 vssd1 vccd1
+ vccd1 _12276_/X sky130_fd_sc_hd__mux4_1
XFILLER_153_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14015_ _15510_/CLK _14015_/D vssd1 vssd1 vccd1 vccd1 _14015_/Q sky130_fd_sc_hd__dfxtp_1
X_11227_ _10527_/C _15015_/Q _11237_/S vssd1 vssd1 vccd1 vccd1 _15015_/D sky130_fd_sc_hd__mux2_1
XFILLER_49_1083 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11158_ _11199_/A _11197_/B _11157_/X vssd1 vssd1 vccd1 vccd1 _11158_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_68_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10109_ _14495_/Q _14743_/Q _10124_/S vssd1 vssd1 vccd1 vccd1 _14495_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11089_ _11307_/A _11087_/X _11088_/X _11048_/Y _11414_/A vssd1 vssd1 vccd1 vccd1
+ _11089_/X sky130_fd_sc_hd__o221a_1
XFILLER_48_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14917_ _15548_/CLK _14917_/D vssd1 vssd1 vccd1 vccd1 _14917_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14848_ _15501_/CLK _14848_/D vssd1 vssd1 vccd1 vccd1 _14848_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14779_ _15596_/CLK _14779_/D vssd1 vssd1 vccd1 vccd1 _14779_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07320_ _15311_/Q _15467_/Q _07335_/S vssd1 vssd1 vccd1 vccd1 _07321_/A sky130_fd_sc_hd__mux2_4
XFILLER_177_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07251_ _07251_/A vssd1 vssd1 vccd1 vccd1 _07264_/B sky130_fd_sc_hd__inv_2
XFILLER_104_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07182_ _15356_/Q _15063_/Q _07188_/S vssd1 vssd1 vccd1 vccd1 _07182_/X sky130_fd_sc_hd__mux2_8
XFILLER_117_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout404 _13241_/A2 vssd1 vssd1 vccd1 vccd1 _13214_/B sky130_fd_sc_hd__buf_6
XFILLER_113_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout415 _10948_/B vssd1 vssd1 vccd1 vccd1 _10944_/B sky130_fd_sc_hd__buf_8
Xfanout426 _13123_/B vssd1 vssd1 vccd1 vccd1 _09522_/A2 sky130_fd_sc_hd__buf_12
XFILLER_99_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09823_ _14189_/Q _13345_/A0 _09823_/S vssd1 vssd1 vccd1 vccd1 _14189_/D sky130_fd_sc_hd__mux2_1
XFILLER_99_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout448 _10244_/S vssd1 vssd1 vccd1 vccd1 _10615_/S sky130_fd_sc_hd__buf_12
Xfanout459 _06769_/Y vssd1 vssd1 vccd1 vccd1 _13217_/A sky130_fd_sc_hd__buf_12
XFILLER_150_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09754_ _14122_/Q _13342_/A0 _09762_/S vssd1 vssd1 vccd1 vccd1 _14122_/D sky130_fd_sc_hd__mux2_1
X_06966_ _14505_/Q _06715_/Y _06716_/Y _13495_/Q vssd1 vssd1 vccd1 vccd1 _06977_/A
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_27_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08705_ _13586_/Q _08749_/A2 _08747_/A2 _13547_/Q _08704_/X vssd1 vssd1 vccd1 vccd1
+ _08709_/B sky130_fd_sc_hd__a221o_1
X_09685_ _14056_/Q _13340_/A0 _09695_/S vssd1 vssd1 vccd1 vccd1 _14056_/D sky130_fd_sc_hd__mux2_1
XTAP_2107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06897_ _15371_/Q _06749_/Y _15370_/Q _06752_/Y _06896_/X vssd1 vssd1 vccd1 vccd1
+ _06897_/X sky130_fd_sc_hd__o221a_1
XFILLER_55_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_93_clk clkbuf_5_24_0_clk/X vssd1 vssd1 vccd1 vccd1 _15620_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_2129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08636_ _13557_/Q _08685_/A2 _08691_/B1 _13493_/Q vssd1 vssd1 vccd1 vccd1 _08636_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_1406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08567_ _13779_/Q _08573_/S _08566_/X vssd1 vssd1 vccd1 vccd1 _13779_/D sky130_fd_sc_hd__o21a_1
XFILLER_70_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07518_ _14748_/Q _13427_/Q _07529_/S vssd1 vssd1 vccd1 vccd1 _13427_/D sky130_fd_sc_hd__mux2_1
XFILLER_168_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08498_ _14612_/Q _14611_/Q vssd1 vssd1 vccd1 vccd1 _13131_/C sky130_fd_sc_hd__nand2_1
XFILLER_23_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07449_ _13337_/A0 _13401_/Q _07501_/S vssd1 vssd1 vccd1 vccd1 _13401_/D sky130_fd_sc_hd__mux2_1
XFILLER_167_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_929 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10460_ _11610_/A wire360/X vssd1 vssd1 vccd1 vccd1 _10462_/A sky130_fd_sc_hd__nand2_1
X_09119_ _09221_/A _09119_/B vssd1 vssd1 vccd1 vccd1 _09119_/X sky130_fd_sc_hd__or2_1
X_10391_ _08240_/A _13799_/Q _13767_/Q _08237_/A vssd1 vssd1 vccd1 vccd1 _10391_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_109_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12130_ _12498_/A _12130_/B vssd1 vssd1 vccd1 vccd1 _12130_/X sky130_fd_sc_hd__and2_1
XFILLER_163_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12061_ _12061_/A _12061_/B vssd1 vssd1 vccd1 vccd1 _12061_/X sky130_fd_sc_hd__and2_1
XFILLER_89_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11012_ _13217_/A _11013_/A _11349_/A vssd1 vssd1 vccd1 vccd1 _11357_/B sky130_fd_sc_hd__a21o_1
XTAP_4010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12963_ _10609_/X _14868_/Q _13038_/S vssd1 vssd1 vccd1 vccd1 _12963_/X sky130_fd_sc_hd__mux2_4
XTAP_4076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_490 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_84_clk clkbuf_5_12_0_clk/X vssd1 vssd1 vccd1 vccd1 _14888_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_4098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14702_ _15607_/CLK _14702_/D vssd1 vssd1 vccd1 vccd1 _14702_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11914_ _15274_/Q _15242_/Q _15210_/Q _15141_/Q _12522_/S _12521_/A vssd1 vssd1 vccd1
+ vccd1 _11915_/B sky130_fd_sc_hd__mux4_1
XFILLER_79_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12894_ _15422_/Q _15607_/Q _12927_/S vssd1 vssd1 vccd1 vccd1 _15422_/D sky130_fd_sc_hd__mux2_1
XTAP_3375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_1076 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14633_ _15636_/CLK _14633_/D vssd1 vssd1 vccd1 vccd1 _14633_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11845_ _15267_/Q _13104_/B2 _11849_/S vssd1 vssd1 vccd1 vccd1 _15267_/D sky130_fd_sc_hd__mux2_1
XTAP_2674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14564_ _15287_/CLK _14564_/D vssd1 vssd1 vccd1 vccd1 _14564_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11776_ _15207_/Q _11777_/B vssd1 vssd1 vccd1 vccd1 _11776_/X sky130_fd_sc_hd__or2_1
XFILLER_9_200 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13515_ _15374_/CLK _13515_/D vssd1 vssd1 vccd1 vccd1 _13515_/Q sky130_fd_sc_hd__dfxtp_1
X_10727_ _15024_/Q _10569_/B _10602_/B _15041_/Q _10732_/C1 vssd1 vssd1 vccd1 vccd1
+ _10727_/X sky130_fd_sc_hd__a221o_1
X_14495_ _14495_/CLK _14495_/D vssd1 vssd1 vccd1 vccd1 _14495_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_186_576 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13446_ _15543_/CLK _13446_/D vssd1 vssd1 vccd1 vccd1 _13446_/Q sky130_fd_sc_hd__dfxtp_2
X_10658_ _14978_/Q _10733_/A2 _10722_/B1 _14946_/Q _10657_/X vssd1 vssd1 vccd1 vccd1
+ _10658_/X sky130_fd_sc_hd__a221o_1
XFILLER_70_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_120 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13377_ _14480_/Q vssd1 vssd1 vccd1 vccd1 _14480_/D sky130_fd_sc_hd__clkbuf_2
X_10589_ _15045_/Q _10734_/A2 _10586_/X _10588_/X vssd1 vssd1 vccd1 vccd1 _10589_/X
+ sky130_fd_sc_hd__o22a_4
X_15116_ _15244_/CLK _15116_/D vssd1 vssd1 vccd1 vccd1 _15116_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_126_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_624 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12328_ _15292_/Q _15260_/Q _15228_/Q _15159_/Q _12543_/S _12544_/A vssd1 vssd1 vccd1
+ vccd1 _12329_/B sky130_fd_sc_hd__mux4_1
XFILLER_47_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15047_ _15553_/CLK _15047_/D vssd1 vssd1 vccd1 vccd1 _15047_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_114_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12259_ _15289_/Q _15257_/Q _15225_/Q _15156_/Q _11993_/S _11992_/A vssd1 vssd1 vccd1
+ vccd1 _12260_/B sky130_fd_sc_hd__mux4_1
XFILLER_141_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06820_ _13576_/Q _13574_/Q _13577_/Q vssd1 vssd1 vccd1 vccd1 _06825_/B sky130_fd_sc_hd__nand3_2
XFILLER_62_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06751_ _13479_/Q vssd1 vssd1 vccd1 vccd1 _06751_/Y sky130_fd_sc_hd__inv_2
XFILLER_83_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_75_clk clkbuf_5_15_0_clk/X vssd1 vssd1 vccd1 vccd1 _15446_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_58_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06682_ _14902_/Q vssd1 vssd1 vccd1 vccd1 _06682_/Y sky130_fd_sc_hd__inv_2
X_09470_ _14449_/Q _08540_/B _13130_/C1 _09469_/X vssd1 vssd1 vccd1 vccd1 _09470_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_36_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_836 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08421_ _08421_/A _08421_/B vssd1 vssd1 vccd1 vccd1 _08421_/Y sky130_fd_sc_hd__nand2_2
XFILLER_52_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08352_ _08244_/A _13762_/Q _15410_/Q _08244_/B vssd1 vssd1 vccd1 vccd1 _08352_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_149_201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07303_ _07294_/Y _07295_/X _07301_/Y _07302_/X vssd1 vssd1 vccd1 vccd1 _07351_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_177_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08283_ _11298_/A _11351_/C1 _08282_/X _08232_/A _13717_/Q vssd1 vssd1 vccd1 vccd1
+ _13717_/D sky130_fd_sc_hd__a32o_1
XFILLER_137_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07234_ _15329_/Q _15485_/Q _07335_/S vssd1 vssd1 vccd1 vccd1 _07235_/B sky130_fd_sc_hd__mux2_8
XFILLER_146_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07165_ _15339_/Q _15046_/Q _07193_/S vssd1 vssd1 vccd1 vccd1 _07165_/X sky130_fd_sc_hd__mux2_4
XFILLER_118_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07096_ _14644_/Q _14676_/Q _07096_/S vssd1 vssd1 vccd1 vccd1 _07096_/X sky130_fd_sc_hd__mux2_1
XFILLER_160_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_432 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_808 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout201 _09763_/Y vssd1 vssd1 vccd1 vccd1 _09790_/S sky130_fd_sc_hd__buf_12
Xfanout212 _09596_/Y vssd1 vssd1 vccd1 vccd1 _09628_/S sky130_fd_sc_hd__buf_12
Xfanout223 _08012_/A2 vssd1 vssd1 vccd1 vccd1 _08022_/B sky130_fd_sc_hd__buf_6
XFILLER_87_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout234 _07614_/A vssd1 vssd1 vccd1 vccd1 _07629_/A sky130_fd_sc_hd__buf_8
XFILLER_99_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout245 _08747_/B1 vssd1 vssd1 vccd1 vccd1 _08691_/B1 sky130_fd_sc_hd__buf_12
XFILLER_59_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout256 _07783_/X vssd1 vssd1 vccd1 vccd1 _07903_/A sky130_fd_sc_hd__buf_8
X_09806_ _14172_/Q _11861_/A1 _09823_/S vssd1 vssd1 vccd1 vccd1 _14172_/D sky130_fd_sc_hd__mux2_1
Xfanout267 _08524_/Y vssd1 vssd1 vccd1 vccd1 _08749_/A2 sky130_fd_sc_hd__buf_12
Xfanout278 _09536_/A2 vssd1 vssd1 vccd1 vccd1 _09558_/A2 sky130_fd_sc_hd__buf_12
XFILLER_115_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07998_ _14758_/Q _07971_/A _07997_/Y _08002_/C1 vssd1 vssd1 vccd1 vccd1 _13565_/D
+ sky130_fd_sc_hd__o211a_1
Xfanout289 _13347_/A0 vssd1 vssd1 vccd1 vccd1 _11847_/A1 sky130_fd_sc_hd__buf_6
XFILLER_75_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09737_ _14105_/Q _13325_/A0 _09757_/S vssd1 vssd1 vccd1 vccd1 _14105_/D sky130_fd_sc_hd__mux2_1
XFILLER_86_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06949_ _06740_/Y _13483_/Q _14491_/Q _06743_/Y vssd1 vssd1 vccd1 vccd1 _06963_/A
+ sky130_fd_sc_hd__a2bb2o_1
Xclkbuf_leaf_66_clk clkbuf_5_11_0_clk/X vssd1 vssd1 vccd1 vccd1 _15014_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_27_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09668_ _14039_/Q _11681_/A0 _09690_/S vssd1 vssd1 vccd1 vccd1 _14039_/D sky130_fd_sc_hd__mux2_1
XFILLER_15_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08619_ _08722_/A _08619_/B _08619_/C vssd1 vssd1 vccd1 vccd1 _08619_/X sky130_fd_sc_hd__or3_1
XTAP_1225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09599_ _13973_/Q _11854_/A1 _09628_/S vssd1 vssd1 vccd1 vccd1 _13973_/D sky130_fd_sc_hd__mux2_1
XTAP_1236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11630_ _11629_/Y _15072_/Q _11641_/S vssd1 vssd1 vccd1 vccd1 _15072_/D sky130_fd_sc_hd__mux2_1
XFILLER_145_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11561_ _11561_/A _11561_/B vssd1 vssd1 vccd1 vccd1 _11563_/B sky130_fd_sc_hd__xor2_2
XFILLER_183_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13300_ _12725_/Y _15632_/Q _13300_/S vssd1 vssd1 vccd1 vccd1 _15632_/D sky130_fd_sc_hd__mux2_1
XFILLER_10_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10512_ _10541_/A _10512_/B vssd1 vssd1 vccd1 vccd1 _10528_/C sky130_fd_sc_hd__nand2b_1
X_14280_ _15669_/CLK _14280_/D vssd1 vssd1 vccd1 vccd1 _14280_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11492_ _11492_/A _11502_/B vssd1 vssd1 vccd1 vccd1 _11505_/D sky130_fd_sc_hd__nor2_1
XFILLER_155_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13231_ _15577_/Q _13219_/S _13230_/X vssd1 vssd1 vccd1 vccd1 _15577_/D sky130_fd_sc_hd__o21a_1
X_10443_ _10537_/B _10443_/B vssd1 vssd1 vccd1 vccd1 _10471_/C sky130_fd_sc_hd__or2_1
XFILLER_10_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13162_ _13217_/A _13162_/B vssd1 vssd1 vccd1 vccd1 _13162_/Y sky130_fd_sc_hd__nand2_1
XFILLER_152_944 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10374_ _07297_/A _10360_/B _10373_/X vssd1 vssd1 vccd1 vccd1 _11476_/A sky130_fd_sc_hd__a21oi_4
XFILLER_136_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_432 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12113_ _12596_/A _12113_/B _12113_/C vssd1 vssd1 vccd1 vccd1 _12113_/X sky130_fd_sc_hd__and3_1
XFILLER_3_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13093_ _15514_/Q _13093_/A2 _13042_/A _13092_/X vssd1 vssd1 vccd1 vccd1 _15514_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_151_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12044_ _12596_/A _12044_/B _12044_/C vssd1 vssd1 vccd1 vccd1 _12044_/X sky130_fd_sc_hd__and3_2
XFILLER_27_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13995_ _14542_/CLK _13995_/D vssd1 vssd1 vccd1 vccd1 _13995_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_57_clk clkbuf_5_11_0_clk/X vssd1 vssd1 vccd1 vccd1 _15021_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_3150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12946_ _13129_/A _12946_/B vssd1 vssd1 vccd1 vccd1 _12946_/Y sky130_fd_sc_hd__nor2_4
XTAP_3161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15665_ _15665_/CLK _15665_/D vssd1 vssd1 vccd1 vccd1 _15665_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_45_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12877_ _15405_/Q _15590_/Q _12933_/S vssd1 vssd1 vccd1 vccd1 _15405_/D sky130_fd_sc_hd__mux2_1
XFILLER_34_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14616_ _15620_/CLK _14616_/D vssd1 vssd1 vccd1 vccd1 _14616_/Q sky130_fd_sc_hd__dfxtp_1
X_11828_ _15250_/Q _11861_/A1 _11849_/S vssd1 vssd1 vccd1 vccd1 _15250_/D sky130_fd_sc_hd__mux2_1
X_15596_ _15596_/CLK _15596_/D vssd1 vssd1 vccd1 vccd1 _15596_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14547_ _15226_/CLK _14547_/D vssd1 vssd1 vccd1 vccd1 _14547_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_187_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11759_ _13082_/B2 _15187_/Q _11774_/S vssd1 vssd1 vccd1 vccd1 _15187_/D sky130_fd_sc_hd__mux2_1
XFILLER_41_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14478_ _15518_/CLK _14478_/D vssd1 vssd1 vccd1 vccd1 _14478_/Q sky130_fd_sc_hd__dfxtp_1
X_13429_ _15381_/CLK _13429_/D vssd1 vssd1 vccd1 vccd1 _13429_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_60_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08970_ _08968_/X _08969_/X _08959_/X vssd1 vssd1 vccd1 vccd1 _08970_/X sky130_fd_sc_hd__o21a_2
XFILLER_142_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07921_ _13545_/Q _07921_/B vssd1 vssd1 vccd1 vccd1 _07921_/X sky130_fd_sc_hd__xor2_1
XFILLER_130_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07852_ _13527_/Q _07858_/D vssd1 vssd1 vccd1 vccd1 _07852_/X sky130_fd_sc_hd__or2_1
XFILLER_57_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06803_ _13732_/Q _12615_/A1 _08405_/B _06665_/Y _06802_/X vssd1 vssd1 vccd1 vccd1
+ _06806_/B sky130_fd_sc_hd__o221a_1
Xinput1 ext_read_data[0] vssd1 vssd1 vccd1 vccd1 input1/X sky130_fd_sc_hd__buf_4
XFILLER_84_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07783_ _07783_/A _07783_/B _07783_/C vssd1 vssd1 vccd1 vccd1 _07783_/X sky130_fd_sc_hd__or3_4
Xclkbuf_leaf_48_clk clkbuf_5_8_0_clk/X vssd1 vssd1 vccd1 vccd1 _15556_/CLK sky130_fd_sc_hd__clkbuf_16
X_09522_ _14097_/Q _09522_/A2 _09522_/B1 _14065_/Q _09532_/A vssd1 vssd1 vccd1 vccd1
+ _09522_/X sky130_fd_sc_hd__a221o_1
X_06734_ _14495_/Q vssd1 vssd1 vccd1 vccd1 _06734_/Y sky130_fd_sc_hd__inv_2
XFILLER_188_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09453_ _13934_/Q _13154_/S vssd1 vssd1 vccd1 vccd1 _09453_/X sky130_fd_sc_hd__and2_1
XFILLER_149_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06665_ _13731_/Q vssd1 vssd1 vccd1 vccd1 _06665_/Y sky130_fd_sc_hd__inv_2
XFILLER_25_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08404_ _13736_/Q _08390_/X _13138_/S vssd1 vssd1 vccd1 vccd1 _13736_/D sky130_fd_sc_hd__mux2_1
X_09384_ _15099_/Q _08519_/B _09519_/B1 _08501_/A vssd1 vssd1 vccd1 vccd1 _09384_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_52_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08335_ _07295_/X _10523_/A2 _08334_/X vssd1 vssd1 vccd1 vccd1 _11440_/A sky130_fd_sc_hd__a21o_4
XFILLER_178_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08266_ _08266_/A vssd1 vssd1 vccd1 vccd1 _08266_/Y sky130_fd_sc_hd__inv_2
X_07217_ _07215_/Y _07213_/X _07211_/X _07210_/Y vssd1 vssd1 vccd1 vccd1 _07356_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_08197_ _13688_/Q _13326_/A0 _08216_/S vssd1 vssd1 vccd1 vccd1 _13688_/D sky130_fd_sc_hd__mux2_1
XFILLER_118_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_1042 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07148_ _14854_/Q _14846_/Q _14838_/Q _14830_/Q _07146_/S _07104_/C vssd1 vssd1 vccd1
+ vccd1 _07149_/B sky130_fd_sc_hd__mux4_1
XFILLER_105_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_1075 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07079_ _07078_/X _13605_/Q _12764_/S vssd1 vssd1 vccd1 vccd1 _07079_/X sky130_fd_sc_hd__mux2_1
XFILLER_117_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_935 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10090_ _14446_/Q _13343_/A0 _10092_/S vssd1 vssd1 vccd1 vccd1 _14446_/D sky130_fd_sc_hd__mux2_1
XFILLER_133_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_39_clk clkbuf_5_12_0_clk/X vssd1 vssd1 vccd1 vccd1 _15587_/CLK sky130_fd_sc_hd__clkbuf_16
X_12800_ _15069_/Q _12834_/B vssd1 vssd1 vccd1 vccd1 _12800_/X sky130_fd_sc_hd__or2_1
XFILLER_56_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13780_ _15397_/CLK _13780_/D vssd1 vssd1 vccd1 vccd1 _13780_/Q sky130_fd_sc_hd__dfxtp_4
X_10992_ _11318_/S _10992_/B vssd1 vssd1 vccd1 vccd1 _10992_/X sky130_fd_sc_hd__or2_1
XFILLER_83_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_1024 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12731_ _15353_/Q _12732_/B vssd1 vssd1 vccd1 vccd1 _12745_/C sky130_fd_sc_hd__and2_2
XTAP_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15450_ _15635_/CLK _15450_/D vssd1 vssd1 vccd1 vccd1 _15450_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12662_ _13420_/Q _12661_/X _12662_/S vssd1 vssd1 vccd1 vccd1 _12663_/B sky130_fd_sc_hd__mux2_1
XTAP_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14401_ _15285_/CLK _14401_/D vssd1 vssd1 vccd1 vccd1 _14401_/Q sky130_fd_sc_hd__dfxtp_1
X_11613_ _11613_/A _11613_/B vssd1 vssd1 vccd1 vccd1 _11613_/Y sky130_fd_sc_hd__xnor2_1
XTAP_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15381_ _15381_/CLK _15381_/D vssd1 vssd1 vccd1 vccd1 _15381_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_184_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12593_ _12586_/X _12588_/X _12590_/X _12592_/X _06671_/A vssd1 vssd1 vccd1 vccd1
+ _12593_/X sky130_fd_sc_hd__o221a_1
XFILLER_168_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14332_ _15281_/CLK _14332_/D vssd1 vssd1 vccd1 vccd1 _14332_/Q sky130_fd_sc_hd__dfxtp_1
X_11544_ _11544_/A _11544_/B vssd1 vssd1 vccd1 vccd1 _11546_/C sky130_fd_sc_hd__nor2_1
XFILLER_128_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14263_ _15276_/CLK _14263_/D vssd1 vssd1 vccd1 vccd1 _14263_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_171_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11475_ _11475_/A _11475_/B vssd1 vssd1 vccd1 vccd1 _11476_/D sky130_fd_sc_hd__nor2_1
XFILLER_183_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13214_ _13214_/A _13214_/B vssd1 vssd1 vccd1 vccd1 _13214_/Y sky130_fd_sc_hd__nor2_1
XFILLER_109_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10426_ _11632_/A vssd1 vssd1 vccd1 vccd1 _10530_/B sky130_fd_sc_hd__inv_2
X_14194_ _15680_/CLK _14194_/D vssd1 vssd1 vccd1 vccd1 _14194_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_124_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13145_ _09466_/A _15543_/Q _13154_/S vssd1 vssd1 vccd1 vccd1 _15543_/D sky130_fd_sc_hd__mux2_1
X_10357_ _08240_/A _13793_/Q _13761_/Q _08237_/A vssd1 vssd1 vccd1 vccd1 _10357_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_151_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13076_ _12981_/X _13104_/A2 _13104_/B1 _07424_/X vssd1 vssd1 vccd1 vccd1 _13076_/X
+ sky130_fd_sc_hd__a22o_1
X_10288_ _14673_/Q _14826_/Q _10735_/S vssd1 vssd1 vccd1 vccd1 _14673_/D sky130_fd_sc_hd__mux2_1
X_12027_ _12023_/X _12024_/X _12582_/A vssd1 vssd1 vccd1 vccd1 _12027_/X sky130_fd_sc_hd__mux2_1
XFILLER_78_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13978_ _15276_/CLK _13978_/D vssd1 vssd1 vccd1 vccd1 _13978_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12929_ _15457_/Q _15643_/Q _12929_/S vssd1 vssd1 vccd1 vccd1 _15457_/D sky130_fd_sc_hd__mux2_1
XFILLER_34_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15648_ _15648_/CLK _15648_/D vssd1 vssd1 vccd1 vccd1 _15648_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15579_ _15579_/CLK _15579_/D vssd1 vssd1 vccd1 vccd1 _15579_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08120_ input31/X input8/X _08133_/S vssd1 vssd1 vccd1 vccd1 _08120_/X sky130_fd_sc_hd__mux2_1
X_08051_ _14744_/Q _13622_/Q _08066_/S vssd1 vssd1 vccd1 vccd1 _13622_/D sky130_fd_sc_hd__mux2_1
XFILLER_174_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07002_ _14718_/Q _07783_/A _08027_/A vssd1 vssd1 vccd1 vccd1 _10099_/B sky130_fd_sc_hd__nor3_4
XFILLER_134_229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08953_ _15276_/Q _15244_/Q _15212_/Q _15143_/Q _09230_/S _09234_/S1 vssd1 vssd1
+ vccd1 vccd1 _08953_/X sky130_fd_sc_hd__mux4_1
XFILLER_88_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07904_ _14765_/Q _07903_/A _07903_/Y _08016_/C1 vssd1 vssd1 vccd1 vccd1 _13540_/D
+ sky130_fd_sc_hd__o211a_1
X_08884_ _13905_/Q _11816_/A1 _08885_/S vssd1 vssd1 vccd1 vccd1 _13905_/D sky130_fd_sc_hd__mux2_1
XFILLER_84_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07835_ _14747_/Q _07830_/A _07834_/Y _12788_/C1 vssd1 vssd1 vccd1 vccd1 _13522_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_3908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07766_ _07764_/Y _07769_/B _07777_/A vssd1 vssd1 vccd1 vccd1 _07766_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_72_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09505_ _13904_/Q _09522_/A2 _09519_/B1 _14419_/Q _08507_/A vssd1 vssd1 vccd1 vccd1
+ _09505_/X sky130_fd_sc_hd__a221o_1
X_06717_ _15386_/Q vssd1 vssd1 vccd1 vccd1 _06717_/Y sky130_fd_sc_hd__inv_2
XFILLER_53_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07697_ _13487_/Q _07697_/B vssd1 vssd1 vccd1 vccd1 _07698_/B sky130_fd_sc_hd__xnor2_1
XFILLER_24_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09436_ _15299_/Q _15267_/Q _15235_/Q _15166_/Q _09444_/S _09446_/A1 vssd1 vssd1
+ vccd1 vccd1 _09436_/X sky130_fd_sc_hd__mux4_1
XFILLER_24_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_5_5_0_clk clkbuf_5_5_0_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_5_5_0_clk/X sky130_fd_sc_hd__clkbuf_8
XFILLER_12_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09367_ _09365_/X _09366_/X _12573_/A _09356_/X vssd1 vssd1 vccd1 vccd1 _09367_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_12_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08318_ _11356_/B _10986_/A _08316_/B _08317_/X vssd1 vssd1 vccd1 vccd1 _08318_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_21_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09298_ _15127_/Q _15095_/Q _15668_/Q _13402_/Q _09484_/S _08519_/A vssd1 vssd1 vccd1
+ vccd1 _09298_/X sky130_fd_sc_hd__mux4_1
XANTENNA_50 _07177_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_61 _07170_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_72 _07147_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_83 _07101_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08249_ _11371_/A _11362_/B vssd1 vssd1 vccd1 vccd1 _08249_/Y sky130_fd_sc_hd__nor2_8
XANTENNA_94 _08638_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11260_ _08376_/X _11259_/X _11297_/S vssd1 vssd1 vccd1 vccd1 _11260_/X sky130_fd_sc_hd__mux2_1
XFILLER_106_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10211_ input5/X _14596_/Q _13284_/S vssd1 vssd1 vccd1 vccd1 _14596_/D sky130_fd_sc_hd__mux2_1
XFILLER_97_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11191_ _11199_/A _11191_/B vssd1 vssd1 vccd1 vccd1 _11191_/Y sky130_fd_sc_hd__nor2_1
XFILLER_106_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10142_ _14527_/Q _13328_/A0 _10159_/S vssd1 vssd1 vccd1 vccd1 _14527_/D sky130_fd_sc_hd__mux2_1
XFILLER_79_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14950_ _15017_/CLK _14950_/D vssd1 vssd1 vccd1 vccd1 _14950_/Q sky130_fd_sc_hd__dfxtp_1
X_10073_ _14429_/Q _12967_/A1 _10092_/S vssd1 vssd1 vccd1 vccd1 _14429_/D sky130_fd_sc_hd__mux2_1
XFILLER_153_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13901_ _15315_/CLK _13901_/D vssd1 vssd1 vccd1 vccd1 _13901_/Q sky130_fd_sc_hd__dfxtp_1
X_14881_ _15452_/CLK _14881_/D vssd1 vssd1 vccd1 vccd1 _14881_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13832_ _15161_/CLK _13832_/D vssd1 vssd1 vccd1 vccd1 _13832_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13763_ _15613_/CLK _13763_/D vssd1 vssd1 vccd1 vccd1 _13763_/Q sky130_fd_sc_hd__dfxtp_1
X_10975_ _11013_/A _13226_/B _11305_/B vssd1 vssd1 vccd1 vccd1 _10979_/B sky130_fd_sc_hd__a21boi_1
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12714_ _13427_/Q _12713_/X _12728_/S vssd1 vssd1 vccd1 vccd1 _12715_/B sky130_fd_sc_hd__mux2_1
X_15502_ _15508_/CLK _15502_/D vssd1 vssd1 vccd1 vccd1 _15502_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13694_ _15315_/CLK _13694_/D vssd1 vssd1 vccd1 vccd1 _13694_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15433_ _15619_/CLK _15433_/D vssd1 vssd1 vccd1 vccd1 _15433_/Q sky130_fd_sc_hd__dfxtp_1
X_12645_ _12657_/C _12645_/B vssd1 vssd1 vccd1 vccd1 _12645_/Y sky130_fd_sc_hd__nor2_1
XFILLER_12_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15364_ _15644_/CLK _15364_/D vssd1 vssd1 vccd1 vccd1 _15364_/Q sky130_fd_sc_hd__dfxtp_2
X_12576_ _14484_/Q _14452_/Q _13873_/Q _14226_/Q _12430_/S _12563_/A vssd1 vssd1 vccd1
+ vccd1 _12576_/X sky130_fd_sc_hd__mux4_1
XFILLER_178_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_894 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14315_ _15336_/CLK _14315_/D vssd1 vssd1 vccd1 vccd1 _14315_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_184_663 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11527_ _11526_/Y _15061_/Q _11614_/S vssd1 vssd1 vccd1 vccd1 _15061_/D sky130_fd_sc_hd__mux2_1
XFILLER_11_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_156_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15295_ _15295_/CLK _15295_/D vssd1 vssd1 vccd1 vccd1 _15295_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_172_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14246_ _15301_/CLK _14246_/D vssd1 vssd1 vccd1 vccd1 _14246_/Q sky130_fd_sc_hd__dfxtp_1
X_11458_ _11472_/A _11458_/B vssd1 vssd1 vccd1 vccd1 _11505_/A sky130_fd_sc_hd__nor2_1
XFILLER_172_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10409_ _11414_/A _13168_/B vssd1 vssd1 vccd1 vccd1 _10555_/A sky130_fd_sc_hd__xnor2_1
X_14177_ _15663_/CLK _14177_/D vssd1 vssd1 vccd1 vccd1 _14177_/Q sky130_fd_sc_hd__dfxtp_1
X_11389_ _11414_/D _11389_/B _11389_/C vssd1 vssd1 vccd1 vccd1 _11390_/C sky130_fd_sc_hd__nand3b_2
XFILLER_125_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13128_ _09382_/A _13124_/X _13126_/X _13127_/X vssd1 vssd1 vccd1 vccd1 _13129_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_139_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13059_ _15497_/Q _13081_/A2 _13105_/B1 _13058_/X vssd1 vssd1 vccd1 vccd1 _15497_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_23_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07620_ _07621_/A _07621_/B vssd1 vssd1 vccd1 vccd1 _07620_/X sky130_fd_sc_hd__and2_1
XFILLER_4_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07551_ _14737_/Q _07644_/A _07550_/Y _08084_/C1 vssd1 vssd1 vccd1 vccd1 _13448_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_35_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_1052 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07482_ _14672_/Q _07490_/B _07482_/C vssd1 vssd1 vccd1 vccd1 _07482_/X sky130_fd_sc_hd__and3_1
XFILLER_50_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09221_ _09221_/A _09221_/B vssd1 vssd1 vccd1 vccd1 _09221_/X sky130_fd_sc_hd__or2_1
XFILLER_50_945 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09152_ _09406_/S1 _09150_/X _09151_/X vssd1 vssd1 vccd1 vccd1 _09152_/X sky130_fd_sc_hd__a21o_1
XFILLER_148_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08103_ _13651_/Q _10344_/S _08096_/X _08102_/X vssd1 vssd1 vccd1 vccd1 _13651_/D
+ sky130_fd_sc_hd__a22o_1
X_09083_ _14463_/Q _14431_/Q _13852_/Q _14205_/Q _09190_/S _09429_/S1 vssd1 vssd1
+ vccd1 vccd1 _09083_/X sky130_fd_sc_hd__mux4_1
XFILLER_108_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08034_ _13575_/Q _14745_/Q _08039_/S vssd1 vssd1 vccd1 vccd1 _13575_/D sky130_fd_sc_hd__mux2_1
XFILLER_163_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09985_ _11872_/A1 _14344_/Q _09996_/S vssd1 vssd1 vccd1 vccd1 _14344_/D sky130_fd_sc_hd__mux2_1
XFILLER_89_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08936_ _08510_/B _08932_/X _08935_/X _08931_/X vssd1 vssd1 vccd1 vccd1 _08949_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_69_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08867_ _13888_/Q _13078_/B2 _08880_/S vssd1 vssd1 vccd1 vccd1 _13888_/D sky130_fd_sc_hd__mux2_1
XFILLER_123_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07818_ _13518_/Q _07825_/D vssd1 vssd1 vccd1 vccd1 _07819_/B sky130_fd_sc_hd__xnor2_1
XTAP_3749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08798_ _13332_/A0 _13824_/Q _08811_/S vssd1 vssd1 vccd1 vccd1 _13824_/D sky130_fd_sc_hd__mux2_1
XFILLER_57_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07749_ _13501_/Q _07757_/D vssd1 vssd1 vccd1 vccd1 _07750_/B sky130_fd_sc_hd__xnor2_1
X_10760_ _15424_/Q _14792_/Q _10765_/S vssd1 vssd1 vccd1 vccd1 _14792_/D sky130_fd_sc_hd__mux2_1
XFILLER_73_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09419_ _09446_/A1 _09419_/A2 _09418_/X _06676_/A vssd1 vssd1 vccd1 vccd1 _09419_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_186_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10691_ _15017_/Q _10717_/A2 _10718_/A2 _14985_/Q _10717_/C1 vssd1 vssd1 vccd1 vccd1
+ _10691_/X sky130_fd_sc_hd__a221o_1
XFILLER_9_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12430_ _14090_/Q _14058_/Q _12430_/S vssd1 vssd1 vccd1 vccd1 _12430_/X sky130_fd_sc_hd__mux2_1
XFILLER_185_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12361_ _14087_/Q _14055_/Q _12541_/S vssd1 vssd1 vccd1 vccd1 _12361_/X sky130_fd_sc_hd__mux2_1
XFILLER_138_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14100_ _15650_/CLK _14100_/D vssd1 vssd1 vccd1 vccd1 _14100_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_154_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11312_ _11312_/A _11312_/B vssd1 vssd1 vccd1 vccd1 _11312_/Y sky130_fd_sc_hd__nand2_1
XFILLER_154_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15080_ _15649_/CLK _15080_/D vssd1 vssd1 vccd1 vccd1 _15080_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_180_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12292_ _14084_/Q _14052_/Q _12614_/S vssd1 vssd1 vccd1 vccd1 _12292_/X sky130_fd_sc_hd__mux2_1
XFILLER_4_323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14031_ _15127_/CLK _14031_/D vssd1 vssd1 vccd1 vccd1 _14031_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_1055 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11243_ _08375_/Y _11242_/Y _11318_/S vssd1 vssd1 vccd1 vccd1 _11243_/X sky130_fd_sc_hd__mux2_1
XFILLER_106_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11174_ _14979_/Q _11164_/S _11173_/X vssd1 vssd1 vccd1 vccd1 _14979_/D sky130_fd_sc_hd__o21a_1
XFILLER_68_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_96 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10125_ _14511_/Q _14759_/Q _10131_/S vssd1 vssd1 vccd1 vccd1 _14511_/D sky130_fd_sc_hd__mux2_1
XFILLER_95_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_831 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_595 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10056_ _14413_/Q _13098_/B2 _10064_/S vssd1 vssd1 vccd1 vccd1 _14413_/D sky130_fd_sc_hd__mux2_1
X_14933_ _14997_/CLK _14933_/D vssd1 vssd1 vccd1 vccd1 _14933_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_169_1022 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14864_ _15619_/CLK _14864_/D vssd1 vssd1 vccd1 vccd1 _14864_/Q sky130_fd_sc_hd__dfxtp_1
X_13815_ _15176_/CLK _13815_/D vssd1 vssd1 vccd1 vccd1 _13815_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_28_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14795_ _15612_/CLK _14795_/D vssd1 vssd1 vccd1 vccd1 hold6/A sky130_fd_sc_hd__dfxtp_1
XFILLER_50_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13746_ _14703_/CLK _13746_/D vssd1 vssd1 vccd1 vccd1 _13746_/Q sky130_fd_sc_hd__dfxtp_1
X_10958_ _11317_/B _10958_/B vssd1 vssd1 vccd1 vccd1 _10958_/Y sky130_fd_sc_hd__nor2_1
XFILLER_32_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13677_ _15622_/CLK _13677_/D vssd1 vssd1 vccd1 vccd1 _13677_/Q sky130_fd_sc_hd__dfxtp_1
X_10889_ _14921_/Q _15552_/Q _13134_/A vssd1 vssd1 vccd1 vccd1 _14921_/D sky130_fd_sc_hd__mux2_1
X_15416_ _15635_/CLK _15416_/D vssd1 vssd1 vccd1 vccd1 _15416_/Q sky130_fd_sc_hd__dfxtp_4
X_12628_ _15338_/Q _12759_/B _12627_/Y _12832_/C1 vssd1 vssd1 vccd1 vccd1 _15338_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_8_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_1072 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15347_ _15630_/CLK _15347_/D vssd1 vssd1 vccd1 vccd1 _15347_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_184_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_172_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12559_ _12559_/A _12559_/B vssd1 vssd1 vccd1 vccd1 _12559_/X sky130_fd_sc_hd__or2_1
XFILLER_117_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15278_ _15278_/CLK _15278_/D vssd1 vssd1 vccd1 vccd1 _15278_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_346 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14229_ _15676_/CLK _14229_/D vssd1 vssd1 vccd1 vccd1 _14229_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout608 _12470_/S vssd1 vssd1 vccd1 vccd1 _12079_/S sky130_fd_sc_hd__buf_12
XFILLER_98_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout619 _12545_/S vssd1 vssd1 vccd1 vccd1 _12543_/S sky130_fd_sc_hd__buf_12
XTAP_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09770_ _14137_/Q _13325_/A0 _09790_/S vssd1 vssd1 vccd1 vccd1 _14137_/D sky130_fd_sc_hd__mux2_1
XTAP_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06982_ _08240_/A _13120_/S _08777_/A _14596_/Q vssd1 vssd1 vccd1 vccd1 _14767_/D
+ sky130_fd_sc_hd__a22o_1
XTAP_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08721_ _15372_/Q _08748_/A2 _08719_/X _08720_/X vssd1 vssd1 vccd1 vccd1 _08722_/C
+ sky130_fd_sc_hd__a211o_1
XTAP_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_1043 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08652_ _10765_/S _08652_/B _08652_/C vssd1 vssd1 vccd1 vccd1 _08652_/X sky130_fd_sc_hd__or3_4
XFILLER_113_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_1087 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07603_ _13462_/Q _13461_/Q _07603_/C _07603_/D vssd1 vssd1 vccd1 vccd1 _07610_/C
+ sky130_fd_sc_hd__and4_2
XFILLER_82_856 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08583_ _15392_/Q _08690_/A2 _08690_/B1 _13437_/Q vssd1 vssd1 vccd1 vccd1 _08583_/X
+ sky130_fd_sc_hd__a22o_1
X_07534_ _14764_/Q _13443_/Q _07535_/S vssd1 vssd1 vccd1 vccd1 _13443_/D sky130_fd_sc_hd__mux2_1
XFILLER_22_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07465_ _13341_/A0 _13405_/Q _07481_/S vssd1 vssd1 vccd1 vccd1 _13405_/D sky130_fd_sc_hd__mux2_1
XFILLER_22_444 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09204_ _14469_/Q _14437_/Q _13858_/Q _14211_/Q _09441_/S _09448_/S1 vssd1 vssd1
+ vccd1 vccd1 _09204_/X sky130_fd_sc_hd__mux4_1
XFILLER_22_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_630 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07396_ _14739_/Q _07395_/X _07500_/S vssd1 vssd1 vccd1 vccd1 _07396_/X sky130_fd_sc_hd__mux2_2
XFILLER_72_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09135_ _09449_/B2 _09131_/X _09134_/X vssd1 vssd1 vccd1 vccd1 _09135_/X sky130_fd_sc_hd__a21o_1
XFILLER_147_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09066_ _15116_/Q _09536_/A2 _09065_/X _09450_/B1 vssd1 vssd1 vccd1 vccd1 _09066_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_136_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08017_ _13571_/Q _13570_/Q _13569_/Q _08017_/D vssd1 vssd1 vccd1 vccd1 _08021_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_135_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_252_clk clkbuf_5_1_0_clk/X vssd1 vssd1 vccd1 vccd1 _15289_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_77_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09968_ _13322_/A0 _14327_/Q _09991_/S vssd1 vssd1 vccd1 vccd1 _14327_/D sky130_fd_sc_hd__mux2_1
X_08919_ _09550_/A1 _08917_/X _08918_/X vssd1 vssd1 vccd1 vccd1 _08920_/C sky130_fd_sc_hd__a21o_1
X_09899_ _11852_/A1 _14260_/Q _09925_/S vssd1 vssd1 vccd1 vccd1 _14260_/D sky130_fd_sc_hd__mux2_1
XTAP_3502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11930_ _15307_/Q _13139_/S _11929_/X vssd1 vssd1 vccd1 vccd1 _15307_/D sky130_fd_sc_hd__a21o_1
XTAP_3524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_119 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_171 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11861_ _15282_/Q _11861_/A1 _11878_/S vssd1 vssd1 vccd1 vccd1 _15282_/D sky130_fd_sc_hd__mux2_1
XTAP_2834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13600_ _15636_/CLK _13600_/D vssd1 vssd1 vccd1 vccd1 _13600_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_2856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10812_ _14844_/Q _07280_/A _12481_/A vssd1 vssd1 vccd1 vccd1 _14844_/D sky130_fd_sc_hd__mux2_1
XTAP_2867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14580_ _15303_/CLK _14580_/D vssd1 vssd1 vccd1 vccd1 _14580_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11792_ _15215_/Q _11858_/A1 _11817_/S vssd1 vssd1 vccd1 vccd1 _15215_/D sky130_fd_sc_hd__mux2_1
XTAP_2889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13531_ _13565_/CLK _13531_/D vssd1 vssd1 vccd1 vccd1 _13531_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10743_ _15407_/Q _14775_/Q _10759_/S vssd1 vssd1 vccd1 vccd1 _14775_/D sky130_fd_sc_hd__mux2_1
XFILLER_158_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_736 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13462_ _15385_/CLK _13462_/D vssd1 vssd1 vccd1 vccd1 _13462_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_186_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10674_ _15062_/Q _10714_/A2 _10671_/X _10673_/X vssd1 vssd1 vccd1 vccd1 _10674_/X
+ sky130_fd_sc_hd__o22a_4
XFILLER_13_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15201_ _15226_/CLK _15201_/D vssd1 vssd1 vccd1 vccd1 _15201_/Q sky130_fd_sc_hd__dfxtp_1
X_12413_ _15328_/Q _13093_/A2 _12412_/X vssd1 vssd1 vccd1 vccd1 _15328_/D sky130_fd_sc_hd__a21o_1
XFILLER_185_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13393_ _15674_/CLK _13393_/D vssd1 vssd1 vccd1 vccd1 _13393_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_167_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15132_ _15673_/CLK _15132_/D vssd1 vssd1 vccd1 vccd1 _15132_/Q sky130_fd_sc_hd__dfxtp_1
X_12344_ _15325_/Q _13149_/S _12343_/X vssd1 vssd1 vccd1 vccd1 _15325_/D sky130_fd_sc_hd__a21o_1
XFILLER_175_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15063_ _15422_/CLK _15063_/D vssd1 vssd1 vccd1 vccd1 _15063_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_182_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12275_ _15322_/Q _13119_/S _12274_/X vssd1 vssd1 vccd1 vccd1 _15322_/D sky130_fd_sc_hd__a21o_1
XFILLER_4_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14014_ _15285_/CLK _14014_/D vssd1 vssd1 vccd1 vccd1 _14014_/Q sky130_fd_sc_hd__dfxtp_1
X_11226_ _10528_/C _15014_/Q _11232_/S vssd1 vssd1 vccd1 vccd1 _15014_/D sky130_fd_sc_hd__mux2_1
XFILLER_49_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_243_clk clkbuf_5_4_0_clk/X vssd1 vssd1 vccd1 vccd1 _14083_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_68_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11157_ _11347_/A _11107_/X _11156_/Y _11414_/A vssd1 vssd1 vccd1 vccd1 _11157_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_136_1076 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_959 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10108_ _14494_/Q _14742_/Q _10124_/S vssd1 vssd1 vccd1 vccd1 _14494_/D sky130_fd_sc_hd__mux2_1
X_11088_ _11033_/Y _11045_/Y _11088_/S vssd1 vssd1 vccd1 vccd1 _11088_/X sky130_fd_sc_hd__mux2_1
XFILLER_49_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10039_ _14396_/Q _11858_/A1 _10064_/S vssd1 vssd1 vccd1 vccd1 _14396_/D sky130_fd_sc_hd__mux2_1
XFILLER_49_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14916_ _15670_/CLK _14916_/D vssd1 vssd1 vccd1 vccd1 _14916_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14847_ _15536_/CLK _14847_/D vssd1 vssd1 vccd1 vccd1 _14847_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14778_ _15596_/CLK _14778_/D vssd1 vssd1 vccd1 vccd1 _14778_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13729_ _15530_/CLK _13729_/D vssd1 vssd1 vccd1 vccd1 _13729_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_90_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07250_ _15325_/Q _15481_/Q _07335_/S vssd1 vssd1 vccd1 vccd1 _07251_/A sky130_fd_sc_hd__mux2_8
XFILLER_149_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07181_ _15355_/Q _15062_/Q _07188_/S vssd1 vssd1 vccd1 vccd1 _07181_/X sky130_fd_sc_hd__mux2_8
XFILLER_173_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout405 _13156_/Y vssd1 vssd1 vccd1 vccd1 _13241_/A2 sky130_fd_sc_hd__buf_8
Xfanout416 _10948_/B vssd1 vssd1 vccd1 vccd1 _10929_/B sky130_fd_sc_hd__clkbuf_4
Xclkbuf_leaf_234_clk clkbuf_5_5_0_clk/X vssd1 vssd1 vccd1 vccd1 _15276_/CLK sky130_fd_sc_hd__clkbuf_16
X_09822_ _14188_/Q _11877_/A1 _09823_/S vssd1 vssd1 vccd1 vccd1 _14188_/D sky130_fd_sc_hd__mux2_1
Xfanout427 _08494_/Y vssd1 vssd1 vccd1 vccd1 _13123_/B sky130_fd_sc_hd__buf_12
XFILLER_59_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout449 _10710_/S vssd1 vssd1 vccd1 vccd1 _10650_/S sky130_fd_sc_hd__buf_12
XFILLER_141_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09753_ _14121_/Q _13341_/A0 _09762_/S vssd1 vssd1 vccd1 vccd1 _14121_/D sky130_fd_sc_hd__mux2_1
X_06965_ _14506_/Q _06713_/Y _14505_/Q _06715_/Y vssd1 vssd1 vccd1 vccd1 _06969_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_39_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08704_ _13451_/Q _08746_/A2 _08750_/A2 _13515_/Q vssd1 vssd1 vccd1 vccd1 _08704_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_104_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09684_ _14055_/Q _13092_/B2 _09695_/S vssd1 vssd1 vccd1 vccd1 _14055_/D sky130_fd_sc_hd__mux2_1
X_06896_ _15370_/Q _06752_/Y _15369_/Q _06755_/Y _06895_/X vssd1 vssd1 vccd1 vccd1
+ _06896_/X sky130_fd_sc_hd__a221o_1
XFILLER_27_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_620 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08635_ _13461_/Q _08684_/A2 _08683_/A2 _13525_/Q _08634_/X vssd1 vssd1 vccd1 vccd1
+ _08635_/X sky130_fd_sc_hd__a221o_1
XFILLER_82_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08566_ _08722_/A _08566_/B _08566_/C vssd1 vssd1 vccd1 vccd1 _08566_/X sky130_fd_sc_hd__or3_1
XTAP_1429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07517_ _14747_/Q _13426_/Q _07529_/S vssd1 vssd1 vccd1 vccd1 _13426_/D sky130_fd_sc_hd__mux2_1
XFILLER_120_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08497_ _08497_/A _13123_/B vssd1 vssd1 vccd1 vccd1 _08538_/A sky130_fd_sc_hd__nand2_8
XFILLER_120_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_167_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_403 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07448_ _14752_/Q _07447_/X _07480_/S vssd1 vssd1 vccd1 vccd1 _07448_/X sky130_fd_sc_hd__mux2_8
XFILLER_156_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07379_ _13650_/Q _07499_/A2 _07499_/B1 _14678_/Q _07378_/X vssd1 vssd1 vccd1 vccd1
+ _07379_/X sky130_fd_sc_hd__a221o_1
XFILLER_109_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09118_ _14367_/Q _15183_/Q _13822_/Q _14561_/Q _09225_/S0 _09429_/S1 vssd1 vssd1
+ vccd1 vccd1 _09119_/B sky130_fd_sc_hd__mux4_1
XFILLER_13_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10390_ _10390_/A _10390_/B _10390_/C vssd1 vssd1 vccd1 vccd1 _10558_/A sky130_fd_sc_hd__or3_4
XFILLER_135_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09049_ _09406_/S1 _09047_/X _09048_/X vssd1 vssd1 vccd1 vccd1 _09049_/X sky130_fd_sc_hd__a21o_1
XFILLER_159_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12060_ _14010_/Q _13978_/Q _12246_/S vssd1 vssd1 vccd1 vccd1 _12061_/B sky130_fd_sc_hd__mux2_1
XFILLER_145_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_225_clk clkbuf_5_7_0_clk/X vssd1 vssd1 vccd1 vccd1 _15673_/CLK sky130_fd_sc_hd__clkbuf_16
X_11011_ _13251_/A _11356_/C vssd1 vssd1 vccd1 vccd1 _11011_/Y sky130_fd_sc_hd__nor2_1
XFILLER_1_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12962_ _15467_/Q _13119_/S _13116_/C _12961_/X vssd1 vssd1 vccd1 vccd1 _15467_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_86_992 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14701_ _14774_/CLK _14701_/D vssd1 vssd1 vccd1 vccd1 _14701_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11913_ _14357_/Q _15173_/Q _13812_/Q _14551_/Q _12522_/S _12521_/A vssd1 vssd1 vccd1
+ vccd1 _11913_/X sky130_fd_sc_hd__mux4_1
XTAP_4099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12893_ _15421_/Q _15606_/Q _12927_/S vssd1 vssd1 vccd1 vccd1 _15421_/D sky130_fd_sc_hd__mux2_1
XTAP_3365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1088 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14632_ _15453_/CLK _14632_/D vssd1 vssd1 vccd1 vccd1 _14632_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11844_ _15266_/Q _11877_/A1 _11849_/S vssd1 vssd1 vccd1 vccd1 _15266_/D sky130_fd_sc_hd__mux2_1
XTAP_2664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14563_ _15218_/CLK _14563_/D vssd1 vssd1 vccd1 vccd1 _14563_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11775_ _13350_/A0 _15203_/Q _11775_/S vssd1 vssd1 vccd1 vccd1 _15203_/D sky130_fd_sc_hd__mux2_1
XFILLER_60_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13514_ _15374_/CLK _13514_/D vssd1 vssd1 vccd1 vccd1 _13514_/Q sky130_fd_sc_hd__dfxtp_1
X_10726_ _15583_/Q _10731_/B vssd1 vssd1 vccd1 vccd1 _10726_/X sky130_fd_sc_hd__and2_1
X_14494_ _15377_/CLK _14494_/D vssd1 vssd1 vccd1 vccd1 _14494_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13445_ _15543_/CLK _13445_/D vssd1 vssd1 vccd1 vccd1 _13445_/Q sky130_fd_sc_hd__dfxtp_2
X_10657_ _15010_/Q _10569_/B _10652_/B _15027_/Q _10732_/C1 vssd1 vssd1 vccd1 vccd1
+ _10657_/X sky130_fd_sc_hd__a221o_1
XFILLER_103_1020 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13376_ _14479_/Q vssd1 vssd1 vccd1 vccd1 _14479_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_186_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_952 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10588_ _13715_/Q _10602_/B _10587_/X vssd1 vssd1 vccd1 vccd1 _10588_/X sky130_fd_sc_hd__a21o_1
XFILLER_138_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12327_ _14375_/Q _15191_/Q _13830_/Q _14569_/Q _12543_/S _12544_/A vssd1 vssd1 vccd1
+ vccd1 _12327_/X sky130_fd_sc_hd__mux4_1
X_15115_ _15656_/CLK _15115_/D vssd1 vssd1 vccd1 vccd1 _15115_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15046_ _15046_/CLK _15046_/D vssd1 vssd1 vccd1 vccd1 _15046_/Q sky130_fd_sc_hd__dfxtp_4
X_12258_ _14372_/Q _15188_/Q _13827_/Q _14566_/Q _11993_/S _11992_/A vssd1 vssd1 vccd1
+ vccd1 _12258_/X sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_216_clk clkbuf_5_18_0_clk/X vssd1 vssd1 vccd1 vccd1 _15527_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_96_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11209_ _10555_/A _14998_/Q _11237_/S vssd1 vssd1 vccd1 vccd1 _14998_/D sky130_fd_sc_hd__mux2_1
X_12189_ _14369_/Q _15185_/Q _13824_/Q _14563_/Q _12472_/S _12498_/A vssd1 vssd1 vccd1
+ vccd1 _12189_/X sky130_fd_sc_hd__mux4_1
XFILLER_68_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_801 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06750_ _14488_/Q vssd1 vssd1 vccd1 vccd1 _06750_/Y sky130_fd_sc_hd__inv_2
XFILLER_48_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_1076 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06681_ _14909_/Q vssd1 vssd1 vccd1 vccd1 _06681_/Y sky130_fd_sc_hd__inv_2
X_08420_ _14595_/Q _13138_/S _08390_/A _08419_/X vssd1 vssd1 vccd1 vccd1 _13742_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_52_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08351_ _11025_/A _11449_/A vssd1 vssd1 vccd1 vccd1 _08355_/A sky130_fd_sc_hd__nor2_1
XFILLER_177_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07302_ _15315_/Q _15471_/Q _07340_/S vssd1 vssd1 vccd1 vccd1 _07302_/X sky130_fd_sc_hd__mux2_8
X_08282_ _10403_/A _08281_/X _11047_/B vssd1 vssd1 vccd1 vccd1 _08282_/X sky130_fd_sc_hd__mux2_2
XFILLER_165_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07233_ _07233_/A vssd1 vssd1 vccd1 vccd1 _07235_/A sky130_fd_sc_hd__inv_2
XFILLER_177_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_227 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07164_ _15338_/Q _15045_/Q _07193_/S vssd1 vssd1 vccd1 vccd1 _07164_/X sky130_fd_sc_hd__mux2_8
XFILLER_117_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07095_ _07094_/X _14764_/Q _07098_/S vssd1 vssd1 vccd1 vccd1 _13610_/D sky130_fd_sc_hd__mux2_1
XFILLER_59_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_207_clk clkbuf_5_16_0_clk/X vssd1 vssd1 vccd1 vccd1 _15679_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_8_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout202 _09763_/Y vssd1 vssd1 vccd1 vccd1 _09795_/S sky130_fd_sc_hd__buf_12
XFILLER_99_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout213 _09562_/Y vssd1 vssd1 vccd1 vccd1 _09589_/S sky130_fd_sc_hd__buf_12
Xfanout224 _07907_/Y vssd1 vssd1 vccd1 vccd1 _08012_/A2 sky130_fd_sc_hd__clkbuf_16
Xfanout235 _07535_/S vssd1 vssd1 vccd1 vccd1 _07529_/S sky130_fd_sc_hd__buf_12
XFILLER_141_691 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout246 _08531_/Y vssd1 vssd1 vccd1 vccd1 _08747_/B1 sky130_fd_sc_hd__buf_12
XFILLER_113_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout257 _07830_/A vssd1 vssd1 vccd1 vccd1 _07874_/A sky130_fd_sc_hd__buf_8
X_09805_ _14171_/Q _13327_/A0 _09823_/S vssd1 vssd1 vccd1 vccd1 _14171_/D sky130_fd_sc_hd__mux2_1
Xfanout268 _08524_/Y vssd1 vssd1 vccd1 vccd1 _08691_/A2 sky130_fd_sc_hd__clkbuf_16
XFILLER_115_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07997_ _08006_/D _07996_/Y _07971_/A vssd1 vssd1 vccd1 vccd1 _07997_/Y sky130_fd_sc_hd__o21ai_1
Xfanout279 _08724_/B vssd1 vssd1 vccd1 vccd1 _09536_/A2 sky130_fd_sc_hd__buf_12
XFILLER_74_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09736_ _14104_/Q _13324_/A0 _09762_/S vssd1 vssd1 vccd1 vccd1 _14104_/D sky130_fd_sc_hd__mux2_1
X_06948_ _06756_/Y _14486_/Q _13478_/Q _06753_/Y vssd1 vssd1 vccd1 vccd1 _06948_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_28_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09667_ _14038_/Q _11680_/A0 _09690_/S vssd1 vssd1 vccd1 vccd1 _14038_/D sky130_fd_sc_hd__mux2_1
X_06879_ _06879_/A _06879_/B _06879_/C vssd1 vssd1 vccd1 vccd1 _06879_/Y sky130_fd_sc_hd__nand3_1
XFILLER_54_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08618_ _14505_/Q _08748_/B1 _08616_/X _08617_/X vssd1 vssd1 vccd1 vccd1 _08619_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_27_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09598_ _13972_/Q _11853_/A1 _09628_/S vssd1 vssd1 vccd1 vccd1 _13972_/D sky130_fd_sc_hd__mux2_1
XTAP_1237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08549_ _15397_/Q _08748_/A2 _08736_/A2 _13442_/Q vssd1 vssd1 vccd1 vccd1 _08549_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_70_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11560_ _11569_/B _13218_/A _11569_/D _13236_/A vssd1 vssd1 vccd1 vccd1 _11561_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_24_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10511_ _13218_/A _13217_/B vssd1 vssd1 vccd1 vccd1 _10511_/Y sky130_fd_sc_hd__nand2_1
XFILLER_7_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11491_ _13202_/B _11491_/B _11491_/C vssd1 vssd1 vccd1 vccd1 _11502_/B sky130_fd_sc_hd__and3_1
XFILLER_155_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13230_ _13229_/A _10532_/B _13241_/A2 _13229_/Y vssd1 vssd1 vccd1 vccd1 _13230_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_7_749 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10442_ _10443_/B vssd1 vssd1 vccd1 vccd1 _10442_/Y sky130_fd_sc_hd__inv_2
XFILLER_137_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13161_ _11356_/B _13159_/Y _13160_/X _13252_/B _15554_/Q vssd1 vssd1 vccd1 vccd1
+ _15554_/D sky130_fd_sc_hd__a32o_1
XFILLER_151_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10373_ _14767_/Q _13795_/Q _13763_/Q _14766_/Q vssd1 vssd1 vccd1 vccd1 _10373_/X
+ sky130_fd_sc_hd__a22o_2
XFILLER_151_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12112_ _12273_/A1 _12111_/X _12110_/X _12503_/C1 vssd1 vssd1 vccd1 vccd1 _12113_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_2_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13092_ _13005_/X _13118_/A2 _13114_/B1 _13092_/B2 vssd1 vssd1 vccd1 vccd1 _13092_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_3_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12043_ _12595_/A1 _12042_/X _12041_/X _12618_/C1 vssd1 vssd1 vccd1 vccd1 _12044_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_120_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_84 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_96 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13994_ _15335_/CLK _13994_/D vssd1 vssd1 vccd1 vccd1 _13994_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12945_ _13024_/B2 _12937_/X _13024_/A2 _07376_/X vssd1 vssd1 vccd1 vccd1 _12945_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_3162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15664_ _15664_/CLK _15664_/D vssd1 vssd1 vccd1 vccd1 _15664_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12876_ _15404_/Q _15589_/Q _12900_/S vssd1 vssd1 vccd1 vccd1 _15404_/D sky130_fd_sc_hd__mux2_1
XTAP_2472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14615_ _15619_/CLK _14615_/D vssd1 vssd1 vccd1 vccd1 _14615_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11827_ _15249_/Q _11860_/A1 _11849_/S vssd1 vssd1 vccd1 vccd1 _15249_/D sky130_fd_sc_hd__mux2_1
XTAP_2494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15595_ _15599_/CLK _15595_/D vssd1 vssd1 vccd1 vccd1 _15595_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14546_ _15259_/CLK _14546_/D vssd1 vssd1 vccd1 vccd1 _14546_/Q sky130_fd_sc_hd__dfxtp_1
X_11758_ _13080_/B2 _15186_/Q _11774_/S vssd1 vssd1 vccd1 vccd1 _15186_/D sky130_fd_sc_hd__mux2_1
XFILLER_119_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10709_ _15069_/Q _10714_/A2 _10706_/X _10708_/X vssd1 vssd1 vccd1 vccd1 _10709_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_186_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11689_ _11689_/A0 _15120_/Q _11703_/S vssd1 vssd1 vccd1 vccd1 _15120_/D sky130_fd_sc_hd__mux2_1
X_14477_ _15523_/CLK _14477_/D vssd1 vssd1 vccd1 vccd1 _14477_/Q sky130_fd_sc_hd__dfxtp_1
X_13428_ _15381_/CLK _13428_/D vssd1 vssd1 vccd1 vccd1 _13428_/Q sky130_fd_sc_hd__dfxtp_2
X_13359_ _14462_/Q vssd1 vssd1 vccd1 vccd1 _14462_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_170_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_742 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07920_ _14737_/Q _08012_/A2 _07919_/X _08084_/C1 vssd1 vssd1 vccd1 vccd1 _13544_/D
+ sky130_fd_sc_hd__o211a_1
X_15029_ _15041_/CLK _15029_/D vssd1 vssd1 vccd1 vccd1 _15029_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_25_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07851_ _13527_/Q _07858_/D vssd1 vssd1 vccd1 vccd1 _07855_/B sky130_fd_sc_hd__nand2_1
XFILLER_111_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06802_ _06663_/Y _08405_/A _12559_/A _13731_/Q vssd1 vssd1 vccd1 vccd1 _06802_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_96_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput2 ext_read_data[10] vssd1 vssd1 vccd1 vccd1 input2/X sky130_fd_sc_hd__buf_6
X_07782_ _07783_/A _07783_/C vssd1 vssd1 vccd1 vccd1 _08074_/B sky130_fd_sc_hd__nor2_4
XFILLER_83_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09521_ _14033_/Q _14001_/Q _09521_/S vssd1 vssd1 vccd1 vccd1 _09521_/X sky130_fd_sc_hd__mux2_1
XFILLER_65_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06733_ _13455_/Q vssd1 vssd1 vccd1 vccd1 _06733_/Y sky130_fd_sc_hd__inv_2
XFILLER_36_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09452_ _13933_/Q _09451_/X _12481_/A vssd1 vssd1 vccd1 vccd1 _13933_/D sky130_fd_sc_hd__mux2_1
X_06664_ _13730_/Q vssd1 vssd1 vccd1 vccd1 _06664_/Y sky130_fd_sc_hd__inv_2
XFILLER_51_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08403_ _13735_/Q _13138_/S _08390_/B _08402_/X vssd1 vssd1 vccd1 vccd1 _13735_/D
+ sky130_fd_sc_hd__o22a_1
X_09383_ _14541_/Q _14154_/Q _14186_/Q _14122_/Q _09535_/S _08494_/B vssd1 vssd1 vccd1
+ vccd1 _09383_/X sky130_fd_sc_hd__mux4_1
X_08334_ _10507_/A1 _13764_/Q _15408_/Q _10515_/B2 vssd1 vssd1 vccd1 vccd1 _08334_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_177_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08265_ _11349_/B _13162_/B _08262_/Y vssd1 vssd1 vccd1 vccd1 _08266_/A sky130_fd_sc_hd__o21a_2
XFILLER_177_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07216_ _07202_/X _07204_/Y _07213_/X _07215_/Y vssd1 vssd1 vccd1 vccd1 _07230_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_119_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08196_ _13687_/Q _11858_/A1 _08221_/S vssd1 vssd1 vccd1 vccd1 _13687_/D sky130_fd_sc_hd__mux2_1
XFILLER_118_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07147_ _14837_/Q _07104_/X _07146_/X _07131_/A vssd1 vssd1 vccd1 vccd1 _07147_/X
+ sky130_fd_sc_hd__a22o_4
XFILLER_134_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_1087 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07078_ _14638_/Q _14670_/Q _07078_/S vssd1 vssd1 vccd1 vccd1 _07078_/X sky130_fd_sc_hd__mux2_2
XFILLER_133_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09719_ _13341_/A0 _14089_/Q _09728_/S vssd1 vssd1 vccd1 vccd1 _14089_/D sky130_fd_sc_hd__mux2_1
X_10991_ _10991_/A _10991_/B vssd1 vssd1 vccd1 vccd1 _10991_/Y sky130_fd_sc_hd__nor2_1
XFILLER_43_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12730_ _15352_/Q _12765_/B _12729_/X _12809_/C1 vssd1 vssd1 vccd1 vccd1 _15352_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12661_ _13587_/Q _12660_/X _12785_/B vssd1 vssd1 vccd1 vccd1 _12661_/X sky130_fd_sc_hd__mux2_1
XTAP_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_166 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11612_ wire360/X _11612_/B vssd1 vssd1 vccd1 vccd1 _11613_/B sky130_fd_sc_hd__xor2_1
XTAP_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14400_ _15133_/CLK _14400_/D vssd1 vssd1 vccd1 vccd1 _14400_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_187_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15380_ _15381_/CLK _15380_/D vssd1 vssd1 vccd1 vccd1 _15380_/Q sky130_fd_sc_hd__dfxtp_1
X_12592_ _12592_/A1 _12591_/X _06670_/A vssd1 vssd1 vccd1 vccd1 _12592_/X sky130_fd_sc_hd__a21o_1
XFILLER_23_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11543_ _11531_/A _11533_/B _11530_/X vssd1 vssd1 vccd1 vccd1 _11543_/Y sky130_fd_sc_hd__a21oi_1
X_14331_ _15663_/CLK _14331_/D vssd1 vssd1 vccd1 vccd1 _14331_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_184_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_156_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14262_ _14537_/CLK _14262_/D vssd1 vssd1 vccd1 vccd1 _14262_/Q sky130_fd_sc_hd__dfxtp_1
X_11474_ _11473_/Y _15056_/Q _11474_/S vssd1 vssd1 vccd1 vccd1 _15056_/D sky130_fd_sc_hd__mux2_1
X_13213_ _15571_/Q _13214_/B _13211_/Y _13212_/X vssd1 vssd1 vccd1 vccd1 _15571_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_183_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10425_ _07225_/A _10457_/A2 _10424_/X vssd1 vssd1 vccd1 vccd1 _11632_/A sky130_fd_sc_hd__a21o_4
X_14193_ _14420_/CLK _14193_/D vssd1 vssd1 vccd1 vccd1 _14193_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_124_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13144_ _13144_/A0 _15542_/Q _13154_/S vssd1 vssd1 vccd1 vccd1 _15542_/D sky130_fd_sc_hd__mux2_1
X_10356_ _10356_/A _10356_/B vssd1 vssd1 vccd1 vccd1 _10366_/A sky130_fd_sc_hd__and2_1
XFILLER_151_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13075_ _15505_/Q _13081_/A2 _13105_/B1 _13074_/X vssd1 vssd1 vccd1 vccd1 _15505_/D
+ sky130_fd_sc_hd__a22o_1
X_10287_ _14672_/Q _14825_/Q _10715_/S vssd1 vssd1 vccd1 vccd1 _14672_/D sky130_fd_sc_hd__mux2_1
XFILLER_140_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12026_ _15114_/Q _15082_/Q _15655_/Q _13389_/Q _12545_/S _12590_/A vssd1 vssd1 vccd1
+ vccd1 _12026_/X sky130_fd_sc_hd__mux4_1
XFILLER_111_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_918 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13977_ _14572_/CLK _13977_/D vssd1 vssd1 vccd1 vccd1 _13977_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12928_ _15456_/Q _15642_/Q _12928_/S vssd1 vssd1 vccd1 vccd1 _15456_/D sky130_fd_sc_hd__mux2_1
XFILLER_34_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_179_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15647_ _15647_/CLK _15647_/D vssd1 vssd1 vccd1 vccd1 _15647_/Q sky130_fd_sc_hd__dfxtp_1
X_12859_ _14753_/Q _15387_/Q _12866_/S vssd1 vssd1 vccd1 vccd1 _15387_/D sky130_fd_sc_hd__mux2_1
XTAP_2291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15578_ _15579_/CLK _15578_/D vssd1 vssd1 vccd1 vccd1 _15578_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14529_ _15253_/CLK _14529_/D vssd1 vssd1 vccd1 vccd1 _14529_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08050_ _14743_/Q _13621_/Q _08066_/S vssd1 vssd1 vccd1 vccd1 _13621_/D sky130_fd_sc_hd__mux2_1
XFILLER_147_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07001_ _14720_/Q _14719_/Q vssd1 vssd1 vccd1 vccd1 _08027_/A sky130_fd_sc_hd__or2_4
XFILLER_127_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08952_ _09391_/A _08952_/B vssd1 vssd1 vccd1 vccd1 _08952_/X sky130_fd_sc_hd__or2_1
XFILLER_130_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07903_ _07903_/A _07903_/B vssd1 vssd1 vccd1 vccd1 _07903_/Y sky130_fd_sc_hd__nand2_1
XFILLER_130_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08883_ _13904_/Q _11881_/A1 _08885_/S vssd1 vssd1 vccd1 vccd1 _13904_/D sky130_fd_sc_hd__mux2_1
X_07834_ _07837_/B _07833_/Y _07830_/A vssd1 vssd1 vccd1 vccd1 _07834_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_56_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07765_ _13505_/Q _13504_/Q _07765_/C vssd1 vssd1 vccd1 vccd1 _07769_/B sky130_fd_sc_hd__and3_1
XFILLER_72_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06716_ _14504_/Q vssd1 vssd1 vccd1 vccd1 _06716_/Y sky130_fd_sc_hd__inv_2
X_09504_ _13968_/Q _13710_/Q _09535_/S vssd1 vssd1 vccd1 vccd1 _09504_/X sky130_fd_sc_hd__mux2_1
X_07696_ _14743_/Q _07713_/A _07695_/Y _07949_/C1 vssd1 vssd1 vccd1 vccd1 _13486_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_53_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09435_ _09435_/A _09435_/B vssd1 vssd1 vccd1 vccd1 _09435_/X sky130_fd_sc_hd__or2_1
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_1020 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09366_ _09524_/A _09359_/X _09362_/X _08501_/A vssd1 vssd1 vccd1 vccd1 _09366_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_40_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08317_ _11356_/C _11399_/A _10999_/B _11088_/S vssd1 vssd1 vccd1 vccd1 _08317_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_162_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09297_ _08519_/A _09295_/X _09296_/X vssd1 vssd1 vccd1 vccd1 _09297_/X sky130_fd_sc_hd__a21o_1
XANTENNA_40 input12/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_51 _07179_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_62 _07171_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_73 _07149_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08248_ _11356_/B _10551_/A vssd1 vssd1 vccd1 vccd1 _10403_/A sky130_fd_sc_hd__nor2_2
XANTENNA_84 _07103_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_181_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_95 _08638_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_772 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08179_ _08133_/S input21/X _08185_/A vssd1 vssd1 vccd1 vccd1 _08179_/X sky130_fd_sc_hd__and3b_1
XFILLER_137_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10210_ input4/X _14595_/Q _13284_/S vssd1 vssd1 vccd1 vccd1 _14595_/D sky130_fd_sc_hd__mux2_1
X_11190_ _14987_/Q _11164_/S _11170_/X _11189_/Y vssd1 vssd1 vccd1 vccd1 _14987_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_137_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10141_ _14526_/Q _13327_/A0 _10159_/S vssd1 vssd1 vccd1 vccd1 _14526_/D sky130_fd_sc_hd__mux2_1
XFILLER_133_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10072_ _14428_/Q _11858_/A1 _10092_/S vssd1 vssd1 vccd1 vccd1 _14428_/D sky130_fd_sc_hd__mux2_1
XFILLER_94_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13900_ _14415_/CLK _13900_/D vssd1 vssd1 vccd1 vccd1 _13900_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_130_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14880_ _15452_/CLK _14880_/D vssd1 vssd1 vccd1 vccd1 _14880_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13831_ _15293_/CLK _13831_/D vssd1 vssd1 vccd1 vccd1 _13831_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_46_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10974_ _11025_/A _11563_/A vssd1 vssd1 vccd1 vccd1 _11305_/B sky130_fd_sc_hd__nand2_1
X_13762_ _14888_/CLK _13762_/D vssd1 vssd1 vccd1 vccd1 _13762_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_46_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15501_ _15501_/CLK _15501_/D vssd1 vssd1 vccd1 vccd1 _15501_/Q sky130_fd_sc_hd__dfxtp_1
X_12713_ _13594_/Q _12712_/X _12785_/B vssd1 vssd1 vccd1 vccd1 _12713_/X sky130_fd_sc_hd__mux2_1
XFILLER_16_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13693_ _15233_/CLK _13693_/D vssd1 vssd1 vccd1 vccd1 _13693_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15432_ _15618_/CLK _15432_/D vssd1 vssd1 vccd1 vccd1 _15432_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12644_ _15341_/Q _12644_/B vssd1 vssd1 vccd1 vccd1 _12645_/B sky130_fd_sc_hd__nor2_1
X_15363_ _15452_/CLK _15363_/D vssd1 vssd1 vccd1 vccd1 _15363_/Q sky130_fd_sc_hd__dfxtp_2
X_12575_ _14258_/Q _14290_/Q _14322_/Q _14354_/Q _12430_/S _12563_/A vssd1 vssd1 vccd1
+ vccd1 _12575_/X sky130_fd_sc_hd__mux4_1
XFILLER_11_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14314_ _14572_/CLK _14314_/D vssd1 vssd1 vccd1 vccd1 _14314_/Q sky130_fd_sc_hd__dfxtp_1
X_11526_ _11544_/A _11526_/B vssd1 vssd1 vccd1 vccd1 _11526_/Y sky130_fd_sc_hd__xnor2_1
X_15294_ _15300_/CLK _15294_/D vssd1 vssd1 vccd1 vccd1 _15294_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11457_ _11457_/A _11457_/B vssd1 vssd1 vccd1 vccd1 _11458_/B sky130_fd_sc_hd__and2_1
X_14245_ _14439_/CLK _14245_/D vssd1 vssd1 vccd1 vccd1 _14245_/Q sky130_fd_sc_hd__dfxtp_1
X_10408_ _11380_/A _11383_/A _10406_/X _10410_/B vssd1 vssd1 vccd1 vccd1 _10408_/Y
+ sky130_fd_sc_hd__o211ai_1
X_14176_ _15662_/CLK _14176_/D vssd1 vssd1 vccd1 vccd1 _14176_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_178_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11388_ _11389_/B _11389_/C _11414_/D vssd1 vssd1 vccd1 vccd1 _11390_/B sky130_fd_sc_hd__a21bo_1
XFILLER_152_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13127_ _14610_/Q _14609_/Q _13127_/C _14608_/Q vssd1 vssd1 vccd1 vccd1 _13127_/X
+ sky130_fd_sc_hd__or4b_1
X_10339_ _14724_/Q _14917_/Q _10343_/S vssd1 vssd1 vccd1 vccd1 _14724_/D sky130_fd_sc_hd__mux2_1
XFILLER_139_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13058_ _12954_/X _13104_/A2 _13104_/B1 _07388_/X vssd1 vssd1 vccd1 vccd1 _13058_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_97_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12009_ _12595_/A1 _12004_/X _12007_/X _12008_/X _08405_/D vssd1 vssd1 vccd1 vccd1
+ _12021_/B sky130_fd_sc_hd__a221o_1
XFILLER_79_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_1020 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07550_ _07559_/D _07549_/Y _07644_/A vssd1 vssd1 vccd1 vccd1 _07550_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_185_1050 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07481_ _13345_/A0 _13409_/Q _07481_/S vssd1 vssd1 vccd1 vccd1 _13409_/D sky130_fd_sc_hd__mux2_1
XFILLER_146_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09220_ _14372_/Q _15188_/Q _13827_/Q _14566_/Q _09132_/S _09225_/S1 vssd1 vssd1
+ vccd1 vccd1 _09221_/B sky130_fd_sc_hd__mux4_1
XFILLER_21_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09151_ _13887_/Q _09445_/A2 _09522_/B1 _14402_/Q _09437_/A1 vssd1 vssd1 vccd1 vccd1
+ _09151_/X sky130_fd_sc_hd__a221o_1
XFILLER_159_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_642 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08102_ input23/X input2/X input10/X input19/X _08094_/S _07104_/C vssd1 vssd1 vccd1
+ vccd1 _08102_/X sky130_fd_sc_hd__mux4_1
X_09082_ _09437_/A1 _09081_/X _09080_/X _09130_/A vssd1 vssd1 vccd1 vccd1 _09082_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_174_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08033_ _08037_/C _08033_/B vssd1 vssd1 vccd1 vccd1 _08039_/S sky130_fd_sc_hd__nor2_4
XFILLER_135_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09984_ _11838_/A1 _14343_/Q _09996_/S vssd1 vssd1 vccd1 vccd1 _14343_/D sky130_fd_sc_hd__mux2_1
XFILLER_107_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08935_ _14456_/Q _09558_/A2 _08934_/X _13049_/A1 vssd1 vssd1 vccd1 vccd1 _08935_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_76_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08866_ _13887_/Q _11689_/A0 _08880_/S vssd1 vssd1 vccd1 vccd1 _13887_/D sky130_fd_sc_hd__mux2_1
XTAP_3706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07817_ _14742_/Q _07903_/A _07816_/Y _07938_/C1 vssd1 vssd1 vccd1 vccd1 _13517_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_123_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08797_ _13331_/A0 _13823_/Q _08811_/S vssd1 vssd1 vccd1 vccd1 _13823_/D sky130_fd_sc_hd__mux2_1
XFILLER_45_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07748_ _14757_/Q _07750_/A _07747_/Y _08002_/C1 vssd1 vssd1 vccd1 vccd1 _13500_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_53_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07679_ _13482_/Q _13481_/Q _07679_/C vssd1 vssd1 vccd1 vccd1 _07687_/C sky130_fd_sc_hd__and3_2
XFILLER_73_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_103 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09418_ _13868_/Q _14221_/Q _09444_/S vssd1 vssd1 vccd1 vccd1 _09418_/X sky130_fd_sc_hd__mux2_1
X_10690_ _14756_/Q _10689_/X _10715_/S vssd1 vssd1 vccd1 vccd1 _14756_/D sky130_fd_sc_hd__mux2_1
XFILLER_179_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09349_ _09532_/A _09349_/B vssd1 vssd1 vccd1 vccd1 _09349_/X sky130_fd_sc_hd__or2_1
XFILLER_40_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12360_ _12540_/A _12360_/B vssd1 vssd1 vccd1 vccd1 _12360_/X sky130_fd_sc_hd__and2_1
XFILLER_120_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11311_ _11347_/A _11311_/B vssd1 vssd1 vccd1 vccd1 _11311_/Y sky130_fd_sc_hd__nand2_1
XFILLER_4_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12291_ _12544_/A _12291_/B vssd1 vssd1 vccd1 vccd1 _12291_/X sky130_fd_sc_hd__and2_1
XFILLER_4_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_335 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14030_ _15334_/CLK _14030_/D vssd1 vssd1 vccd1 vccd1 _14030_/Q sky130_fd_sc_hd__dfxtp_1
X_11242_ _11242_/A _11242_/B vssd1 vssd1 vccd1 vccd1 _11242_/Y sky130_fd_sc_hd__nor2_1
XFILLER_107_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_1067 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_892 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11173_ _11414_/A _11032_/X _11170_/X vssd1 vssd1 vccd1 vccd1 _11173_/X sky130_fd_sc_hd__a21o_1
XFILLER_171_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_147 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10124_ _14510_/Q _14758_/Q _10124_/S vssd1 vssd1 vccd1 vccd1 _14510_/D sky130_fd_sc_hd__mux2_1
XFILLER_79_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_106 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10055_ _14412_/Q _13341_/A0 _10059_/S vssd1 vssd1 vccd1 vccd1 _14412_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14932_ _15556_/CLK _14932_/D vssd1 vssd1 vccd1 vccd1 _14932_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_76_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14863_ _14863_/CLK _14863_/D vssd1 vssd1 vccd1 vccd1 _14863_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_169_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13814_ _15212_/CLK _13814_/D vssd1 vssd1 vccd1 vccd1 _13814_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14794_ _15647_/CLK _14794_/D vssd1 vssd1 vccd1 vccd1 _14794_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13745_ _14868_/CLK _13745_/D vssd1 vssd1 vccd1 vccd1 _13745_/Q sky130_fd_sc_hd__dfxtp_1
X_10957_ _11023_/A _11584_/A vssd1 vssd1 vccd1 vccd1 _10958_/B sky130_fd_sc_hd__and2_1
XFILLER_31_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13676_ _15645_/CLK _13676_/D vssd1 vssd1 vccd1 vccd1 _13676_/Q sky130_fd_sc_hd__dfxtp_1
X_10888_ _14920_/Q _15551_/Q _12320_/A vssd1 vssd1 vccd1 vccd1 _14920_/D sky130_fd_sc_hd__mux2_1
XFILLER_188_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15415_ _15634_/CLK _15415_/D vssd1 vssd1 vccd1 vccd1 _15415_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_31_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12627_ _12759_/B _12627_/B vssd1 vssd1 vccd1 vccd1 _12627_/Y sky130_fd_sc_hd__nand2_1
XFILLER_185_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15346_ _15453_/CLK _15346_/D vssd1 vssd1 vccd1 vccd1 _15346_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_89_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12558_ _15302_/Q _15270_/Q _15238_/Q _15169_/Q _12568_/S _12567_/A vssd1 vssd1 vccd1
+ vccd1 _12559_/B sky130_fd_sc_hd__mux4_1
XFILLER_106_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11509_ _11508_/X _15059_/Q _11614_/S vssd1 vssd1 vccd1 vccd1 _15059_/D sky130_fd_sc_hd__mux2_1
XFILLER_129_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15277_ _15277_/CLK _15277_/D vssd1 vssd1 vccd1 vccd1 _15277_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12489_ _15299_/Q _15267_/Q _15235_/Q _15166_/Q _12489_/S0 _12489_/S1 vssd1 vssd1
+ vccd1 vccd1 _12490_/B sky130_fd_sc_hd__mux4_1
XFILLER_176_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14228_ _15172_/CLK _14228_/D vssd1 vssd1 vccd1 vccd1 _14228_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_132_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14159_ _15200_/CLK _14159_/D vssd1 vssd1 vccd1 vccd1 _14159_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout609 _12470_/S vssd1 vssd1 vccd1 vccd1 _12246_/S sky130_fd_sc_hd__buf_12
XTAP_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_5_4_0_clk clkbuf_5_5_0_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_5_4_0_clk/X sky130_fd_sc_hd__clkbuf_8
XTAP_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06981_ _13138_/S _08477_/C vssd1 vssd1 vccd1 vccd1 _08777_/A sky130_fd_sc_hd__and2_4
XTAP_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08720_ _13417_/Q _08736_/A2 _08748_/B1 _14490_/Q vssd1 vssd1 vccd1 vccd1 _08720_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08651_ _14500_/Q _08693_/A2 _08649_/X _08650_/X vssd1 vssd1 vccd1 vccd1 _08652_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_27_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07602_ _13461_/Q _07599_/B _13462_/Q vssd1 vssd1 vccd1 vccd1 _07602_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_113_1099 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08582_ _13533_/Q _08750_/A2 _08691_/B1 _13501_/Q _08581_/X vssd1 vssd1 vccd1 vccd1
+ _08582_/X sky130_fd_sc_hd__a221o_1
XFILLER_183_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07533_ _14763_/Q _13442_/Q _07535_/S vssd1 vssd1 vccd1 vccd1 _13442_/D sky130_fd_sc_hd__mux2_1
XFILLER_34_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07464_ _14756_/Q _07463_/X _07480_/S vssd1 vssd1 vccd1 vccd1 _07464_/X sky130_fd_sc_hd__mux2_8
XFILLER_50_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09203_ _14243_/Q _14275_/Q _14307_/Q _14339_/Q _09438_/S0 _09448_/S1 vssd1 vssd1
+ vccd1 vccd1 _09203_/X sky130_fd_sc_hd__mux4_1
X_07395_ _13654_/Q _07499_/A2 _07499_/B1 _14682_/Q _07394_/X vssd1 vssd1 vccd1 vccd1
+ _07395_/X sky130_fd_sc_hd__a221o_1
XFILLER_176_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09134_ _15119_/Q _09536_/A2 _13130_/B1 _15087_/Q _09133_/X vssd1 vssd1 vccd1 vccd1
+ _09134_/X sky130_fd_sc_hd__a221o_1
XFILLER_175_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09065_ _15084_/Q _13130_/B1 _08520_/B _09064_/X vssd1 vssd1 vccd1 vccd1 _09065_/X
+ sky130_fd_sc_hd__a22o_1
X_08016_ _14763_/Q _08022_/B _08015_/Y _08016_/C1 vssd1 vssd1 vccd1 vccd1 _13570_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_135_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xmax_cap371 _08361_/B vssd1 vssd1 vccd1 vccd1 _11457_/A sky130_fd_sc_hd__buf_6
XFILLER_150_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09967_ _13321_/A0 _14326_/Q _09996_/S vssd1 vssd1 vccd1 vccd1 _14326_/D sky130_fd_sc_hd__mux2_1
X_08918_ _14068_/Q _13123_/B _08508_/Y _14036_/Q _09532_/A vssd1 vssd1 vccd1 vccd1
+ _08918_/X sky130_fd_sc_hd__a221o_1
XFILLER_94_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09898_ _11818_/A _09964_/B vssd1 vssd1 vccd1 vccd1 _09898_/Y sky130_fd_sc_hd__nand2b_4
XTAP_3503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08849_ _13872_/Q _13110_/B2 _08851_/S vssd1 vssd1 vccd1 vccd1 _13872_/D sky130_fd_sc_hd__mux2_1
XFILLER_85_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_183 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11860_ _15281_/Q _11860_/A1 _11878_/S vssd1 vssd1 vccd1 vccd1 _15281_/D sky130_fd_sc_hd__mux2_1
XTAP_2824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10811_ _14843_/Q _07284_/A _12900_/S vssd1 vssd1 vccd1 vccd1 _14843_/D sky130_fd_sc_hd__mux2_1
X_11791_ _15214_/Q _11857_/A1 _11817_/S vssd1 vssd1 vccd1 vccd1 _15214_/D sky130_fd_sc_hd__mux2_1
XFILLER_72_378 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13530_ _14506_/CLK _13530_/D vssd1 vssd1 vccd1 vccd1 _13530_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10742_ _15406_/Q _14774_/Q _10764_/S vssd1 vssd1 vccd1 vccd1 _14774_/D sky130_fd_sc_hd__mux2_1
XFILLER_129_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13461_ _13627_/CLK _13461_/D vssd1 vssd1 vccd1 vccd1 _13461_/Q sky130_fd_sc_hd__dfxtp_2
X_10673_ _14981_/Q _10718_/A2 _10722_/B1 _14949_/Q _10672_/X vssd1 vssd1 vccd1 vccd1
+ _10673_/X sky130_fd_sc_hd__a221o_2
XFILLER_9_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15200_ _15200_/CLK _15200_/D vssd1 vssd1 vccd1 vccd1 _15200_/Q sky130_fd_sc_hd__dfxtp_1
X_12412_ _12573_/A _12412_/B _12412_/C vssd1 vssd1 vccd1 vccd1 _12412_/X sky130_fd_sc_hd__and3_1
XFILLER_173_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13392_ _15658_/CLK _13392_/D vssd1 vssd1 vccd1 vccd1 _13392_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15131_ _15328_/CLK _15131_/D vssd1 vssd1 vccd1 vccd1 _15131_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_182_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12343_ _12573_/A _12343_/B _12343_/C vssd1 vssd1 vccd1 vccd1 _12343_/X sky130_fd_sc_hd__and3_2
XFILLER_154_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15062_ _15067_/CLK _15062_/D vssd1 vssd1 vccd1 vccd1 _15062_/Q sky130_fd_sc_hd__dfxtp_4
X_12274_ _12596_/A _12274_/B _12274_/C vssd1 vssd1 vccd1 vccd1 _12274_/X sky130_fd_sc_hd__and3_2
XFILLER_114_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_572 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11225_ _10527_/D _15013_/Q _11232_/S vssd1 vssd1 vccd1 vccd1 _15013_/D sky130_fd_sc_hd__mux2_1
XFILLER_4_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14013_ _15133_/CLK _14013_/D vssd1 vssd1 vccd1 vccd1 _14013_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_122_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11156_ _11347_/A _11156_/B vssd1 vssd1 vccd1 vccd1 _11156_/Y sky130_fd_sc_hd__nand2_1
XFILLER_110_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10107_ _14493_/Q _14741_/Q _10131_/S vssd1 vssd1 vccd1 vccd1 _14493_/D sky130_fd_sc_hd__mux2_1
XFILLER_136_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_371 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11087_ _11041_/Y _11044_/Y _11356_/B vssd1 vssd1 vccd1 vccd1 _11087_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10038_ _14395_/Q _11649_/A0 _10064_/S vssd1 vssd1 vccd1 vccd1 _14395_/D sky130_fd_sc_hd__mux2_1
XFILLER_49_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14915_ _15552_/CLK _14915_/D vssd1 vssd1 vccd1 vccd1 _14915_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14846_ _15510_/CLK _14846_/D vssd1 vssd1 vccd1 vccd1 _14846_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14777_ _15599_/CLK _14777_/D vssd1 vssd1 vccd1 vccd1 _14777_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11989_ _13879_/Q _14394_/Q _11993_/S vssd1 vssd1 vccd1 vccd1 _11989_/X sky130_fd_sc_hd__mux2_1
XFILLER_90_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13728_ _15041_/CLK _13728_/D vssd1 vssd1 vccd1 vccd1 _13728_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13659_ _14774_/CLK _13659_/D vssd1 vssd1 vccd1 vccd1 _13659_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_83_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07180_ _15354_/Q _15061_/Q _07188_/S vssd1 vssd1 vccd1 vccd1 _07180_/X sky130_fd_sc_hd__mux2_8
XFILLER_9_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15329_ _15517_/CLK _15329_/D vssd1 vssd1 vccd1 vccd1 _15329_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout406 _13156_/Y vssd1 vssd1 vccd1 vccd1 _13252_/B sky130_fd_sc_hd__buf_8
Xfanout417 _10894_/X vssd1 vssd1 vccd1 vccd1 _10948_/B sky130_fd_sc_hd__buf_6
X_09821_ _14187_/Q _11876_/A1 _09823_/S vssd1 vssd1 vccd1 vccd1 _14187_/D sky130_fd_sc_hd__mux2_1
XFILLER_98_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout428 _09419_/A2 vssd1 vssd1 vccd1 vccd1 _09449_/A1 sky130_fd_sc_hd__buf_12
Xfanout439 _07499_/B1 vssd1 vssd1 vccd1 vccd1 _07483_/B1 sky130_fd_sc_hd__clkbuf_16
XFILLER_141_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09752_ _14120_/Q _13340_/A0 _09762_/S vssd1 vssd1 vccd1 vccd1 _14120_/D sky130_fd_sc_hd__mux2_1
X_06964_ _06946_/X _06963_/Y _06945_/A vssd1 vssd1 vccd1 vccd1 _06964_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_104_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08703_ _13799_/Q _12932_/S _08698_/X _08702_/X vssd1 vssd1 vccd1 vccd1 _13799_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_55_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09683_ _14054_/Q _11838_/A1 _09695_/S vssd1 vssd1 vccd1 vccd1 _14054_/D sky130_fd_sc_hd__mux2_1
XFILLER_67_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06895_ _15369_/Q _06755_/Y _15368_/Q _06757_/Y vssd1 vssd1 vccd1 vccd1 _06895_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_55_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08634_ _13596_/Q _08691_/A2 _08693_/B1 _13628_/Q vssd1 vssd1 vccd1 vccd1 _08634_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_42_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08565_ _14513_/Q _08748_/B1 _08563_/X _08564_/X vssd1 vssd1 vccd1 vccd1 _08566_/C
+ sky130_fd_sc_hd__a211o_1
X_07516_ _14746_/Q _13425_/Q _07529_/S vssd1 vssd1 vccd1 vccd1 _13425_/D sky130_fd_sc_hd__mux2_1
X_08496_ _08910_/S _13125_/A vssd1 vssd1 vccd1 vccd1 _08724_/B sky130_fd_sc_hd__nor2_8
XFILLER_161_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07447_ _13667_/Q _07483_/A2 _07483_/B1 _14695_/Q _07446_/X vssd1 vssd1 vccd1 vccd1
+ _07447_/X sky130_fd_sc_hd__a221o_1
XFILLER_22_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_170_clk clkbuf_5_23_0_clk/X vssd1 vssd1 vccd1 vccd1 _15544_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_167_247 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_973 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07378_ _14646_/Q _07498_/B _07498_/C vssd1 vssd1 vccd1 vccd1 _07378_/X sky130_fd_sc_hd__and3_1
XFILLER_164_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09117_ _15284_/Q _15252_/Q _15220_/Q _15151_/Q _09225_/S0 _09225_/S1 vssd1 vssd1
+ vccd1 vccd1 _09117_/X sky130_fd_sc_hd__mux4_1
XFILLER_136_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09048_ _13882_/Q _09445_/A2 _09522_/B1 _14397_/Q _09445_/C1 vssd1 vssd1 vccd1 vccd1
+ _09048_/X sky130_fd_sc_hd__a221o_1
XFILLER_164_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11010_ _11259_/S _11312_/A _11324_/B _11007_/X vssd1 vssd1 vccd1 vccd1 _11010_/Y
+ sky130_fd_sc_hd__a31oi_2
XFILLER_131_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_43 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12961_ _13324_/A0 _13039_/A2 _12960_/X _12944_/A vssd1 vssd1 vccd1 vccd1 _12961_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_4056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14700_ _15438_/CLK _14700_/D vssd1 vssd1 vccd1 vccd1 _14700_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11912_ _11908_/X _11909_/X _12617_/S vssd1 vssd1 vccd1 vccd1 _11912_/X sky130_fd_sc_hd__mux2_1
XTAP_3355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15680_ _15680_/CLK _15680_/D vssd1 vssd1 vccd1 vccd1 _15680_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12892_ _15420_/Q _15605_/Q _12929_/S vssd1 vssd1 vccd1 vccd1 _15420_/D sky130_fd_sc_hd__mux2_1
XTAP_2621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14631_ _15354_/CLK _14631_/D vssd1 vssd1 vccd1 vccd1 _14631_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_166_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11843_ _15265_/Q _11876_/A1 _11849_/S vssd1 vssd1 vccd1 vccd1 _15265_/D sky130_fd_sc_hd__mux2_1
XFILLER_54_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14562_ _15184_/CLK _14562_/D vssd1 vssd1 vccd1 vccd1 _14562_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11774_ _11816_/A1 _15202_/Q _11774_/S vssd1 vssd1 vccd1 vccd1 _15202_/D sky130_fd_sc_hd__mux2_1
XTAP_1964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13513_ _15461_/CLK _13513_/D vssd1 vssd1 vccd1 vccd1 _13513_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10725_ _14763_/Q _10724_/X _10735_/S vssd1 vssd1 vccd1 vccd1 _14763_/D sky130_fd_sc_hd__mux2_1
XFILLER_13_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_161_clk clkbuf_5_19_0_clk/X vssd1 vssd1 vccd1 vccd1 _15650_/CLK sky130_fd_sc_hd__clkbuf_16
X_14493_ _14493_/CLK _14493_/D vssd1 vssd1 vccd1 vccd1 _14493_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_186_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13444_ _15461_/CLK _13444_/D vssd1 vssd1 vccd1 vccd1 _13444_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_186_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10656_ _15569_/Q _10706_/B vssd1 vssd1 vccd1 vccd1 _10656_/X sky130_fd_sc_hd__and2_1
XFILLER_16_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_1032 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13375_ _14478_/Q vssd1 vssd1 vccd1 vccd1 _14478_/D sky130_fd_sc_hd__clkbuf_2
X_10587_ _15555_/Q _10731_/B _10733_/B1 _14932_/Q vssd1 vssd1 vccd1 vccd1 _10587_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_10_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15114_ _15679_/CLK _15114_/D vssd1 vssd1 vccd1 vccd1 _15114_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12326_ _12322_/X _12323_/X _12536_/A vssd1 vssd1 vccd1 vccd1 _12326_/X sky130_fd_sc_hd__mux2_1
XFILLER_126_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15045_ _15306_/CLK _15045_/D vssd1 vssd1 vccd1 vccd1 _15045_/Q sky130_fd_sc_hd__dfxtp_4
X_12257_ _12253_/X _12254_/X _12260_/A vssd1 vssd1 vccd1 vccd1 _12257_/X sky130_fd_sc_hd__mux2_1
XFILLER_141_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11208_ _10556_/B _14997_/Q _11237_/S vssd1 vssd1 vccd1 vccd1 _14997_/D sky130_fd_sc_hd__mux2_1
X_12188_ _12184_/X _12185_/X _12490_/A vssd1 vssd1 vccd1 vccd1 _12188_/X sky130_fd_sc_hd__mux2_1
XFILLER_95_201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11139_ _14971_/Q _11138_/Y _11164_/S vssd1 vssd1 vccd1 vccd1 _14971_/D sky130_fd_sc_hd__mux2_1
XFILLER_1_691 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1088 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06680_ _14907_/Q vssd1 vssd1 vccd1 vccd1 _06680_/Y sky130_fd_sc_hd__inv_2
XFILLER_36_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_131 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14829_ _15647_/CLK _14829_/D vssd1 vssd1 vccd1 vccd1 _14829_/Q sky130_fd_sc_hd__dfxtp_1
X_08350_ _13724_/Q _11346_/A2 _11351_/C1 _08349_/X vssd1 vssd1 vccd1 vccd1 _13724_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_51_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07301_ _07301_/A vssd1 vssd1 vccd1 vccd1 _07301_/Y sky130_fd_sc_hd__inv_2
XFILLER_149_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08281_ _08266_/Y _08280_/Y _11088_/S vssd1 vssd1 vccd1 vccd1 _08281_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_152_clk clkbuf_5_24_0_clk/X vssd1 vssd1 vccd1 vccd1 _15617_/CLK sky130_fd_sc_hd__clkbuf_16
X_07232_ _13930_/Q _15517_/Q _15527_/Q vssd1 vssd1 vccd1 vccd1 _07233_/A sky130_fd_sc_hd__mux2_8
XFILLER_165_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_239 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07163_ _07163_/A _07163_/B vssd1 vssd1 vccd1 vccd1 _07163_/X sky130_fd_sc_hd__and2_4
XFILLER_30_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_1059 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07094_ _07093_/X _13610_/Q _12662_/S vssd1 vssd1 vccd1 vccd1 _07094_/X sky130_fd_sc_hd__mux2_1
XFILLER_117_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout203 _09730_/Y vssd1 vssd1 vccd1 vccd1 _09757_/S sky130_fd_sc_hd__buf_12
XFILLER_120_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout214 _09562_/Y vssd1 vssd1 vccd1 vccd1 _09594_/S sky130_fd_sc_hd__buf_12
Xfanout225 _07964_/A vssd1 vssd1 vccd1 vccd1 _07971_/A sky130_fd_sc_hd__buf_6
XFILLER_59_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout236 _07505_/X vssd1 vssd1 vccd1 vccd1 _07535_/S sky130_fd_sc_hd__buf_12
XFILLER_113_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09804_ _14170_/Q _13326_/A0 _09823_/S vssd1 vssd1 vccd1 vccd1 _14170_/D sky130_fd_sc_hd__mux2_1
XFILLER_8_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_523 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout247 _08530_/Y vssd1 vssd1 vccd1 vccd1 _08747_/A2 sky130_fd_sc_hd__buf_12
Xfanout258 _07783_/X vssd1 vssd1 vccd1 vccd1 _07830_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_75_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout269 _08513_/Y vssd1 vssd1 vccd1 vccd1 _08748_/B1 sky130_fd_sc_hd__buf_12
X_07996_ _13564_/Q _13563_/Q _07995_/D _13565_/Q vssd1 vssd1 vccd1 vccd1 _07996_/Y
+ sky130_fd_sc_hd__a31oi_1
XFILLER_28_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09735_ _14103_/Q _13323_/A0 _09757_/S vssd1 vssd1 vccd1 vccd1 _14103_/D sky130_fd_sc_hd__mux2_1
XFILLER_74_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06947_ _06742_/Y _13482_/Q _06745_/Y _13481_/Q _06946_/X vssd1 vssd1 vccd1 vccd1
+ _06947_/X sky130_fd_sc_hd__a221o_1
X_09666_ _14037_/Q _11854_/A1 _09695_/S vssd1 vssd1 vccd1 vccd1 _14037_/D sky130_fd_sc_hd__mux2_1
XFILLER_54_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06878_ _06692_/Y _13506_/Q _14509_/Q _06707_/Y vssd1 vssd1 vccd1 vccd1 _06878_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_83_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08617_ _15387_/Q _08748_/A2 _08736_/A2 _13432_/Q vssd1 vssd1 vccd1 vccd1 _08617_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_1205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_827 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09597_ _13971_/Q _13319_/A0 _09627_/S vssd1 vssd1 vccd1 vccd1 _13971_/D sky130_fd_sc_hd__mux2_1
XTAP_1227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08548_ _13538_/Q _08750_/A2 _08747_/A2 _13570_/Q _08547_/X vssd1 vssd1 vccd1 vccd1
+ _08552_/B sky130_fd_sc_hd__a221o_1
X_08479_ hold8/A _08465_/B _08478_/X _13120_/S vssd1 vssd1 vccd1 vccd1 _08479_/X sky130_fd_sc_hd__a211o_1
Xclkbuf_leaf_143_clk clkbuf_5_28_0_clk/X vssd1 vssd1 vccd1 vccd1 _15399_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_24_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10510_ _13217_/B _13218_/A vssd1 vssd1 vccd1 vccd1 _10512_/B sky130_fd_sc_hd__nand2b_1
X_11490_ _11505_/C _11484_/B _11502_/A vssd1 vssd1 vccd1 vccd1 _11493_/A sky130_fd_sc_hd__a21o_1
XFILLER_168_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_537 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10441_ _11624_/A _11626_/A vssd1 vssd1 vccd1 vccd1 _10443_/B sky130_fd_sc_hd__and2_1
X_10372_ _11431_/A _11436_/B vssd1 vssd1 vccd1 vccd1 _10382_/B sky130_fd_sc_hd__xor2_2
X_13160_ _13251_/A _13159_/B _13219_/S vssd1 vssd1 vccd1 vccd1 _13160_/X sky130_fd_sc_hd__o21a_1
XFILLER_156_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12111_ _12094_/X _12095_/X _12260_/A vssd1 vssd1 vccd1 vccd1 _12111_/X sky130_fd_sc_hd__mux2_1
X_13091_ _15513_/Q _10877_/S _13042_/A _13090_/X vssd1 vssd1 vccd1 vccd1 _15513_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_123_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12042_ _12025_/X _12026_/X _12594_/S vssd1 vssd1 vccd1 vccd1 _12042_/X sky130_fd_sc_hd__mux2_1
XFILLER_85_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13993_ _15654_/CLK _13993_/D vssd1 vssd1 vccd1 vccd1 _13993_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12944_ _12944_/A _13116_/B vssd1 vssd1 vccd1 vccd1 _12944_/Y sky130_fd_sc_hd__nor2_4
XTAP_3141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15663_ _15663_/CLK _15663_/D vssd1 vssd1 vccd1 vccd1 _15663_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_130 _14745_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12875_ _15403_/Q _15588_/Q _12900_/S vssd1 vssd1 vccd1 vccd1 _15403_/D sky130_fd_sc_hd__mux2_1
XTAP_3196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14614_ _14649_/CLK _14614_/D vssd1 vssd1 vccd1 vccd1 _14614_/Q sky130_fd_sc_hd__dfxtp_4
X_11826_ _15248_/Q _12967_/A1 _11849_/S vssd1 vssd1 vccd1 vccd1 _15248_/D sky130_fd_sc_hd__mux2_1
XFILLER_61_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15594_ _15599_/CLK _15594_/D vssd1 vssd1 vccd1 vccd1 _15594_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14545_ _15161_/CLK _14545_/D vssd1 vssd1 vccd1 vccd1 _14545_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_134_clk clkbuf_5_29_0_clk/X vssd1 vssd1 vccd1 vccd1 _14513_/CLK sky130_fd_sc_hd__clkbuf_16
X_11757_ _13332_/A0 _15185_/Q _11774_/S vssd1 vssd1 vccd1 vccd1 _15185_/D sky130_fd_sc_hd__mux2_1
XTAP_1794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10708_ _14988_/Q _10718_/A2 _10722_/B1 _14956_/Q _10707_/X vssd1 vssd1 vccd1 vccd1
+ _10708_/X sky130_fd_sc_hd__a221o_1
XFILLER_159_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14476_ _15081_/CLK _14476_/D vssd1 vssd1 vccd1 vccd1 _14476_/Q sky130_fd_sc_hd__dfxtp_1
X_11688_ _13074_/B2 _15119_/Q _11703_/S vssd1 vssd1 vccd1 vccd1 _15119_/D sky130_fd_sc_hd__mux2_1
X_13427_ _15381_/CLK _13427_/D vssd1 vssd1 vccd1 vccd1 _13427_/Q sky130_fd_sc_hd__dfxtp_2
X_10639_ _15055_/Q _10734_/A2 _10636_/X _10638_/X vssd1 vssd1 vccd1 vccd1 _10639_/X
+ sky130_fd_sc_hd__o22a_2
XFILLER_155_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13358_ _14461_/Q vssd1 vssd1 vccd1 vccd1 _14461_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_142_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12309_ _13957_/Q _13699_/Q _12614_/S vssd1 vssd1 vccd1 vccd1 _12310_/B sky130_fd_sc_hd__mux2_1
XFILLER_114_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13289_ _12645_/Y _15621_/Q _13291_/S vssd1 vssd1 vccd1 vccd1 _15621_/D sky130_fd_sc_hd__mux2_1
XFILLER_46_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15028_ _15041_/CLK _15028_/D vssd1 vssd1 vccd1 vccd1 _15028_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_102_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07850_ _14751_/Q _07874_/A _07849_/Y _07949_/C1 vssd1 vssd1 vccd1 vccd1 _13526_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_57_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06801_ _06663_/Y _08405_/A _12618_/C1 _13729_/Q vssd1 vssd1 vccd1 vccd1 _06801_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_56_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07781_ _08027_/A _14717_/Q _14718_/Q vssd1 vssd1 vccd1 vccd1 _07783_/C sky130_fd_sc_hd__or3b_4
Xinput3 ext_read_data[11] vssd1 vssd1 vccd1 vccd1 input3/X sky130_fd_sc_hd__buf_6
XFILLER_110_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09520_ _09523_/A1 _09518_/X _09519_/X vssd1 vssd1 vccd1 vccd1 _09524_/B sky130_fd_sc_hd__a21o_1
XFILLER_49_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06732_ _13487_/Q vssd1 vssd1 vccd1 vccd1 _06732_/Y sky130_fd_sc_hd__inv_2
XFILLER_36_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09451_ _14607_/Q _09440_/X _09449_/X _09450_/X vssd1 vssd1 vccd1 vccd1 _09451_/X
+ sky130_fd_sc_hd__o22a_1
X_06663_ _13733_/Q vssd1 vssd1 vccd1 vccd1 _06663_/Y sky130_fd_sc_hd__inv_2
XFILLER_149_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08402_ _13140_/S _08469_/A vssd1 vssd1 vccd1 vccd1 _08402_/X sky130_fd_sc_hd__or2_2
XFILLER_101_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09382_ _09382_/A _09382_/B _09382_/C vssd1 vssd1 vccd1 vccd1 _09382_/X sky130_fd_sc_hd__and3_1
XFILLER_178_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08333_ _11025_/A _11431_/A vssd1 vssd1 vccd1 vccd1 _10986_/B sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_125_clk clkbuf_5_31_0_clk/X vssd1 vssd1 vccd1 vccd1 _13632_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_33_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08264_ _07336_/A _10481_/B _08263_/X vssd1 vssd1 vccd1 vccd1 _13162_/B sky130_fd_sc_hd__a21oi_4
XFILLER_178_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07215_ _07215_/A vssd1 vssd1 vccd1 vccd1 _07215_/Y sky130_fd_sc_hd__inv_2
X_08195_ _13686_/Q _11857_/A1 _08221_/S vssd1 vssd1 vccd1 vccd1 _13686_/D sky130_fd_sc_hd__mux2_1
XFILLER_119_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07146_ _14853_/Q _14845_/Q _07146_/S vssd1 vssd1 vccd1 vccd1 _07146_/X sky130_fd_sc_hd__mux2_1
XFILLER_117_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07077_ _07076_/X _14758_/Q _07077_/S vssd1 vssd1 vccd1 vccd1 _13604_/D sky130_fd_sc_hd__mux2_1
XFILLER_69_1099 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07979_ _07981_/B _07978_/X _07971_/A vssd1 vssd1 vccd1 vccd1 _07979_/X sky130_fd_sc_hd__a21bo_1
XFILLER_75_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09718_ _13340_/A0 _14088_/Q _09728_/S vssd1 vssd1 vccd1 vccd1 _14088_/D sky130_fd_sc_hd__mux2_1
XFILLER_132_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10990_ _10990_/A _11242_/B vssd1 vssd1 vccd1 vccd1 _10992_/B sky130_fd_sc_hd__nor2_1
XFILLER_56_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09649_ _14022_/Q _11838_/A1 _09661_/S vssd1 vssd1 vccd1 vccd1 _14022_/D sky130_fd_sc_hd__mux2_1
XTAP_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_1048 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12660_ _15050_/Q _12659_/Y _12834_/B vssd1 vssd1 vccd1 vccd1 _12660_/X sky130_fd_sc_hd__mux2_1
XFILLER_150_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11611_ _11611_/A _11611_/B vssd1 vssd1 vccd1 vccd1 _11613_/A sky130_fd_sc_hd__nor2_1
XTAP_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_116_clk _15447_/CLK vssd1 vssd1 vccd1 vccd1 _15637_/CLK sky130_fd_sc_hd__clkbuf_16
X_12591_ _14097_/Q _14065_/Q _12591_/S vssd1 vssd1 vccd1 vccd1 _12591_/X sky130_fd_sc_hd__mux2_1
X_14330_ _14462_/CLK _14330_/D vssd1 vssd1 vccd1 vccd1 _14330_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_184_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11542_ _11542_/A _11542_/B vssd1 vssd1 vccd1 vccd1 _11576_/A sky130_fd_sc_hd__nand2_1
XFILLER_129_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14261_ _14606_/CLK _14261_/D vssd1 vssd1 vccd1 vccd1 _14261_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_183_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11473_ _11505_/B _11473_/B vssd1 vssd1 vccd1 vccd1 _11473_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_13_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13212_ _13233_/A _11521_/A _13219_/S vssd1 vssd1 vccd1 vccd1 _13212_/X sky130_fd_sc_hd__o21a_1
XFILLER_13_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10424_ _08240_/A _13776_/Q _13744_/Q _08237_/A vssd1 vssd1 vccd1 vccd1 _10424_/X
+ sky130_fd_sc_hd__a22o_1
X_14192_ _15678_/CLK _14192_/D vssd1 vssd1 vccd1 vccd1 _14192_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_152_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13143_ _09342_/S _15541_/Q _13154_/S vssd1 vssd1 vccd1 vccd1 _15541_/D sky130_fd_sc_hd__mux2_1
X_10355_ _13199_/B _11496_/A vssd1 vssd1 vccd1 vccd1 _10356_/B sky130_fd_sc_hd__or2_1
XFILLER_152_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10286_ _14671_/Q _14824_/Q _10630_/S vssd1 vssd1 vccd1 vccd1 _14671_/D sky130_fd_sc_hd__mux2_1
XFILLER_140_938 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13074_ _12978_/X _13104_/A2 _13104_/B1 _13074_/B2 vssd1 vssd1 vccd1 vccd1 _13074_/X
+ sky130_fd_sc_hd__a22o_1
X_12025_ _14524_/Q _14137_/Q _14169_/Q _14105_/Q _12591_/S _12590_/A vssd1 vssd1 vccd1
+ vccd1 _12025_/X sky130_fd_sc_hd__mux4_1
XFILLER_38_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13976_ _15278_/CLK _13976_/D vssd1 vssd1 vccd1 vccd1 _13976_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12927_ hold9/A _15641_/Q _12927_/S vssd1 vssd1 vccd1 vccd1 _15455_/D sky130_fd_sc_hd__mux2_1
XFILLER_34_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_164 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_218 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15646_ _15646_/CLK _15646_/D vssd1 vssd1 vccd1 vccd1 _15646_/Q sky130_fd_sc_hd__dfxtp_1
X_12858_ _14752_/Q _15386_/Q _12871_/S vssd1 vssd1 vccd1 vccd1 _15386_/D sky130_fd_sc_hd__mux2_1
XFILLER_34_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11809_ _15232_/Q _13342_/A0 _11817_/S vssd1 vssd1 vccd1 vccd1 _15232_/D sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_107_clk clkbuf_5_26_0_clk/X vssd1 vssd1 vccd1 vccd1 _15453_/CLK sky130_fd_sc_hd__clkbuf_16
X_15577_ _15577_/CLK _15577_/D vssd1 vssd1 vccd1 vccd1 _15577_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12789_ _15361_/Q _15360_/Q _12789_/C vssd1 vssd1 vccd1 vccd1 _13309_/B sky130_fd_sc_hd__and3_1
XTAP_1591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14528_ _15674_/CLK _14528_/D vssd1 vssd1 vccd1 vccd1 _14528_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_175_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14459_ _15211_/CLK _14459_/D vssd1 vssd1 vccd1 vccd1 _14459_/Q sky130_fd_sc_hd__dfxtp_1
X_07000_ _14724_/Q _07504_/B _10098_/A vssd1 vssd1 vccd1 vccd1 _08074_/A sky130_fd_sc_hd__nor3_4
XFILLER_134_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08951_ _14359_/Q _15175_/Q _13814_/Q _14553_/Q _09230_/S _09234_/S1 vssd1 vssd1
+ vccd1 vccd1 _08952_/B sky130_fd_sc_hd__mux4_1
XFILLER_97_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07902_ _07913_/D _07902_/B vssd1 vssd1 vccd1 vccd1 _07903_/B sky130_fd_sc_hd__nand2b_1
X_08882_ _13903_/Q _13347_/A0 _08885_/S vssd1 vssd1 vccd1 vccd1 _13903_/D sky130_fd_sc_hd__mux2_1
XFILLER_111_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07833_ _13521_/Q _07836_/D _13522_/Q vssd1 vssd1 vccd1 vccd1 _07833_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_57_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07764_ _13505_/Q _07764_/B vssd1 vssd1 vccd1 vccd1 _07764_/Y sky130_fd_sc_hd__nor2_1
XFILLER_112_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09503_ _08668_/D _09499_/X _09502_/X _09498_/X vssd1 vssd1 vccd1 vccd1 _09516_/B
+ sky130_fd_sc_hd__a211o_1
X_06715_ _13496_/Q vssd1 vssd1 vccd1 vccd1 _06715_/Y sky130_fd_sc_hd__inv_2
XFILLER_65_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07695_ _07693_/Y _07697_/B _07713_/A vssd1 vssd1 vccd1 vccd1 _07695_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_52_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_432 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09434_ _14382_/Q _15198_/Q _13837_/Q _14576_/Q _09444_/S _09446_/A1 vssd1 vssd1
+ vccd1 vccd1 _09435_/B sky130_fd_sc_hd__mux4_1
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_988 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09365_ _08519_/B _09363_/X _09364_/X _08668_/D vssd1 vssd1 vccd1 vccd1 _09365_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_36_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08316_ _10986_/A _08316_/B vssd1 vssd1 vccd1 vccd1 _08316_/Y sky130_fd_sc_hd__nor2_1
XFILLER_138_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_30 _14749_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_177_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09296_ _13894_/Q _09522_/A2 _08512_/B _14409_/Q _13123_/A vssd1 vssd1 vccd1 vccd1
+ _09296_/X sky130_fd_sc_hd__a221o_1
XFILLER_165_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_41 input16/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_52 _07188_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_63 _07171_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08247_ _11356_/C _10895_/B vssd1 vssd1 vccd1 vccd1 _10551_/A sky130_fd_sc_hd__nand2_2
XANTENNA_74 _07151_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_85 _07107_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_96 _08991_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08178_ _13676_/Q _10695_/S _08155_/X _08177_/X vssd1 vssd1 vccd1 vccd1 _13676_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_4_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07129_ _07131_/A _07129_/B vssd1 vssd1 vccd1 vccd1 _07129_/X sky130_fd_sc_hd__and2_4
XFILLER_133_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10140_ _14525_/Q _13326_/A0 _10159_/S vssd1 vssd1 vccd1 vccd1 _14525_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10071_ _14427_/Q _11649_/A0 _10097_/S vssd1 vssd1 vccd1 vccd1 _14427_/D sky130_fd_sc_hd__mux2_1
XFILLER_88_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_767 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_88 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13830_ _15292_/CLK _13830_/D vssd1 vssd1 vccd1 vccd1 _13830_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13761_ _14888_/CLK _13761_/D vssd1 vssd1 vccd1 vccd1 _13761_/Q sky130_fd_sc_hd__dfxtp_1
X_10973_ _11330_/A _10971_/Y _10972_/X vssd1 vssd1 vccd1 vccd1 _10973_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_55_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15500_ _15500_/CLK _15500_/D vssd1 vssd1 vccd1 vccd1 _15500_/Q sky130_fd_sc_hd__dfxtp_1
X_12712_ _15057_/Q _12711_/X _12792_/B vssd1 vssd1 vccd1 vccd1 _12712_/X sky130_fd_sc_hd__mux2_1
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13692_ _15285_/CLK _13692_/D vssd1 vssd1 vccd1 vccd1 _13692_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15431_ _15617_/CLK _15431_/D vssd1 vssd1 vccd1 vccd1 _15431_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_30_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12643_ _15341_/Q _12644_/B vssd1 vssd1 vccd1 vccd1 _12657_/C sky130_fd_sc_hd__and2_2
XFILLER_31_638 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_178_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15362_ _15452_/CLK _15362_/D vssd1 vssd1 vccd1 vccd1 _15362_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_62_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12574_ _15335_/Q _13093_/A2 _12573_/X vssd1 vssd1 vccd1 vccd1 _15335_/D sky130_fd_sc_hd__a21o_1
XFILLER_62_96 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14313_ _15544_/CLK _14313_/D vssd1 vssd1 vccd1 vccd1 _14313_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_184_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11525_ _11544_/A _11526_/B vssd1 vssd1 vccd1 vccd1 _11531_/B sky130_fd_sc_hd__nand2b_1
XFILLER_8_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15293_ _15293_/CLK _15293_/D vssd1 vssd1 vccd1 vccd1 _15293_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14244_ _15289_/CLK _14244_/D vssd1 vssd1 vccd1 vccd1 _14244_/Q sky130_fd_sc_hd__dfxtp_1
X_11456_ _11457_/A _11457_/B vssd1 vssd1 vccd1 vccd1 _11472_/A sky130_fd_sc_hd__nor2_1
XFILLER_156_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_171_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10407_ _13171_/B _11414_/D vssd1 vssd1 vccd1 vccd1 _10410_/B sky130_fd_sc_hd__nand2_1
XFILLER_152_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14175_ _15661_/CLK _14175_/D vssd1 vssd1 vccd1 vccd1 _14175_/Q sky130_fd_sc_hd__dfxtp_1
X_11387_ _11386_/X _15047_/Q _11641_/S vssd1 vssd1 vccd1 vccd1 _15047_/D sky130_fd_sc_hd__mux2_1
XFILLER_113_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13126_ _14609_/Q _13125_/X _08536_/A _14608_/Q vssd1 vssd1 vccd1 vccd1 _13126_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10338_ _14723_/Q _14916_/Q _10343_/S vssd1 vssd1 vccd1 vccd1 _14723_/D sky130_fd_sc_hd__mux2_1
XTAP_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13057_ _15496_/Q _10877_/S _13042_/A _13056_/X vssd1 vssd1 vccd1 vccd1 _15496_/D
+ sky130_fd_sc_hd__a22o_1
X_10269_ _14654_/Q _14807_/Q _10630_/S vssd1 vssd1 vccd1 vccd1 _14654_/D sky130_fd_sc_hd__mux2_1
X_12008_ _06670_/A _12005_/X _06671_/A vssd1 vssd1 vccd1 vccd1 _12008_/X sky130_fd_sc_hd__o21a_1
XFILLER_94_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13959_ _15293_/CLK _13959_/D vssd1 vssd1 vccd1 vccd1 _13959_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_432 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07480_ _14760_/Q _07479_/X _07480_/S vssd1 vssd1 vccd1 vccd1 _07480_/X sky130_fd_sc_hd__mux2_8
XFILLER_50_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15629_ _15632_/CLK _15629_/D vssd1 vssd1 vccd1 vccd1 _15629_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_188_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09150_ _13951_/Q _13693_/Q _09407_/S vssd1 vssd1 vccd1 vccd1 _09150_/X sky130_fd_sc_hd__mux2_1
XFILLER_188_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08101_ input10/X input19/X _08145_/S vssd1 vssd1 vccd1 vccd1 _08159_/B sky130_fd_sc_hd__mux2_1
XFILLER_174_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09081_ _15282_/Q _15250_/Q _15218_/Q _15149_/Q _09190_/S _09429_/S1 vssd1 vssd1
+ vccd1 vccd1 _09081_/X sky130_fd_sc_hd__mux4_1
XFILLER_174_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08032_ _14737_/Q _08027_/X _08031_/X _12832_/C1 vssd1 vssd1 vccd1 vccd1 _13574_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_174_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09983_ _11870_/A1 _14342_/Q _09996_/S vssd1 vssd1 vccd1 vccd1 _14342_/D sky130_fd_sc_hd__mux2_1
XFILLER_66_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08934_ _14424_/Q _08540_/B _08520_/B _08933_/X vssd1 vssd1 vccd1 vccd1 _08934_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_57_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08865_ _13886_/Q _13074_/B2 _08880_/S vssd1 vssd1 vccd1 vccd1 _13886_/D sky130_fd_sc_hd__mux2_1
XTAP_3707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07816_ _07816_/A _07816_/B vssd1 vssd1 vccd1 vccd1 _07816_/Y sky130_fd_sc_hd__nand2_1
XTAP_3729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08796_ _13330_/A0 _13822_/Q _08811_/S vssd1 vssd1 vccd1 vccd1 _13822_/D sky130_fd_sc_hd__mux2_1
XFILLER_84_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07747_ _07745_/Y _07757_/D _07750_/A vssd1 vssd1 vccd1 vccd1 _07747_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_25_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07678_ _13481_/Q _07679_/C _13482_/Q vssd1 vssd1 vccd1 vccd1 _07678_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_26_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09417_ _14253_/Q _14285_/Q _14317_/Q _14349_/Q _09444_/S _09446_/A1 vssd1 vssd1
+ vccd1 vccd1 _09417_/X sky130_fd_sc_hd__mux4_1
XFILLER_40_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_159 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09348_ _14378_/Q _15194_/Q _13833_/Q _14572_/Q _09521_/S _09523_/A1 vssd1 vssd1
+ vccd1 vccd1 _09349_/B sky130_fd_sc_hd__mux4_1
XFILLER_21_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09279_ _15094_/Q _08540_/B _09278_/X _08501_/A vssd1 vssd1 vccd1 vccd1 _09279_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_138_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11310_ _15035_/Q _11302_/A _08321_/X _11303_/A _11309_/Y vssd1 vssd1 vccd1 vccd1
+ _15035_/D sky130_fd_sc_hd__o221a_1
X_12290_ _14020_/Q _13988_/Q _12543_/S vssd1 vssd1 vccd1 vccd1 _12291_/B sky130_fd_sc_hd__mux2_1
XFILLER_107_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11241_ _10420_/A _11239_/Y _11240_/Y _11240_/B _15026_/Q vssd1 vssd1 vccd1 vccd1
+ _15026_/D sky130_fd_sc_hd__a32o_1
XFILLER_4_347 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_1079 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11172_ _14978_/Q _11164_/S _11171_/X vssd1 vssd1 vccd1 vccd1 _14978_/D sky130_fd_sc_hd__o21a_1
XFILLER_122_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10123_ _14509_/Q _14757_/Q _10124_/S vssd1 vssd1 vccd1 vccd1 _14509_/D sky130_fd_sc_hd__mux2_1
XFILLER_79_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10054_ _14411_/Q _11873_/A1 _10064_/S vssd1 vssd1 vccd1 vccd1 _14411_/D sky130_fd_sc_hd__mux2_1
XFILLER_94_118 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14931_ _15556_/CLK _14931_/D vssd1 vssd1 vccd1 vccd1 _14931_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_76_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14862_ _15462_/CLK _14862_/D vssd1 vssd1 vccd1 vccd1 _14862_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13813_ _15142_/CLK _13813_/D vssd1 vssd1 vccd1 vccd1 _13813_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14793_ _15644_/CLK _14793_/D vssd1 vssd1 vccd1 vccd1 _14793_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13744_ _14649_/CLK _13744_/D vssd1 vssd1 vccd1 vccd1 _13744_/Q sky130_fd_sc_hd__dfxtp_1
X_10956_ _11013_/A _13233_/B vssd1 vssd1 vccd1 vccd1 _11317_/B sky130_fd_sc_hd__and2_1
XFILLER_17_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13675_ _15612_/CLK _13675_/D vssd1 vssd1 vccd1 vccd1 _13675_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10887_ _14919_/Q _15550_/Q _13134_/A vssd1 vssd1 vccd1 vccd1 _14919_/D sky130_fd_sc_hd__mux2_1
XFILLER_176_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15414_ _15596_/CLK _15414_/D vssd1 vssd1 vccd1 vccd1 _15414_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_176_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12626_ _13415_/Q _12640_/S _12625_/X vssd1 vssd1 vccd1 vccd1 _12627_/B sky130_fd_sc_hd__o21ai_1
XFILLER_188_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15345_ _15453_/CLK _15345_/D vssd1 vssd1 vccd1 vccd1 _15345_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_129_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12557_ _14385_/Q _15201_/Q _13840_/Q _14579_/Q _12568_/S _12567_/A vssd1 vssd1 vccd1
+ vccd1 _12557_/X sky130_fd_sc_hd__mux4_1
XFILLER_145_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11508_ _11546_/A _11508_/B vssd1 vssd1 vccd1 vccd1 _11508_/X sky130_fd_sc_hd__xor2_1
XFILLER_156_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15276_ _15276_/CLK _15276_/D vssd1 vssd1 vccd1 vccd1 _15276_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_1006 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12488_ _14382_/Q _15198_/Q _13837_/Q _14576_/Q _12489_/S0 _12489_/S1 vssd1 vssd1
+ vccd1 vccd1 _12488_/X sky130_fd_sc_hd__mux4_1
XFILLER_156_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14227_ _14485_/CLK _14227_/D vssd1 vssd1 vccd1 vccd1 _14227_/Q sky130_fd_sc_hd__dfxtp_1
X_11439_ _11476_/B _11439_/B vssd1 vssd1 vccd1 vccd1 _11440_/B sky130_fd_sc_hd__xnor2_4
XFILLER_125_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14158_ _15334_/CLK _14158_/D vssd1 vssd1 vccd1 vccd1 _14158_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13109_ _15522_/Q _10877_/S _13042_/A _13108_/X vssd1 vssd1 vccd1 vccd1 _15522_/D
+ sky130_fd_sc_hd__a22o_1
XTAP_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14089_ _15654_/CLK _14089_/D vssd1 vssd1 vccd1 vccd1 _14089_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06980_ _06879_/B _06877_/X _06882_/Y _06979_/X vssd1 vssd1 vccd1 vccd1 _13578_/D
+ sky130_fd_sc_hd__a22o_2
XFILLER_79_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08650_ _13491_/Q _08691_/B1 _08693_/B1 _13626_/Q vssd1 vssd1 vccd1 vccd1 _08650_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_187_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07601_ _14750_/Q _07607_/A _07600_/Y _07949_/C1 vssd1 vssd1 vccd1 vccd1 _13461_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_82_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08581_ _13469_/Q _08746_/A2 _08693_/B1 _13636_/Q vssd1 vssd1 vccd1 vccd1 _08581_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_19_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07532_ _14762_/Q _13441_/Q _07535_/S vssd1 vssd1 vccd1 vccd1 _13441_/D sky130_fd_sc_hd__mux2_1
XFILLER_35_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07463_ _13671_/Q _07499_/A2 _07499_/B1 _14699_/Q _07462_/X vssd1 vssd1 vccd1 vccd1
+ _07463_/X sky130_fd_sc_hd__a221o_1
XFILLER_139_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09202_ _09437_/A1 _09199_/X _09201_/X _09405_/A vssd1 vssd1 vccd1 vccd1 _09202_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_179_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07394_ _14650_/Q _07498_/B _07498_/C vssd1 vssd1 vccd1 vccd1 _07394_/X sky130_fd_sc_hd__and3_1
X_09133_ _09429_/S1 _09449_/A1 _09132_/X _09450_/B1 vssd1 vssd1 vccd1 vccd1 _09133_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_72_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09064_ _15657_/Q _13391_/Q _09230_/S vssd1 vssd1 vccd1 vccd1 _09064_/X sky130_fd_sc_hd__mux2_1
XFILLER_136_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08015_ _08018_/B _08014_/Y _08022_/B vssd1 vssd1 vccd1 vccd1 _08015_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_116_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_532 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09966_ _11853_/A1 _14325_/Q _09996_/S vssd1 vssd1 vccd1 vccd1 _14325_/D sky130_fd_sc_hd__mux2_1
XFILLER_131_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08917_ _14004_/Q _13972_/Q _09557_/S vssd1 vssd1 vccd1 vccd1 _08917_/X sky130_fd_sc_hd__mux2_1
XTAP_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09897_ _13350_/A0 _14259_/Q _09897_/S vssd1 vssd1 vccd1 vccd1 _14259_/D sky130_fd_sc_hd__mux2_1
XFILLER_134_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_96_clk clkbuf_5_24_0_clk/X vssd1 vssd1 vccd1 vccd1 _15645_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08848_ _13871_/Q _11847_/A1 _08851_/S vssd1 vssd1 vccd1 vccd1 _13871_/D sky130_fd_sc_hd__mux2_1
XFILLER_73_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08779_ _08779_/A _08779_/B _08779_/C vssd1 vssd1 vccd1 vccd1 _08779_/X sky130_fd_sc_hd__or3_1
XTAP_2825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10810_ _14842_/Q _07289_/X _12481_/A vssd1 vssd1 vccd1 vccd1 _14842_/D sky130_fd_sc_hd__mux2_1
XTAP_2847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11790_ _15213_/Q _13323_/A0 _11816_/S vssd1 vssd1 vccd1 vccd1 _15213_/D sky130_fd_sc_hd__mux2_1
XTAP_2869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10741_ _15405_/Q _14773_/Q _10765_/S vssd1 vssd1 vccd1 vccd1 _14773_/D sky130_fd_sc_hd__mux2_1
XFILLER_13_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13460_ _15383_/CLK _13460_/D vssd1 vssd1 vccd1 vccd1 _13460_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10672_ _15013_/Q _10717_/A2 _10652_/B _15030_/Q _10717_/C1 vssd1 vssd1 vccd1 vccd1
+ _10672_/X sky130_fd_sc_hd__a221o_1
XFILLER_159_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12411_ _12595_/A1 _12410_/X _12409_/X _12618_/C1 vssd1 vssd1 vccd1 vccd1 _12412_/C
+ sky130_fd_sc_hd__a211o_1
X_13391_ _15657_/CLK _13391_/D vssd1 vssd1 vccd1 vccd1 _13391_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_139_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_20_clk clkbuf_5_3_0_clk/X vssd1 vssd1 vccd1 vccd1 _15664_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_182_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15130_ _15130_/CLK _15130_/D vssd1 vssd1 vccd1 vccd1 _15130_/Q sky130_fd_sc_hd__dfxtp_1
X_12342_ _12618_/A1 _12341_/X _12340_/X _12618_/C1 vssd1 vssd1 vccd1 vccd1 _12343_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_126_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15061_ _15067_/CLK _15061_/D vssd1 vssd1 vccd1 vccd1 _15061_/Q sky130_fd_sc_hd__dfxtp_4
X_12273_ _12273_/A1 _12272_/X _12271_/X _12503_/C1 vssd1 vssd1 vccd1 vccd1 _12274_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_107_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14012_ _14415_/CLK _14012_/D vssd1 vssd1 vccd1 vccd1 _14012_/Q sky130_fd_sc_hd__dfxtp_1
X_11224_ _10528_/D _15012_/Q _11232_/S vssd1 vssd1 vccd1 vccd1 _15012_/D sky130_fd_sc_hd__mux2_1
XFILLER_107_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_175_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11155_ _11129_/A _11105_/B _11129_/Y vssd1 vssd1 vccd1 vccd1 _11197_/B sky130_fd_sc_hd__a21oi_2
XFILLER_110_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10106_ _14492_/Q _14740_/Q _10131_/S vssd1 vssd1 vccd1 vccd1 _14492_/D sky130_fd_sc_hd__mux2_1
XFILLER_95_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11086_ _11084_/X _11085_/X _11297_/S vssd1 vssd1 vccd1 vccd1 _11086_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_87_clk clkbuf_5_13_0_clk/X vssd1 vssd1 vccd1 vccd1 _15612_/CLK sky130_fd_sc_hd__clkbuf_16
X_10037_ _14394_/Q _11681_/A0 _10059_/S vssd1 vssd1 vccd1 vccd1 _14394_/D sky130_fd_sc_hd__mux2_1
X_14914_ _15670_/CLK _14914_/D vssd1 vssd1 vccd1 vccd1 _14914_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14845_ _15587_/CLK _14845_/D vssd1 vssd1 vccd1 vccd1 _14845_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14776_ _15626_/CLK _14776_/D vssd1 vssd1 vccd1 vccd1 _14776_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11988_ _11992_/A _11988_/B vssd1 vssd1 vccd1 vccd1 _11988_/X sky130_fd_sc_hd__and2_1
XFILLER_90_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13727_ _15020_/CLK _13727_/D vssd1 vssd1 vccd1 vccd1 _13727_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10939_ _14954_/Q _10455_/A _10944_/B vssd1 vssd1 vccd1 vccd1 _14954_/D sky130_fd_sc_hd__mux2_1
XFILLER_16_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_1027 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13658_ _14774_/CLK _13658_/D vssd1 vssd1 vccd1 vccd1 _13658_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12609_ _12613_/A _12609_/B vssd1 vssd1 vccd1 vccd1 _12609_/X sky130_fd_sc_hd__and2_1
XFILLER_158_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13589_ _15453_/CLK _13589_/D vssd1 vssd1 vccd1 vccd1 _13589_/Q sky130_fd_sc_hd__dfxtp_2
Xclkbuf_leaf_11_clk clkbuf_5_2_0_clk/X vssd1 vssd1 vccd1 vccd1 _15218_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_76_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15328_ _15328_/CLK _15328_/D vssd1 vssd1 vccd1 vccd1 _15328_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15259_ _15259_/CLK _15259_/D vssd1 vssd1 vccd1 vccd1 _15259_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_173_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout407 _11641_/S vssd1 vssd1 vccd1 vccd1 _11614_/S sky130_fd_sc_hd__clkbuf_16
X_09820_ _14186_/Q _13342_/A0 _09828_/S vssd1 vssd1 vccd1 vccd1 _14186_/D sky130_fd_sc_hd__mux2_1
Xfanout418 _10733_/B1 vssd1 vssd1 vccd1 vccd1 _10722_/B1 sky130_fd_sc_hd__buf_12
Xfanout429 _08497_/A vssd1 vssd1 vccd1 vccd1 _09419_/A2 sky130_fd_sc_hd__buf_12
XFILLER_140_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09751_ _14119_/Q _13092_/B2 _09762_/S vssd1 vssd1 vccd1 vccd1 _14119_/D sky130_fd_sc_hd__mux2_1
X_06963_ _06963_/A _06963_/B vssd1 vssd1 vccd1 vccd1 _06963_/Y sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_78_clk clkbuf_5_15_0_clk/X vssd1 vssd1 vccd1 vccd1 _15608_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_95_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08702_ _13420_/Q _08535_/X _08699_/X _08701_/X _10765_/S vssd1 vssd1 vccd1 vccd1
+ _08702_/X sky130_fd_sc_hd__a2111o_1
XFILLER_104_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09682_ _14053_/Q _13337_/A0 _09695_/S vssd1 vssd1 vccd1 vccd1 _14053_/D sky130_fd_sc_hd__mux2_1
X_06894_ _15383_/Q _07595_/A vssd1 vssd1 vccd1 vccd1 _06894_/X sky130_fd_sc_hd__and2_1
XFILLER_27_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08633_ _13789_/Q _08626_/S _08632_/X vssd1 vssd1 vccd1 vccd1 _13789_/D sky130_fd_sc_hd__o21a_1
XFILLER_54_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08564_ _15395_/Q _08748_/A2 _08736_/A2 _13440_/Q vssd1 vssd1 vccd1 vccd1 _08564_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_81_154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07515_ _14745_/Q _13424_/Q _07529_/S vssd1 vssd1 vccd1 vccd1 _13424_/D sky130_fd_sc_hd__mux2_1
XFILLER_81_187 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_744 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08495_ _08668_/B _08519_/B vssd1 vssd1 vccd1 vccd1 _13125_/A sky130_fd_sc_hd__nand2_8
X_07446_ _14663_/Q _07474_/B _07498_/C vssd1 vssd1 vccd1 vccd1 _07446_/X sky130_fd_sc_hd__and3_1
XFILLER_149_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07377_ _11852_/A1 _13383_/Q _07481_/S vssd1 vssd1 vccd1 vccd1 _13383_/D sky130_fd_sc_hd__mux2_1
XFILLER_129_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09116_ _13917_/Q _09115_/X _12504_/A vssd1 vssd1 vccd1 vccd1 _13917_/D sky130_fd_sc_hd__mux2_1
XFILLER_108_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_175_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09047_ _13946_/Q _13688_/Q _09047_/S vssd1 vssd1 vccd1 vccd1 _09047_/X sky130_fd_sc_hd__mux2_1
XFILLER_124_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09949_ _11761_/A0 _14309_/Q _09963_/S vssd1 vssd1 vccd1 vccd1 _14309_/D sky130_fd_sc_hd__mux2_1
XFILLER_49_129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_69_clk clkbuf_5_14_0_clk/X vssd1 vssd1 vccd1 vccd1 _15067_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_93_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12960_ _10604_/X _14867_/Q _13038_/S vssd1 vssd1 vccd1 vccd1 _12960_/X sky130_fd_sc_hd__mux2_2
XTAP_4046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11911_ _15109_/Q _15077_/Q _15650_/Q _13384_/Q _12614_/S _12383_/A vssd1 vssd1 vccd1
+ vccd1 _11911_/X sky130_fd_sc_hd__mux4_1
XTAP_4079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12891_ _15419_/Q _15604_/Q _12932_/S vssd1 vssd1 vccd1 vccd1 _15419_/D sky130_fd_sc_hd__mux2_1
XFILLER_72_110 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14630_ _15634_/CLK _14630_/D vssd1 vssd1 vccd1 vccd1 _14630_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_166_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11842_ _15264_/Q _13342_/A0 _11850_/S vssd1 vssd1 vccd1 vccd1 _15264_/D sky130_fd_sc_hd__mux2_1
XTAP_2644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_64 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14561_ _15220_/CLK _14561_/D vssd1 vssd1 vccd1 vccd1 _14561_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11773_ _13348_/A0 _15201_/Q _11775_/S vssd1 vssd1 vccd1 vccd1 _15201_/D sky130_fd_sc_hd__mux2_1
XTAP_1954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13512_ _15372_/CLK _13512_/D vssd1 vssd1 vccd1 vccd1 _13512_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10724_ _15072_/Q _10734_/A2 _10721_/X _10723_/X vssd1 vssd1 vccd1 vccd1 _10724_/X
+ sky130_fd_sc_hd__o22a_4
XFILLER_159_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14492_ _15374_/CLK _14492_/D vssd1 vssd1 vccd1 vccd1 _14492_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_5_3_0_clk clkbuf_5_3_0_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_5_3_0_clk/X sky130_fd_sc_hd__clkbuf_8
X_13443_ _15461_/CLK _13443_/D vssd1 vssd1 vccd1 vccd1 _13443_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_174_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10655_ _14749_/Q _10654_/X _10710_/S vssd1 vssd1 vccd1 vccd1 _14749_/D sky130_fd_sc_hd__mux2_1
XFILLER_142_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13374_ _14477_/Q vssd1 vssd1 vccd1 vccd1 _14477_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_103_1044 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10586_ _14996_/Q _10569_/B _10733_/A2 _14964_/Q _10732_/C1 vssd1 vssd1 vccd1 vccd1
+ _10586_/X sky130_fd_sc_hd__a221o_1
XFILLER_62_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15113_ _15211_/CLK _15113_/D vssd1 vssd1 vccd1 vccd1 _15113_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_420 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12325_ _15127_/Q _15095_/Q _15668_/Q _13402_/Q _12543_/S _12544_/A vssd1 vssd1 vccd1
+ vccd1 _12325_/X sky130_fd_sc_hd__mux4_1
XFILLER_103_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15044_ _15306_/CLK _15044_/D vssd1 vssd1 vccd1 vccd1 _15044_/Q sky130_fd_sc_hd__dfxtp_1
X_12256_ _15124_/Q _15092_/Q _15665_/Q _13399_/Q _12269_/S _12268_/A vssd1 vssd1 vccd1
+ vccd1 _12256_/X sky130_fd_sc_hd__mux4_1
XFILLER_107_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11207_ _10556_/C _14996_/Q _11237_/S vssd1 vssd1 vccd1 vccd1 _14996_/D sky130_fd_sc_hd__mux2_1
X_12187_ _15121_/Q _15089_/Q _15662_/Q _13396_/Q _12489_/S0 _12465_/S1 vssd1 vssd1
+ vccd1 vccd1 _12187_/X sky130_fd_sc_hd__mux4_1
XFILLER_95_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11138_ _11344_/A _11189_/B _11137_/X vssd1 vssd1 vccd1 vccd1 _11138_/Y sky130_fd_sc_hd__a21oi_1
X_11069_ _11356_/B _10999_/Y _11068_/X vssd1 vssd1 vccd1 vccd1 _11069_/X sky130_fd_sc_hd__a21o_1
Xclkbuf_leaf_0_clk clkbuf_5_0_0_clk/X vssd1 vssd1 vccd1 vccd1 _15277_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_37_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14828_ _15622_/CLK _14828_/D vssd1 vssd1 vccd1 vccd1 _14828_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14759_ _15607_/CLK _14759_/D vssd1 vssd1 vccd1 vccd1 _14759_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_177_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07300_ _13916_/Q _15503_/Q _07339_/S vssd1 vssd1 vccd1 vccd1 _07301_/A sky130_fd_sc_hd__mux2_8
X_08280_ _11356_/C _13165_/B _10999_/A vssd1 vssd1 vccd1 vccd1 _08280_/Y sky130_fd_sc_hd__o21bai_2
XFILLER_177_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07231_ _07356_/A _07231_/B _07231_/C _07230_/X vssd1 vssd1 vccd1 vccd1 _07355_/A
+ sky130_fd_sc_hd__or4b_1
XFILLER_146_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07162_ _14861_/Q _14853_/Q _14845_/Q _14837_/Q _07146_/S _08151_/S vssd1 vssd1 vccd1
+ vccd1 _07163_/B sky130_fd_sc_hd__mux4_1
XFILLER_146_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07093_ _14643_/Q _14675_/Q _07096_/S vssd1 vssd1 vccd1 vccd1 _07093_/X sky130_fd_sc_hd__mux2_2
XFILLER_173_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout204 _09730_/Y vssd1 vssd1 vccd1 vccd1 _09762_/S sky130_fd_sc_hd__buf_12
Xfanout215 _08853_/Y vssd1 vssd1 vccd1 vccd1 _08880_/S sky130_fd_sc_hd__buf_12
XFILLER_119_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout226 _07907_/Y vssd1 vssd1 vccd1 vccd1 _07964_/A sky130_fd_sc_hd__buf_8
XFILLER_99_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09803_ _14169_/Q _13325_/A0 _09823_/S vssd1 vssd1 vccd1 vccd1 _14169_/D sky130_fd_sc_hd__mux2_1
Xfanout237 _07004_/X vssd1 vssd1 vccd1 vccd1 _07098_/S sky130_fd_sc_hd__buf_12
Xfanout248 _08530_/Y vssd1 vssd1 vccd1 vccd1 _08685_/A2 sky130_fd_sc_hd__clkbuf_16
XFILLER_86_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07995_ _13565_/Q _13564_/Q _13563_/Q _07995_/D vssd1 vssd1 vccd1 vccd1 _08006_/D
+ sky130_fd_sc_hd__and4_2
XFILLER_59_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout259 _07370_/X vssd1 vssd1 vccd1 vccd1 _07481_/S sky130_fd_sc_hd__buf_12
X_09734_ _14102_/Q _11680_/A0 _09757_/S vssd1 vssd1 vccd1 vccd1 _14102_/D sky130_fd_sc_hd__mux2_1
X_06946_ _06738_/Y _13484_/Q _06740_/Y _13483_/Q vssd1 vssd1 vccd1 vccd1 _06946_/X
+ sky130_fd_sc_hd__a22o_2
XFILLER_95_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09665_ _14036_/Q _11853_/A1 _09695_/S vssd1 vssd1 vccd1 vccd1 _14036_/D sky130_fd_sc_hd__mux2_1
XFILLER_83_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06877_ _06882_/C _06877_/B vssd1 vssd1 vccd1 vccd1 _06877_/X sky130_fd_sc_hd__or2_1
XFILLER_28_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08616_ _13560_/Q _08685_/A2 _08691_/B1 _13496_/Q vssd1 vssd1 vccd1 vccd1 _08616_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_43_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09596_ _11710_/A _09696_/B vssd1 vssd1 vccd1 vccd1 _09596_/Y sky130_fd_sc_hd__nor2_8
XFILLER_82_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08547_ _13474_/Q _08746_/A2 _08747_/B1 _13506_/Q vssd1 vssd1 vccd1 vccd1 _08547_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_11_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08478_ _14607_/Q _08487_/B _08477_/X _08449_/A vssd1 vssd1 vccd1 vccd1 _08478_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_11_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07429_ _13332_/A0 _13396_/Q _07481_/S vssd1 vssd1 vccd1 vccd1 _13396_/D sky130_fd_sc_hd__mux2_1
XFILLER_183_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10440_ _11624_/A _11626_/A vssd1 vssd1 vccd1 vccd1 _10537_/B sky130_fd_sc_hd__nor2_1
XFILLER_136_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10371_ _07301_/A _10360_/B _10370_/X vssd1 vssd1 vccd1 vccd1 _11436_/B sky130_fd_sc_hd__a21oi_4
XFILLER_152_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12110_ _12103_/X _12105_/X _12107_/X _12109_/X _12501_/C1 vssd1 vssd1 vccd1 vccd1
+ _12110_/X sky130_fd_sc_hd__o221a_1
XFILLER_136_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13090_ _13002_/X _13118_/A2 _13114_/B1 _07452_/X vssd1 vssd1 vccd1 vccd1 _13090_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_6_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12041_ _12034_/X _12036_/X _12038_/X _12040_/X _06671_/A vssd1 vssd1 vccd1 vccd1
+ _12041_/X sky130_fd_sc_hd__o221a_1
XFILLER_46_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13992_ _15334_/CLK _13992_/D vssd1 vssd1 vccd1 vccd1 _13992_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_77_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12943_ _12943_/A _12943_/B _12943_/C vssd1 vssd1 vccd1 vccd1 _13116_/B sky130_fd_sc_hd__or3_2
XTAP_3131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_120 _07161_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15662_ _15662_/CLK _15662_/D vssd1 vssd1 vccd1 vccd1 _15662_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12874_ _15402_/Q _15587_/Q _12900_/S vssd1 vssd1 vccd1 vccd1 _15402_/D sky130_fd_sc_hd__mux2_1
XTAP_3186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_131 _14745_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11825_ _15247_/Q _11858_/A1 _11850_/S vssd1 vssd1 vccd1 vccd1 _15247_/D sky130_fd_sc_hd__mux2_1
X_14613_ _15648_/CLK _14613_/D vssd1 vssd1 vccd1 vccd1 _14613_/Q sky130_fd_sc_hd__dfxtp_4
X_15593_ _15626_/CLK _15593_/D vssd1 vssd1 vccd1 vccd1 _15593_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14544_ _15331_/CLK _14544_/D vssd1 vssd1 vccd1 vccd1 _14544_/Q sky130_fd_sc_hd__dfxtp_1
X_11756_ _13331_/A0 _15184_/Q _11774_/S vssd1 vssd1 vccd1 vccd1 _15184_/D sky130_fd_sc_hd__mux2_1
XTAP_1784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1027 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10707_ _15020_/Q _10717_/A2 _10652_/B _15037_/Q _10717_/C1 vssd1 vssd1 vccd1 vccd1
+ _10707_/X sky130_fd_sc_hd__a221o_1
XFILLER_186_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14475_ _14485_/CLK _14475_/D vssd1 vssd1 vccd1 vccd1 _14475_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_186_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11687_ _13329_/A0 _15118_/Q _11703_/S vssd1 vssd1 vccd1 vccd1 _15118_/D sky130_fd_sc_hd__mux2_1
XFILLER_128_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13426_ _15381_/CLK _13426_/D vssd1 vssd1 vccd1 vccd1 _13426_/Q sky130_fd_sc_hd__dfxtp_1
X_10638_ _14974_/Q _10718_/A2 _10722_/B1 _14942_/Q _10637_/X vssd1 vssd1 vccd1 vccd1
+ _10638_/X sky130_fd_sc_hd__a221o_2
XFILLER_139_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13357_ _14460_/Q vssd1 vssd1 vccd1 vccd1 _14460_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_6_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10569_ _10581_/A _10569_/B vssd1 vssd1 vccd1 vccd1 _10569_/Y sky130_fd_sc_hd__nand2_2
XFILLER_155_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12308_ _12595_/A1 _12303_/X _12306_/X _12307_/X _08405_/D vssd1 vssd1 vccd1 vccd1
+ _12320_/B sky130_fd_sc_hd__a221o_2
X_13288_ _12637_/Y _15620_/Q _13288_/S vssd1 vssd1 vccd1 vccd1 _15620_/D sky130_fd_sc_hd__mux2_1
XFILLER_64_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15027_ _15582_/CLK _15027_/D vssd1 vssd1 vccd1 vccd1 _15027_/Q sky130_fd_sc_hd__dfxtp_1
X_12239_ _12503_/A1 _12234_/X _12237_/X _12238_/X _08449_/A vssd1 vssd1 vccd1 vccd1
+ _12251_/B sky130_fd_sc_hd__a221o_1
XFILLER_114_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_799 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_1104 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06800_ _06799_/A _06797_/A _08773_/A _15615_/Q vssd1 vssd1 vccd1 vccd1 _06806_/A
+ sky130_fd_sc_hd__o211a_2
X_07780_ _07787_/A _08817_/B _13509_/Q vssd1 vssd1 vccd1 vccd1 _07780_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_110_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput4 ext_read_data[12] vssd1 vssd1 vccd1 vccd1 input4/X sky130_fd_sc_hd__clkbuf_8
X_06731_ _13456_/Q vssd1 vssd1 vccd1 vccd1 _06731_/Y sky130_fd_sc_hd__inv_2
XFILLER_65_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09450_ _09405_/A _09443_/X _09446_/X _09450_/B1 vssd1 vssd1 vccd1 vccd1 _09450_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_92_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06662_ _14899_/Q vssd1 vssd1 vccd1 vccd1 _06771_/C sky130_fd_sc_hd__inv_2
XFILLER_188_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08401_ _13734_/Q _10871_/S _08400_/X vssd1 vssd1 vccd1 vccd1 _13734_/D sky130_fd_sc_hd__o21a_1
XFILLER_51_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09381_ _08494_/B _09379_/X _09380_/X vssd1 vssd1 vccd1 vccd1 _09382_/C sky130_fd_sc_hd__a21o_1
XFILLER_51_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_1099 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08332_ _13722_/Q _08232_/A _11351_/C1 _08331_/X vssd1 vssd1 vccd1 vccd1 _13722_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_178_833 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08263_ _10507_/A1 _13772_/Q _15400_/Q _10515_/B2 vssd1 vssd1 vccd1 vccd1 _08263_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_177_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07214_ _15333_/Q _15489_/Q _07335_/S vssd1 vssd1 vccd1 vccd1 _07215_/A sky130_fd_sc_hd__mux2_8
X_08194_ _13685_/Q _11681_/A0 _08216_/S vssd1 vssd1 vccd1 vccd1 _13685_/D sky130_fd_sc_hd__mux2_1
XFILLER_118_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07145_ _14836_/Q _07104_/X _07144_/X _07131_/A vssd1 vssd1 vccd1 vccd1 _07145_/X
+ sky130_fd_sc_hd__a22o_4
XFILLER_145_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07076_ _07075_/X _13604_/Q _12764_/S vssd1 vssd1 vccd1 vccd1 _07076_/X sky130_fd_sc_hd__mux2_1
XFILLER_133_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_1048 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07978_ _13560_/Q _07984_/D vssd1 vssd1 vccd1 vccd1 _07978_/X sky130_fd_sc_hd__or2_1
XFILLER_28_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09717_ _13092_/B2 _14087_/Q _09728_/S vssd1 vssd1 vccd1 vccd1 _14087_/D sky130_fd_sc_hd__mux2_1
X_06929_ _06929_/A _06929_/B _06927_/X vssd1 vssd1 vccd1 vccd1 _06929_/X sky130_fd_sc_hd__or3b_1
X_09648_ _14021_/Q _13337_/A0 _09661_/S vssd1 vssd1 vccd1 vccd1 _14021_/D sky130_fd_sc_hd__mux2_1
XTAP_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09579_ _13955_/Q _13335_/A0 _09589_/S vssd1 vssd1 vccd1 vccd1 _13955_/D sky130_fd_sc_hd__mux2_1
XTAP_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11610_ _11610_/A _11610_/B vssd1 vssd1 vccd1 vccd1 _11612_/B sky130_fd_sc_hd__xnor2_2
XTAP_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12590_ _12590_/A _12590_/B vssd1 vssd1 vccd1 vccd1 _12590_/X sky130_fd_sc_hd__and2_1
XFILLER_143_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11541_ _13217_/B _11541_/B vssd1 vssd1 vccd1 vccd1 _11542_/B sky130_fd_sc_hd__nand2_1
XFILLER_23_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14260_ _15289_/CLK _14260_/D vssd1 vssd1 vccd1 vccd1 _14260_/Q sky130_fd_sc_hd__dfxtp_1
X_11472_ _11472_/A _11472_/B vssd1 vssd1 vccd1 vccd1 _11473_/B sky130_fd_sc_hd__nor2_1
XFILLER_51_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13211_ _13233_/A _11521_/A _11536_/C vssd1 vssd1 vccd1 vccd1 _13211_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_52_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10423_ _11349_/C vssd1 vssd1 vccd1 vccd1 _11633_/A sky130_fd_sc_hd__clkinv_4
X_14191_ _15094_/CLK _14191_/D vssd1 vssd1 vccd1 vccd1 _14191_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_733 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13142_ _08777_/A _08777_/B _08767_/Y _13129_/A _15539_/Q vssd1 vssd1 vccd1 vccd1
+ _15539_/D sky130_fd_sc_hd__a32o_1
X_10354_ _13199_/B _11496_/A vssd1 vssd1 vccd1 vccd1 _10356_/A sky130_fd_sc_hd__nand2_1
XFILLER_83_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13073_ _15504_/Q _13105_/A2 _13105_/B1 _13072_/X vssd1 vssd1 vccd1 vccd1 _15504_/D
+ sky130_fd_sc_hd__a22o_1
X_10285_ _14670_/Q _14823_/Q _10285_/S vssd1 vssd1 vccd1 vccd1 _14670_/D sky130_fd_sc_hd__mux2_1
XFILLER_2_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12024_ _14460_/Q _14428_/Q _13849_/Q _14202_/Q _12079_/S _12080_/A vssd1 vssd1 vccd1
+ vccd1 _12024_/X sky130_fd_sc_hd__mux4_1
XFILLER_78_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_51 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout590 _12486_/S1 vssd1 vssd1 vccd1 vccd1 _12489_/S1 sky130_fd_sc_hd__buf_12
XFILLER_47_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13975_ _15253_/CLK _13975_/D vssd1 vssd1 vccd1 vccd1 _13975_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_964 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12926_ _15454_/Q _15640_/Q _12927_/S vssd1 vssd1 vccd1 vccd1 _15454_/D sky130_fd_sc_hd__mux2_1
XFILLER_62_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15645_ _15645_/CLK _15645_/D vssd1 vssd1 vccd1 vccd1 _15645_/Q sky130_fd_sc_hd__dfxtp_1
X_12857_ _14751_/Q _15385_/Q _12866_/S vssd1 vssd1 vccd1 vccd1 _15385_/D sky130_fd_sc_hd__mux2_1
XTAP_2271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11808_ _15231_/Q _11874_/A1 _11817_/S vssd1 vssd1 vccd1 vccd1 _15231_/D sky130_fd_sc_hd__mux2_1
X_12788_ _15360_/Q _12765_/B _12784_/X _12787_/X _12788_/C1 vssd1 vssd1 vccd1 vccd1
+ _15360_/D sky130_fd_sc_hd__o221a_1
XTAP_1570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15576_ _15613_/CLK _15576_/D vssd1 vssd1 vccd1 vccd1 _15576_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_42_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14527_ _15658_/CLK _14527_/D vssd1 vssd1 vccd1 vccd1 _14527_/Q sky130_fd_sc_hd__dfxtp_1
X_11739_ _15168_/Q _11847_/A1 _11742_/S vssd1 vssd1 vccd1 vccd1 _15168_/D sky130_fd_sc_hd__mux2_1
XFILLER_186_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14458_ _15273_/CLK _14458_/D vssd1 vssd1 vccd1 vccd1 _14458_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13409_ _15675_/CLK _13409_/D vssd1 vssd1 vccd1 vccd1 _13409_/Q sky130_fd_sc_hd__dfxtp_1
X_14389_ _15617_/CLK _14389_/D vssd1 vssd1 vccd1 vccd1 _14389_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08950_ _13909_/Q _10877_/S _08949_/X vssd1 vssd1 vccd1 vccd1 _13909_/D sky130_fd_sc_hd__a21o_1
XFILLER_9_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07901_ _13539_/Q _07900_/C _07900_/D _13540_/Q vssd1 vssd1 vccd1 vccd1 _07902_/B
+ sky130_fd_sc_hd__a31o_1
X_08881_ _13902_/Q _13346_/A0 _08885_/S vssd1 vssd1 vccd1 vccd1 _13902_/D sky130_fd_sc_hd__mux2_1
XFILLER_155_1092 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07832_ _13522_/Q _13521_/Q _07836_/D vssd1 vssd1 vccd1 vccd1 _07837_/B sky130_fd_sc_hd__and3_1
XFILLER_84_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07763_ _14761_/Q _07777_/A _07762_/Y _08012_/C1 vssd1 vssd1 vccd1 vccd1 _13504_/D
+ sky130_fd_sc_hd__o211a_1
X_09502_ _14483_/Q _09558_/A2 _13130_/B1 _14451_/Q _09501_/X vssd1 vssd1 vccd1 vccd1
+ _09502_/X sky130_fd_sc_hd__a221o_1
X_06714_ _15387_/Q vssd1 vssd1 vccd1 vccd1 _06714_/Y sky130_fd_sc_hd__inv_2
XFILLER_112_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07694_ _13486_/Q _13485_/Q _07717_/A vssd1 vssd1 vccd1 vccd1 _07697_/B sky130_fd_sc_hd__and3_2
XFILLER_25_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09433_ _13932_/Q _13081_/A2 _09432_/X vssd1 vssd1 vccd1 vccd1 _13932_/D sky130_fd_sc_hd__a21o_1
XFILLER_52_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09364_ _14540_/Q _14153_/Q _14185_/Q _14121_/Q _09521_/S _09523_/A1 vssd1 vssd1
+ vccd1 vccd1 _09364_/X sky130_fd_sc_hd__mux4_1
XFILLER_52_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_1044 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08315_ _11356_/C _13178_/B vssd1 vssd1 vccd1 vccd1 _08316_/B sky130_fd_sc_hd__nor2_1
X_09295_ _13958_/Q _13700_/Q _09484_/S vssd1 vssd1 vccd1 vccd1 _09295_/X sky130_fd_sc_hd__mux2_1
XANTENNA_20 _14606_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_31 _14749_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_42 input19/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_53 _07191_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08246_ _07332_/X _10481_/B _08245_/X vssd1 vssd1 vccd1 vccd1 _10895_/B sky130_fd_sc_hd__a21o_4
XFILLER_123_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_64 _06865_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_75 _07153_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_86 _07903_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_97 _11563_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08177_ _08133_/S input20/X _08185_/A vssd1 vssd1 vccd1 vccd1 _08177_/X sky130_fd_sc_hd__and3b_1
XFILLER_21_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_891 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07128_ _14844_/Q _14836_/Q _08094_/S vssd1 vssd1 vccd1 vccd1 _07129_/B sky130_fd_sc_hd__mux2_1
XFILLER_137_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07059_ _07058_/X _14752_/Q _07077_/S vssd1 vssd1 vccd1 vccd1 _13598_/D sky130_fd_sc_hd__mux2_1
XFILLER_115_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10070_ _14426_/Q _13323_/A0 _10092_/S vssd1 vssd1 vccd1 vccd1 _14426_/D sky130_fd_sc_hd__mux2_1
XFILLER_121_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_663 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_463 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13760_ _14888_/CLK _13760_/D vssd1 vssd1 vccd1 vccd1 _13760_/Q sky130_fd_sc_hd__dfxtp_1
X_10972_ _11259_/S _10972_/B vssd1 vssd1 vccd1 vccd1 _10972_/X sky130_fd_sc_hd__or2_1
XFILLER_44_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12711_ _12723_/C _12711_/B vssd1 vssd1 vccd1 vccd1 _12711_/X sky130_fd_sc_hd__and2b_1
XFILLER_188_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13691_ _14093_/CLK _13691_/D vssd1 vssd1 vccd1 vccd1 _13691_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_71 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15430_ _15434_/CLK _15430_/D vssd1 vssd1 vccd1 vccd1 _15430_/Q sky130_fd_sc_hd__dfxtp_1
X_12642_ _15340_/Q _12759_/B _12641_/X _12832_/C1 vssd1 vssd1 vccd1 vccd1 _15340_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_188_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15361_ _15641_/CLK _15361_/D vssd1 vssd1 vccd1 vccd1 _15361_/Q sky130_fd_sc_hd__dfxtp_2
X_12573_ _12573_/A _12573_/B _12573_/C vssd1 vssd1 vccd1 vccd1 _12573_/X sky130_fd_sc_hd__and3_1
XFILLER_129_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11524_ _11546_/A _11508_/B _11546_/B _11523_/Y vssd1 vssd1 vccd1 vccd1 _11526_/B
+ sky130_fd_sc_hd__a31o_1
X_14312_ _15669_/CLK _14312_/D vssd1 vssd1 vccd1 vccd1 _14312_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15292_ _15292_/CLK _15292_/D vssd1 vssd1 vccd1 vccd1 _15292_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_178_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14243_ _15306_/CLK _14243_/D vssd1 vssd1 vccd1 vccd1 _14243_/Q sky130_fd_sc_hd__dfxtp_1
X_11455_ _11475_/B _11455_/B vssd1 vssd1 vccd1 vccd1 _11457_/B sky130_fd_sc_hd__xnor2_1
XFILLER_184_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10406_ _11371_/A _13165_/B _11383_/A _11380_/A _10405_/X vssd1 vssd1 vccd1 vccd1
+ _10406_/X sky130_fd_sc_hd__a221o_1
X_14174_ _15253_/CLK _14174_/D vssd1 vssd1 vccd1 vccd1 _14174_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_178_1070 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11386_ _11401_/A _11386_/B vssd1 vssd1 vccd1 vccd1 _11386_/X sky130_fd_sc_hd__xor2_1
XFILLER_152_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13125_ _13125_/A _13125_/B _14610_/Q vssd1 vssd1 vccd1 vccd1 _13125_/X sky130_fd_sc_hd__or3b_1
XFILLER_113_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10337_ _14722_/Q _14915_/Q _10343_/S vssd1 vssd1 vccd1 vccd1 _14722_/D sky130_fd_sc_hd__mux2_1
XTAP_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13056_ _12951_/X _13118_/A2 _13114_/B1 _07384_/X vssd1 vssd1 vccd1 vccd1 _13056_/X
+ sky130_fd_sc_hd__a22o_1
X_10268_ _14653_/Q hold7/X _10285_/S vssd1 vssd1 vccd1 vccd1 _14653_/D sky130_fd_sc_hd__mux2_1
XFILLER_105_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12007_ _12594_/S _12007_/B vssd1 vssd1 vccd1 vccd1 _12007_/X sky130_fd_sc_hd__or2_1
XFILLER_39_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10199_ input12/X _14584_/Q _13284_/S vssd1 vssd1 vccd1 vccd1 _14584_/D sky130_fd_sc_hd__mux2_1
XFILLER_38_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_1060 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13958_ _15127_/CLK _13958_/D vssd1 vssd1 vccd1 vccd1 _13958_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12909_ _15437_/Q _15623_/Q _12933_/S vssd1 vssd1 vccd1 vccd1 _15437_/D sky130_fd_sc_hd__mux2_1
XFILLER_34_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13889_ _14415_/CLK _13889_/D vssd1 vssd1 vccd1 vccd1 _13889_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15628_ _15628_/CLK _15628_/D vssd1 vssd1 vccd1 vccd1 _15628_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_107_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15559_ _15613_/CLK _15559_/D vssd1 vssd1 vccd1 vccd1 _15559_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_147_313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08100_ _13650_/Q _10344_/S _08096_/X _08099_/X vssd1 vssd1 vccd1 vccd1 _13650_/D
+ sky130_fd_sc_hd__a22o_1
X_09080_ _09221_/A _09080_/B vssd1 vssd1 vccd1 vccd1 _09080_/X sky130_fd_sc_hd__or2_1
XFILLER_148_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08031_ _13574_/Q _06861_/Y _08030_/Y _13573_/Q _08028_/B vssd1 vssd1 vccd1 vccd1
+ _08031_/X sky130_fd_sc_hd__a221o_1
XFILLER_174_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09982_ _13086_/B2 _14341_/Q _09996_/S vssd1 vssd1 vccd1 vccd1 _14341_/D sky130_fd_sc_hd__mux2_1
XFILLER_107_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08933_ _13845_/Q _14198_/Q _09484_/S vssd1 vssd1 vccd1 vccd1 _08933_/X sky130_fd_sc_hd__mux2_1
XFILLER_88_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08864_ _13885_/Q _13072_/B2 _08880_/S vssd1 vssd1 vccd1 vccd1 _13885_/D sky130_fd_sc_hd__mux2_1
XFILLER_130_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07815_ _07825_/D _07815_/B vssd1 vssd1 vccd1 vccd1 _07816_/B sky130_fd_sc_hd__nand2b_1
XFILLER_57_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08795_ _13329_/A0 _13821_/Q _08811_/S vssd1 vssd1 vccd1 vccd1 _13821_/D sky130_fd_sc_hd__mux2_1
XFILLER_72_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_912 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07746_ _13500_/Q _13499_/Q _07746_/C vssd1 vssd1 vccd1 vccd1 _07757_/D sky130_fd_sc_hd__and3_2
XFILLER_38_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07677_ _14738_/Q _07676_/A _07676_/Y _08084_/C1 vssd1 vssd1 vccd1 vccd1 _13481_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_26_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09416_ _09437_/A1 _09415_/X _09414_/X _09405_/A vssd1 vssd1 vccd1 vccd1 _09416_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_25_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_274 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09347_ _13928_/Q _13154_/S _09346_/X vssd1 vssd1 vccd1 vccd1 _13928_/D sky130_fd_sc_hd__a21o_1
XFILLER_166_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09278_ _15126_/Q _09558_/A2 _13130_/C1 _09277_/X vssd1 vssd1 vccd1 vccd1 _09278_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_181_603 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08229_ _08240_/A _13802_/Q _13770_/Q _08237_/A vssd1 vssd1 vccd1 vccd1 _08229_/X
+ sky130_fd_sc_hd__a22o_2
XFILLER_126_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11240_ _11240_/A _11240_/B vssd1 vssd1 vccd1 vccd1 _11240_/Y sky130_fd_sc_hd__nor2_1
XFILLER_162_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_255_clk clkbuf_5_0_0_clk/X vssd1 vssd1 vccd1 vccd1 _15209_/CLK sky130_fd_sc_hd__clkbuf_16
X_11171_ _08233_/B _10982_/X _11170_/X vssd1 vssd1 vccd1 vccd1 _11171_/X sky130_fd_sc_hd__a21o_1
XFILLER_121_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10122_ _14508_/Q _14756_/Q _10124_/S vssd1 vssd1 vccd1 vccd1 _14508_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_543 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10053_ _14410_/Q _11872_/A1 _10064_/S vssd1 vssd1 vccd1 vccd1 _14410_/D sky130_fd_sc_hd__mux2_1
X_14930_ _15046_/CLK _14930_/D vssd1 vssd1 vccd1 vccd1 _14930_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14861_ _14861_/CLK _14861_/D vssd1 vssd1 vccd1 vccd1 _14861_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_180_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13812_ _14197_/CLK _13812_/D vssd1 vssd1 vccd1 vccd1 _13812_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14792_ _15645_/CLK _14792_/D vssd1 vssd1 vccd1 vccd1 _14792_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10955_ _11259_/S _10955_/B vssd1 vssd1 vccd1 vccd1 _10955_/Y sky130_fd_sc_hd__nor2_1
X_13743_ _14861_/CLK _13743_/D vssd1 vssd1 vccd1 vccd1 _13743_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13674_ _15606_/CLK _13674_/D vssd1 vssd1 vccd1 vccd1 _13674_/Q sky130_fd_sc_hd__dfxtp_1
X_10886_ _14918_/Q _15549_/Q _12320_/A vssd1 vssd1 vccd1 vccd1 _14918_/D sky130_fd_sc_hd__mux2_1
X_15413_ _15599_/CLK _15413_/D vssd1 vssd1 vccd1 vccd1 _15413_/Q sky130_fd_sc_hd__dfxtp_2
X_12625_ _13582_/Q _06861_/B _12624_/X _12647_/B vssd1 vssd1 vccd1 vccd1 _12625_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_169_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_633 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15344_ _15624_/CLK _15344_/D vssd1 vssd1 vccd1 vccd1 _15344_/Q sky130_fd_sc_hd__dfxtp_2
X_12556_ _12552_/X _12553_/X _12559_/A vssd1 vssd1 vccd1 vccd1 _12556_/X sky130_fd_sc_hd__mux2_1
XFILLER_89_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11507_ _11507_/A _11507_/B vssd1 vssd1 vccd1 vccd1 _11508_/B sky130_fd_sc_hd__or2_4
XFILLER_144_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15275_ _15275_/CLK _15275_/D vssd1 vssd1 vccd1 vccd1 _15275_/Q sky130_fd_sc_hd__dfxtp_1
X_12487_ _12483_/X _12484_/X _12490_/A vssd1 vssd1 vccd1 vccd1 _12487_/X sky130_fd_sc_hd__mux2_1
XFILLER_171_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11438_ _13229_/A _11476_/C vssd1 vssd1 vccd1 vccd1 _11439_/B sky130_fd_sc_hd__or2_4
X_14226_ _14420_/CLK _14226_/D vssd1 vssd1 vccd1 vccd1 _14226_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_137_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_246_clk clkbuf_5_4_0_clk/X vssd1 vssd1 vccd1 vccd1 _15212_/CLK sky130_fd_sc_hd__clkbuf_16
X_14157_ _15675_/CLK _14157_/D vssd1 vssd1 vccd1 vccd1 _14157_/Q sky130_fd_sc_hd__dfxtp_1
X_11369_ _11641_/S _11369_/B _11369_/C vssd1 vssd1 vccd1 vccd1 _11369_/X sky130_fd_sc_hd__or3_1
XFILLER_153_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13108_ _13029_/X _13044_/X _13114_/B1 _07488_/X vssd1 vssd1 vccd1 vccd1 _13108_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_140_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14088_ _15334_/CLK _14088_/D vssd1 vssd1 vccd1 vccd1 _14088_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13039_ _07500_/X _13039_/A2 _13038_/X _12944_/A vssd1 vssd1 vccd1 vccd1 _13039_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_21_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07600_ _07607_/A _07600_/B vssd1 vssd1 vccd1 vccd1 _07600_/Y sky130_fd_sc_hd__nand2_1
XFILLER_26_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08580_ _13781_/Q _08626_/S _08579_/X vssd1 vssd1 vccd1 vccd1 _13781_/D sky130_fd_sc_hd__o21a_1
XFILLER_66_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07531_ _14761_/Q _13440_/Q _07535_/S vssd1 vssd1 vccd1 vccd1 _13440_/D sky130_fd_sc_hd__mux2_1
XFILLER_50_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07462_ _14667_/Q _07474_/B _07482_/C vssd1 vssd1 vccd1 vccd1 _07462_/X sky130_fd_sc_hd__and3_1
XFILLER_50_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09201_ _09435_/A _09201_/B vssd1 vssd1 vccd1 vccd1 _09201_/X sky130_fd_sc_hd__or2_1
X_07393_ _13323_/A0 _13387_/Q _07481_/S vssd1 vssd1 vccd1 vccd1 _13387_/D sky130_fd_sc_hd__mux2_1
XFILLER_176_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09132_ _15660_/Q _13394_/Q _09132_/S vssd1 vssd1 vccd1 vccd1 _09132_/X sky130_fd_sc_hd__mux2_1
XFILLER_147_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09063_ _14526_/Q _14139_/Q _14171_/Q _14107_/Q _09230_/S _09234_/S1 vssd1 vssd1
+ vccd1 vccd1 _09063_/X sky130_fd_sc_hd__mux4_1
XFILLER_135_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08014_ _13569_/Q _08017_/D _13570_/Q vssd1 vssd1 vccd1 vccd1 _08014_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_135_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_237_clk clkbuf_5_5_0_clk/X vssd1 vssd1 vccd1 vccd1 _15202_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_144_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09965_ _11852_/A1 _14324_/Q _09991_/S vssd1 vssd1 vccd1 vccd1 _14324_/D sky130_fd_sc_hd__mux2_1
XFILLER_98_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08916_ _09546_/S1 _08914_/X _08915_/X vssd1 vssd1 vccd1 vccd1 _08920_/B sky130_fd_sc_hd__a21o_1
XFILLER_134_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09896_ _13349_/A0 _14258_/Q _09897_/S vssd1 vssd1 vccd1 vccd1 _14258_/D sky130_fd_sc_hd__mux2_1
XFILLER_97_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08847_ _13870_/Q _11879_/A1 _08851_/S vssd1 vssd1 vccd1 vccd1 _13870_/D sky130_fd_sc_hd__mux2_1
XFILLER_111_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08778_ _13125_/B _14613_/Q _13125_/A _08778_/D vssd1 vssd1 vccd1 vccd1 _08779_/C
+ sky130_fd_sc_hd__or4_1
XTAP_2804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07729_ _14752_/Q _07750_/A _07728_/Y _07987_/C1 vssd1 vssd1 vccd1 vccd1 _13495_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_2848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10740_ _15404_/Q _14772_/Q _10759_/S vssd1 vssd1 vccd1 vccd1 _14772_/D sky130_fd_sc_hd__mux2_1
XFILLER_129_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10671_ _15572_/Q _10706_/B vssd1 vssd1 vccd1 vccd1 _10671_/X sky130_fd_sc_hd__and2_1
XFILLER_159_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12410_ _12393_/X _12394_/X _12594_/S vssd1 vssd1 vccd1 vccd1 _12410_/X sky130_fd_sc_hd__mux2_1
XFILLER_22_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13390_ _15656_/CLK _13390_/D vssd1 vssd1 vccd1 vccd1 _13390_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_166_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12341_ _12324_/X _12325_/X _12536_/A vssd1 vssd1 vccd1 vccd1 _12341_/X sky130_fd_sc_hd__mux2_1
XFILLER_166_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15060_ _15067_/CLK _15060_/D vssd1 vssd1 vccd1 vccd1 _15060_/Q sky130_fd_sc_hd__dfxtp_4
X_12272_ _12255_/X _12256_/X _12582_/A vssd1 vssd1 vccd1 vccd1 _12272_/X sky130_fd_sc_hd__mux2_1
XFILLER_181_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14011_ _14083_/CLK _14011_/D vssd1 vssd1 vccd1 vccd1 _14011_/Q sky130_fd_sc_hd__dfxtp_1
X_11223_ _10528_/A _15011_/Q _11232_/S vssd1 vssd1 vccd1 vccd1 _15011_/D sky130_fd_sc_hd__mux2_1
XFILLER_49_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_228_clk clkbuf_5_6_0_clk/X vssd1 vssd1 vccd1 vccd1 _15510_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_153_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11154_ _14974_/Q _10984_/Y _11153_/X vssd1 vssd1 vccd1 vccd1 _14974_/D sky130_fd_sc_hd__a21o_1
XFILLER_136_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10105_ _14491_/Q _14739_/Q _10131_/S vssd1 vssd1 vccd1 vccd1 _14491_/D sky130_fd_sc_hd__mux2_1
XFILLER_110_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11085_ _11034_/Y _11036_/Y _11330_/A vssd1 vssd1 vccd1 vccd1 _11085_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10036_ _14393_/Q _11680_/A0 _10059_/S vssd1 vssd1 vccd1 vccd1 _14393_/D sky130_fd_sc_hd__mux2_1
X_14913_ _15544_/CLK _14913_/D vssd1 vssd1 vccd1 vccd1 _14913_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14844_ _15497_/CLK _14844_/D vssd1 vssd1 vccd1 vccd1 _14844_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14775_ _15592_/CLK _14775_/D vssd1 vssd1 vccd1 vccd1 _14775_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11987_ _13943_/Q _13685_/Q _12079_/S vssd1 vssd1 vccd1 vccd1 _11988_/B sky130_fd_sc_hd__mux2_1
XFILLER_32_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13726_ _15020_/CLK _13726_/D vssd1 vssd1 vccd1 vccd1 _13726_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10938_ _14953_/Q _10951_/B _10937_/Y _13226_/B vssd1 vssd1 vccd1 vccd1 _14953_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_143_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13657_ _14774_/CLK _13657_/D vssd1 vssd1 vccd1 vccd1 _13657_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10869_ _14901_/Q hold3/X _12906_/S vssd1 vssd1 vccd1 vccd1 _14901_/D sky130_fd_sc_hd__mux2_1
XFILLER_176_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12608_ _13970_/Q _13712_/Q _12612_/S vssd1 vssd1 vccd1 vccd1 _12609_/B sky130_fd_sc_hd__mux2_1
XPHY_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13588_ _15624_/CLK _13588_/D vssd1 vssd1 vccd1 vccd1 _13588_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_158_986 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15327_ _15670_/CLK _15327_/D vssd1 vssd1 vccd1 vccd1 _15327_/Q sky130_fd_sc_hd__dfxtp_2
X_12539_ _13967_/Q _13709_/Q _12541_/S vssd1 vssd1 vccd1 vccd1 _12540_/B sky130_fd_sc_hd__mux2_1
XFILLER_129_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15258_ _15666_/CLK _15258_/D vssd1 vssd1 vccd1 vccd1 _15258_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_172_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_219_clk clkbuf_5_18_0_clk/X vssd1 vssd1 vccd1 vccd1 _15517_/CLK sky130_fd_sc_hd__clkbuf_16
X_14209_ _15235_/CLK _14209_/D vssd1 vssd1 vccd1 vccd1 _14209_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_28_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15189_ _15666_/CLK _15189_/D vssd1 vssd1 vccd1 vccd1 _15189_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_126_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout408 _11641_/S vssd1 vssd1 vccd1 vccd1 _11474_/S sky130_fd_sc_hd__buf_4
XFILLER_63_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout419 _10576_/X vssd1 vssd1 vccd1 vccd1 _10733_/B1 sky130_fd_sc_hd__buf_12
XFILLER_141_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09750_ _14118_/Q _13338_/A0 _09762_/S vssd1 vssd1 vccd1 vccd1 _14118_/D sky130_fd_sc_hd__mux2_1
X_06962_ _14491_/Q _06743_/Y _14490_/Q _06746_/Y _06961_/X vssd1 vssd1 vccd1 vccd1
+ _06963_/B sky130_fd_sc_hd__o221a_1
XFILLER_79_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08701_ _13579_/Q _08667_/X _08668_/X _13578_/Q _08700_/X vssd1 vssd1 vccd1 vccd1
+ _08701_/X sky130_fd_sc_hd__a221o_1
X_09681_ _14052_/Q _11761_/A0 _09695_/S vssd1 vssd1 vccd1 vccd1 _14052_/D sky130_fd_sc_hd__mux2_1
X_06893_ _15383_/Q _07595_/A _15382_/Q _07595_/B vssd1 vssd1 vccd1 vccd1 _06910_/S
+ sky130_fd_sc_hd__o22a_1
XFILLER_39_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_366 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08632_ _08722_/A _08632_/B _08632_/C vssd1 vssd1 vccd1 vccd1 _08632_/X sky130_fd_sc_hd__or3_1
XFILLER_82_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08563_ _13568_/Q _08747_/A2 _08747_/B1 _13504_/Q vssd1 vssd1 vccd1 vccd1 _08563_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_35_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07514_ _14744_/Q _13423_/Q _07529_/S vssd1 vssd1 vccd1 vccd1 _13423_/D sky130_fd_sc_hd__mux2_1
XFILLER_35_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08494_ _09512_/S _08494_/B vssd1 vssd1 vccd1 vccd1 _08494_/Y sky130_fd_sc_hd__nor2_8
XFILLER_120_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_199 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07445_ _13336_/A0 _13400_/Q _07501_/S vssd1 vssd1 vccd1 vccd1 _13400_/D sky130_fd_sc_hd__mux2_1
XFILLER_50_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07376_ _14734_/Q _07375_/X _07500_/S vssd1 vssd1 vccd1 vccd1 _07376_/X sky130_fd_sc_hd__mux2_8
X_09115_ _06676_/A _09104_/X _09113_/X _09114_/X vssd1 vssd1 vccd1 vccd1 _09115_/X
+ sky130_fd_sc_hd__o22a_2
XFILLER_135_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09046_ _09406_/S1 _09044_/X _09045_/X vssd1 vssd1 vccd1 vccd1 _09046_/X sky130_fd_sc_hd__a21o_1
XFILLER_164_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_79 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09948_ _11868_/A1 _14308_/Q _09958_/S vssd1 vssd1 vccd1 vccd1 _14308_/D sky130_fd_sc_hd__mux2_1
XTAP_4003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09879_ _13078_/B2 _14241_/Q _09892_/S vssd1 vssd1 vccd1 vccd1 _14241_/D sky130_fd_sc_hd__mux2_1
XTAP_4047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11910_ _14519_/Q _14132_/Q _14164_/Q _14100_/Q _08405_/A _12563_/A vssd1 vssd1 vccd1
+ vccd1 _11910_/X sky130_fd_sc_hd__mux4_1
XTAP_3335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12890_ _15418_/Q _15603_/Q _12929_/S vssd1 vssd1 vccd1 vccd1 _15418_/D sky130_fd_sc_hd__mux2_1
XTAP_3346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_122 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11841_ _15263_/Q _11874_/A1 _11850_/S vssd1 vssd1 vccd1 vccd1 _15263_/D sky130_fd_sc_hd__mux2_1
XTAP_2634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_572 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11772_ _11847_/A1 _15200_/Q _11775_/S vssd1 vssd1 vccd1 vccd1 _15200_/D sky130_fd_sc_hd__mux2_1
X_14560_ _15298_/CLK _14560_/D vssd1 vssd1 vccd1 vccd1 _14560_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13511_ _15372_/CLK _13511_/D vssd1 vssd1 vccd1 vccd1 _13511_/Q sky130_fd_sc_hd__dfxtp_2
X_10723_ _15040_/Q _10602_/B _10722_/X vssd1 vssd1 vccd1 vccd1 _10723_/X sky130_fd_sc_hd__a21o_1
XFILLER_186_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14491_ _15399_/CLK _14491_/D vssd1 vssd1 vccd1 vccd1 _14491_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_13_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10654_ _10651_/X _10652_/X _10653_/X _10714_/A2 _15058_/Q vssd1 vssd1 vccd1 vccd1
+ _10654_/X sky130_fd_sc_hd__o32a_2
XFILLER_9_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13442_ _14493_/CLK _13442_/D vssd1 vssd1 vccd1 vccd1 _13442_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_155_912 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_900 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13373_ _14476_/Q vssd1 vssd1 vccd1 vccd1 _14476_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_127_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10585_ _14735_/Q _10584_/X _10730_/S vssd1 vssd1 vccd1 vccd1 _14735_/D sky130_fd_sc_hd__mux2_1
XFILLER_103_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15112_ _15649_/CLK _15112_/D vssd1 vssd1 vccd1 vccd1 _15112_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_155_967 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12324_ _14537_/Q _14150_/Q _14182_/Q _14118_/Q _12543_/S _12544_/A vssd1 vssd1 vccd1
+ vccd1 _12324_/X sky130_fd_sc_hd__mux4_1
XFILLER_186_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12255_ _14534_/Q _14147_/Q _14179_/Q _14115_/Q _12269_/S _12268_/A vssd1 vssd1 vccd1
+ vccd1 _12255_/X sky130_fd_sc_hd__mux4_1
X_15043_ _15046_/CLK _15043_/D vssd1 vssd1 vccd1 vccd1 _15043_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_119_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11206_ _10555_/D _14995_/Q _11237_/S vssd1 vssd1 vccd1 vccd1 _14995_/D sky130_fd_sc_hd__mux2_1
XFILLER_107_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12186_ _14531_/Q _14144_/Q _14176_/Q _14112_/Q _12472_/S _12465_/S1 vssd1 vssd1
+ vccd1 vccd1 _12186_/X sky130_fd_sc_hd__mux4_1
XFILLER_122_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11137_ _11129_/A _11031_/A _11136_/X _08233_/B vssd1 vssd1 vccd1 vccd1 _11137_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_95_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11068_ _11088_/S _10996_/B _11307_/A vssd1 vssd1 vccd1 vccd1 _11068_/X sky130_fd_sc_hd__a21o_1
XFILLER_48_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_83 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10019_ _11873_/A1 _14377_/Q _10029_/S vssd1 vssd1 vccd1 vccd1 _14377_/D sky130_fd_sc_hd__mux2_1
XFILLER_110_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14827_ _15645_/CLK _14827_/D vssd1 vssd1 vccd1 vccd1 _14827_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14758_ _15607_/CLK _14758_/D vssd1 vssd1 vccd1 vccd1 _14758_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_60_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13709_ _15259_/CLK _13709_/D vssd1 vssd1 vccd1 vccd1 _13709_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_177_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14689_ _15592_/CLK _14689_/D vssd1 vssd1 vccd1 vccd1 _14689_/Q sky130_fd_sc_hd__dfxtp_1
X_07230_ _07205_/X _07230_/B _07230_/C _07230_/D vssd1 vssd1 vccd1 vccd1 _07230_/X
+ sky130_fd_sc_hd__and4b_1
X_07161_ _07163_/A _07161_/B vssd1 vssd1 vccd1 vccd1 _07161_/X sky130_fd_sc_hd__and2_4
XFILLER_9_771 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_956 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07092_ _07091_/X _14763_/Q _07098_/S vssd1 vssd1 vccd1 vccd1 _13609_/D sky130_fd_sc_hd__mux2_1
XFILLER_133_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout205 _09696_/X vssd1 vssd1 vccd1 vccd1 _09723_/S sky130_fd_sc_hd__buf_12
XFILLER_87_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout216 _08853_/Y vssd1 vssd1 vccd1 vccd1 _08885_/S sky130_fd_sc_hd__buf_12
XFILLER_101_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09802_ _14168_/Q _13324_/A0 _09828_/S vssd1 vssd1 vccd1 vccd1 _14168_/D sky130_fd_sc_hd__mux2_1
XFILLER_87_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout227 _07676_/A vssd1 vssd1 vccd1 vccd1 _07777_/A sky130_fd_sc_hd__buf_6
Xfanout238 _07004_/X vssd1 vssd1 vccd1 vccd1 _07077_/S sky130_fd_sc_hd__buf_12
X_07994_ _14757_/Q _07971_/A _07993_/Y vssd1 vssd1 vccd1 vccd1 _13564_/D sky130_fd_sc_hd__o21a_1
Xfanout249 _08521_/Y vssd1 vssd1 vccd1 vccd1 _08750_/A2 sky130_fd_sc_hd__buf_12
XFILLER_115_38 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09733_ _14101_/Q _13321_/A0 _09762_/S vssd1 vssd1 vccd1 vccd1 _14101_/D sky130_fd_sc_hd__mux2_1
X_06945_ _06945_/A vssd1 vssd1 vccd1 vccd1 _06945_/Y sky130_fd_sc_hd__inv_2
XFILLER_86_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09664_ _14035_/Q _13319_/A0 _09690_/S vssd1 vssd1 vccd1 vccd1 _14035_/D sky130_fd_sc_hd__mux2_1
X_06876_ _06692_/Y _13506_/Q _06882_/A _06875_/X _06879_/C vssd1 vssd1 vccd1 vccd1
+ _06877_/B sky130_fd_sc_hd__o221a_1
XFILLER_54_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_5_19_0_clk clkbuf_4_9_0_clk/X vssd1 vssd1 vccd1 vccd1 clkbuf_5_19_0_clk/X
+ sky130_fd_sc_hd__clkbuf_8
X_08615_ _13464_/Q _08684_/A2 _08693_/B1 _13631_/Q _08614_/X vssd1 vssd1 vccd1 vccd1
+ _08619_/B sky130_fd_sc_hd__a221o_1
XFILLER_131_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09595_ _11743_/C _14714_/Q _14716_/Q vssd1 vssd1 vccd1 vccd1 _09696_/B sky130_fd_sc_hd__or3b_4
XFILLER_83_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08546_ _13776_/Q _08573_/S _08542_/X _08545_/X vssd1 vssd1 vccd1 vccd1 _13776_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_23_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08477_ _14597_/Q _08756_/B _08477_/C vssd1 vssd1 vccd1 vccd1 _08477_/X sky130_fd_sc_hd__and3_2
XFILLER_126_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07428_ _14747_/Q _07427_/X _07480_/S vssd1 vssd1 vccd1 vccd1 _07428_/X sky130_fd_sc_hd__mux2_8
XFILLER_156_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_383 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_772 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07359_ _07195_/Y _07197_/B _07231_/C _07358_/Y _15529_/Q vssd1 vssd1 vccd1 vccd1
+ _07359_/X sky130_fd_sc_hd__o221a_1
XFILLER_6_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10370_ _10520_/A1 _13797_/Q _13765_/Q _10520_/B2 vssd1 vssd1 vccd1 vccd1 _10370_/X
+ sky130_fd_sc_hd__a22o_2
XFILLER_152_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09029_ _13881_/Q _09522_/A2 _09519_/B1 _14396_/Q _08507_/A vssd1 vssd1 vccd1 vccd1
+ _09029_/X sky130_fd_sc_hd__a221o_1
XFILLER_156_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12040_ _12592_/A1 _12039_/X _06670_/A vssd1 vssd1 vccd1 vccd1 _12040_/X sky130_fd_sc_hd__a21o_1
XFILLER_85_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13991_ _15293_/CLK _13991_/D vssd1 vssd1 vccd1 vccd1 _13991_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_93_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12942_ _08405_/D _13318_/C _09662_/B _08405_/A _12941_/Y vssd1 vssd1 vccd1 vccd1
+ _12943_/C sky130_fd_sc_hd__a221o_1
XFILLER_86_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15661_ _15661_/CLK _15661_/D vssd1 vssd1 vccd1 vccd1 _15661_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_73_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_110 input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12873_ _15401_/Q _15586_/Q _12932_/S vssd1 vssd1 vccd1 vccd1 _15401_/D sky130_fd_sc_hd__mux2_1
XTAP_3176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_121 _07117_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_132 _15344_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14612_ _14612_/CLK _14612_/D vssd1 vssd1 vccd1 vccd1 _14612_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_2453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11824_ _15246_/Q _11857_/A1 _11850_/S vssd1 vssd1 vccd1 vccd1 _15246_/D sky130_fd_sc_hd__mux2_1
XTAP_2464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15592_ _15592_/CLK _15592_/D vssd1 vssd1 vccd1 vccd1 _15592_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14543_ _15674_/CLK _14543_/D vssd1 vssd1 vccd1 vccd1 _14543_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11755_ _13330_/A0 _15183_/Q _11774_/S vssd1 vssd1 vccd1 vccd1 _15183_/D sky130_fd_sc_hd__mux2_1
XFILLER_14_564 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10706_ _15579_/Q _10706_/B vssd1 vssd1 vccd1 vccd1 _10706_/X sky130_fd_sc_hd__and2_1
XFILLER_159_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14474_ _15192_/CLK _14474_/D vssd1 vssd1 vccd1 vccd1 _14474_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_174_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11686_ _13328_/A0 _15117_/Q _11703_/S vssd1 vssd1 vccd1 vccd1 _15117_/D sky130_fd_sc_hd__mux2_1
X_13425_ _15354_/CLK _13425_/D vssd1 vssd1 vccd1 vccd1 _13425_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10637_ _15006_/Q _10717_/A2 _10652_/B _13725_/Q _10717_/C1 vssd1 vssd1 vccd1 vccd1
+ _10637_/X sky130_fd_sc_hd__a221o_1
XFILLER_155_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13356_ _14459_/Q vssd1 vssd1 vccd1 vccd1 _14459_/D sky130_fd_sc_hd__clkbuf_2
X_10568_ _10581_/A _10569_/B vssd1 vssd1 vccd1 vccd1 _10568_/X sky130_fd_sc_hd__and2_2
XFILLER_128_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12307_ _12615_/B1 _12304_/X _12616_/C1 vssd1 vssd1 vccd1 vccd1 _12307_/X sky130_fd_sc_hd__o21a_1
X_10499_ _10507_/A1 _13753_/Q _15419_/Q _10515_/B2 vssd1 vssd1 vccd1 vccd1 _10499_/X
+ sky130_fd_sc_hd__a22o_1
X_13287_ _12629_/X _15619_/Q _13291_/S vssd1 vssd1 vccd1 vccd1 _15619_/D sky130_fd_sc_hd__mux2_1
XFILLER_142_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15026_ _15584_/CLK _15026_/D vssd1 vssd1 vccd1 vccd1 _15026_/Q sky130_fd_sc_hd__dfxtp_1
X_12238_ _08453_/A _12235_/X _08451_/A vssd1 vssd1 vccd1 vccd1 _12238_/X sky130_fd_sc_hd__o21a_1
XFILLER_170_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12169_ _12500_/B1 _12166_/X _12501_/C1 vssd1 vssd1 vccd1 vccd1 _12169_/X sky130_fd_sc_hd__o21a_1
XFILLER_96_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06730_ _14497_/Q vssd1 vssd1 vccd1 vccd1 _06730_/Y sky130_fd_sc_hd__clkinv_2
Xinput5 ext_read_data[13] vssd1 vssd1 vccd1 vccd1 input5/X sky130_fd_sc_hd__clkbuf_8
XFILLER_36_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_1050 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06661_ _14900_/Q vssd1 vssd1 vccd1 vccd1 _06661_/Y sky130_fd_sc_hd__inv_2
XFILLER_91_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08400_ _13140_/S _08469_/A _08400_/C vssd1 vssd1 vccd1 vccd1 _08400_/X sky130_fd_sc_hd__or3_1
X_09380_ _14090_/Q _13123_/B _08508_/Y _14058_/Q _09532_/A vssd1 vssd1 vccd1 vccd1
+ _09380_/X sky130_fd_sc_hd__a221o_1
XFILLER_80_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08331_ _08259_/Y _08320_/Y _08330_/X _11329_/A vssd1 vssd1 vccd1 vccd1 _08331_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_51_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_322 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08262_ _11349_/B _13159_/B vssd1 vssd1 vccd1 vccd1 _08262_/Y sky130_fd_sc_hd__nand2_1
XFILLER_20_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07213_ _13934_/Q _15521_/Q _07334_/S vssd1 vssd1 vccd1 vccd1 _07213_/X sky130_fd_sc_hd__mux2_8
X_08193_ _13684_/Q _11680_/A0 _08216_/S vssd1 vssd1 vccd1 vccd1 _13684_/D sky130_fd_sc_hd__mux2_1
XFILLER_146_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07144_ _14852_/Q _14844_/Q _08094_/S vssd1 vssd1 vccd1 vccd1 _07144_/X sky130_fd_sc_hd__mux2_1
XFILLER_69_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_775 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07075_ _14637_/Q _14669_/Q _07078_/S vssd1 vssd1 vccd1 vccd1 _07075_/X sky130_fd_sc_hd__mux2_1
XFILLER_145_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_13 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_5_2_0_clk clkbuf_5_3_0_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_5_2_0_clk/X sky130_fd_sc_hd__clkbuf_8
XFILLER_75_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07977_ _13560_/Q _07984_/D vssd1 vssd1 vccd1 vccd1 _07981_/B sky130_fd_sc_hd__nand2_1
XFILLER_75_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09716_ _11838_/A1 _14086_/Q _09728_/S vssd1 vssd1 vccd1 vccd1 _14086_/D sky130_fd_sc_hd__mux2_1
X_06928_ _06687_/Y _13476_/Q _06704_/Y _13469_/Q _06883_/X vssd1 vssd1 vccd1 vccd1
+ _06931_/A sky130_fd_sc_hd__o221a_1
XFILLER_28_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09647_ _14020_/Q _11761_/A0 _09661_/S vssd1 vssd1 vccd1 vccd1 _14020_/D sky130_fd_sc_hd__mux2_1
XFILLER_82_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06859_ _14730_/Q _14729_/Q vssd1 vssd1 vccd1 vccd1 _06861_/B sky130_fd_sc_hd__and2_4
XFILLER_27_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09578_ _13954_/Q _13082_/B2 _09589_/S vssd1 vssd1 vccd1 vccd1 _13954_/D sky130_fd_sc_hd__mux2_1
XTAP_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08529_ _13125_/B _08529_/B vssd1 vssd1 vccd1 vccd1 _08530_/B sky130_fd_sc_hd__or2_4
XFILLER_169_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11540_ _13217_/B _11541_/B vssd1 vssd1 vccd1 vccd1 _11542_/A sky130_fd_sc_hd__or2_2
XFILLER_184_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11471_ _11471_/A _11471_/B vssd1 vssd1 vccd1 vccd1 _11505_/B sky130_fd_sc_hd__nor2_1
XFILLER_167_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13210_ _13208_/Y _13209_/X _15570_/Q _13241_/A2 vssd1 vssd1 vccd1 vccd1 _15570_/D
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_13_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10422_ _07227_/A _10481_/B _10421_/X vssd1 vssd1 vccd1 vccd1 _11349_/C sky130_fd_sc_hd__a21o_4
X_14190_ _15676_/CLK _14190_/D vssd1 vssd1 vccd1 vccd1 _14190_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10353_ _07280_/A _10360_/B _10352_/X vssd1 vssd1 vccd1 vccd1 _11496_/A sky130_fd_sc_hd__a21oi_4
X_13141_ _08530_/B _08779_/B _15538_/Q _13129_/A vssd1 vssd1 vccd1 vccd1 _15538_/D
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_174_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13072_ _12975_/X _13104_/A2 _13104_/B1 _13072_/B2 vssd1 vssd1 vccd1 vccd1 _13072_/X
+ sky130_fd_sc_hd__a22o_1
X_10284_ _14669_/Q _14822_/Q _10285_/S vssd1 vssd1 vccd1 vccd1 _14669_/D sky130_fd_sc_hd__mux2_1
XFILLER_152_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12023_ _14234_/Q _14266_/Q _14298_/Q _14330_/Q _12079_/S _12080_/A vssd1 vssd1 vccd1
+ vccd1 _12023_/X sky130_fd_sc_hd__mux4_1
XFILLER_78_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout580 _08405_/B vssd1 vssd1 vccd1 vccd1 _12615_/B1 sky130_fd_sc_hd__buf_12
XFILLER_76_63 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout591 _14599_/Q vssd1 vssd1 vccd1 vccd1 _12486_/S1 sky130_fd_sc_hd__buf_6
XFILLER_120_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13974_ _14462_/CLK _13974_/D vssd1 vssd1 vccd1 vccd1 _13974_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_1016 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12925_ _15453_/Q _15639_/Q _12929_/S vssd1 vssd1 vccd1 vccd1 _15453_/D sky130_fd_sc_hd__mux2_1
XFILLER_73_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15644_ _15644_/CLK _15644_/D vssd1 vssd1 vccd1 vccd1 _15644_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12856_ _14750_/Q _15384_/Q _12866_/S vssd1 vssd1 vccd1 vccd1 _15384_/D sky130_fd_sc_hd__mux2_1
XFILLER_33_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11807_ _15230_/Q _13340_/A0 _11817_/S vssd1 vssd1 vccd1 vccd1 _15230_/D sky130_fd_sc_hd__mux2_1
XTAP_2294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15575_ _15579_/CLK _15575_/D vssd1 vssd1 vccd1 vccd1 _15575_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12787_ _06861_/B _12786_/X _12785_/X _12764_/S vssd1 vssd1 vccd1 vccd1 _12787_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14526_ _15657_/CLK _14526_/D vssd1 vssd1 vccd1 vccd1 _14526_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_42_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11738_ _15167_/Q _11879_/A1 _11742_/S vssd1 vssd1 vccd1 vccd1 _15167_/D sky130_fd_sc_hd__mux2_1
XFILLER_31_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14457_ _15244_/CLK _14457_/D vssd1 vssd1 vccd1 vccd1 _14457_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_175_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11669_ _13344_/A0 _15101_/Q _11670_/S vssd1 vssd1 vccd1 vccd1 _15101_/D sky130_fd_sc_hd__mux2_1
X_13408_ _15674_/CLK _13408_/D vssd1 vssd1 vccd1 vccd1 _13408_/Q sky130_fd_sc_hd__dfxtp_1
X_14388_ _15619_/CLK _14388_/D vssd1 vssd1 vccd1 vccd1 _14388_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_183_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13339_ _13339_/A0 _15669_/Q _13350_/S vssd1 vssd1 vccd1 vccd1 _15669_/D sky130_fd_sc_hd__mux2_1
XFILLER_51_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15009_ _15570_/CLK _15009_/D vssd1 vssd1 vccd1 vccd1 _15009_/Q sky130_fd_sc_hd__dfxtp_1
X_07900_ _13540_/Q _13539_/Q _07900_/C _07900_/D vssd1 vssd1 vccd1 vccd1 _07913_/D
+ sky130_fd_sc_hd__and4_2
XFILLER_29_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08880_ _13901_/Q _13104_/B2 _08880_/S vssd1 vssd1 vccd1 vccd1 _13901_/D sky130_fd_sc_hd__mux2_1
X_07831_ _14746_/Q _07830_/A _07830_/Y _12788_/C1 vssd1 vssd1 vccd1 vccd1 _13521_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_116_1055 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07762_ _07760_/Y _07764_/B _07777_/A vssd1 vssd1 vccd1 vccd1 _07762_/Y sky130_fd_sc_hd__o21ai_1
X_09501_ _08494_/B _08519_/B _09500_/X _13049_/A1 vssd1 vssd1 vccd1 vccd1 _09501_/X
+ sky130_fd_sc_hd__a31o_1
X_06713_ _13497_/Q vssd1 vssd1 vccd1 vccd1 _06713_/Y sky130_fd_sc_hd__inv_2
XFILLER_38_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07693_ _13485_/Q _07717_/A _13486_/Q vssd1 vssd1 vccd1 vccd1 _07693_/Y sky130_fd_sc_hd__a21oi_1
X_09432_ _09430_/X _09431_/X _12481_/A _09421_/X vssd1 vssd1 vccd1 vccd1 _09432_/X
+ sky130_fd_sc_hd__o211a_1
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09363_ _15130_/Q _15098_/Q _15671_/Q _13405_/Q _09521_/S _09523_/A1 vssd1 vssd1
+ vccd1 vccd1 _09363_/X sky130_fd_sc_hd__mux4_1
XFILLER_12_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_1083 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08314_ _11037_/A _11419_/A vssd1 vssd1 vccd1 vccd1 _10986_/A sky130_fd_sc_hd__nor2_1
XFILLER_166_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09294_ _08519_/A _09292_/X _09293_/X vssd1 vssd1 vccd1 vccd1 _09294_/X sky130_fd_sc_hd__a21o_1
XANTENNA_10 _10624_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_21 _13787_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_32 _14750_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_43 input20/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08245_ _10515_/B2 _15430_/Q _13774_/Q _10507_/A1 vssd1 vssd1 vccd1 vccd1 _08245_/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA_54 _07164_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_65 _07127_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_76 _07155_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_87 _13072_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_98 _10634_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08176_ _13675_/Q _10285_/S _08155_/X _08175_/X vssd1 vssd1 vccd1 vccd1 _13675_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_107_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07127_ _07131_/A _07127_/B vssd1 vssd1 vccd1 vccd1 _07127_/X sky130_fd_sc_hd__and2_4
XFILLER_119_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07058_ _07057_/X _13598_/Q _12764_/S vssd1 vssd1 vccd1 vccd1 _07058_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_714 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10971_ _11258_/B _11242_/A vssd1 vssd1 vccd1 vccd1 _10971_/Y sky130_fd_sc_hd__nor2_1
XFILLER_90_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12710_ _15350_/Q _12710_/B vssd1 vssd1 vccd1 vccd1 _12711_/B sky130_fd_sc_hd__or2_1
XFILLER_15_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13690_ _15184_/CLK _13690_/D vssd1 vssd1 vccd1 vccd1 _13690_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_147 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12641_ _12743_/A _12641_/B vssd1 vssd1 vccd1 vccd1 _12641_/X sky130_fd_sc_hd__or2_1
XFILLER_70_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15360_ _15378_/CLK _15360_/D vssd1 vssd1 vccd1 vccd1 _15360_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_168_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12572_ _12595_/A1 _12571_/X _12570_/X _12618_/C1 vssd1 vssd1 vccd1 vccd1 _12573_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_50_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14311_ _15275_/CLK _14311_/D vssd1 vssd1 vccd1 vccd1 _14311_/Q sky130_fd_sc_hd__dfxtp_1
X_11523_ _11501_/A _11515_/B _11512_/X vssd1 vssd1 vccd1 vccd1 _11523_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_156_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15291_ _15291_/CLK _15291_/D vssd1 vssd1 vccd1 vccd1 _15291_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14242_ _14468_/CLK _14242_/D vssd1 vssd1 vccd1 vccd1 _14242_/Q sky130_fd_sc_hd__dfxtp_1
X_11454_ _11476_/A _11476_/B _11476_/C _13229_/A vssd1 vssd1 vccd1 vccd1 _11455_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_171_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10405_ _11362_/B _13162_/B _13165_/B _11371_/A _10404_/X vssd1 vssd1 vccd1 vccd1
+ _10405_/X sky130_fd_sc_hd__o221a_1
XFILLER_164_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14173_ _15674_/CLK _14173_/D vssd1 vssd1 vccd1 vccd1 _14173_/Q sky130_fd_sc_hd__dfxtp_1
X_11385_ _11423_/A _11423_/B vssd1 vssd1 vccd1 vccd1 _11386_/B sky130_fd_sc_hd__and2_1
XFILLER_178_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13124_ _08668_/B _08724_/C _08532_/B _13123_/Y vssd1 vssd1 vccd1 vccd1 _13124_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_139_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10336_ _14721_/Q _14914_/Q _10343_/S vssd1 vssd1 vccd1 vccd1 _14721_/D sky130_fd_sc_hd__mux2_1
XFILLER_180_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_406 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_4_9_0_clk clkbuf_4_9_0_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_9_0_clk/X sky130_fd_sc_hd__clkbuf_8
XTAP_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13055_ _15495_/Q _13139_/S _13042_/A _13054_/X vssd1 vssd1 vccd1 vccd1 _15495_/D
+ sky130_fd_sc_hd__a22o_1
X_10267_ _14652_/Q _14805_/Q _10343_/S vssd1 vssd1 vccd1 vccd1 _14652_/D sky130_fd_sc_hd__mux2_1
XFILLER_121_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12006_ _15278_/Q _15246_/Q _15214_/Q _15145_/Q _12407_/S _12406_/A vssd1 vssd1 vccd1
+ vccd1 _12007_/B sky130_fd_sc_hd__mux4_1
XFILLER_78_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10198_ input1/X _14583_/Q _13284_/S vssd1 vssd1 vccd1 vccd1 _14583_/D sky130_fd_sc_hd__mux2_1
XFILLER_94_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13957_ _15094_/CLK _13957_/D vssd1 vssd1 vccd1 vccd1 _13957_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_46_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_1072 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12908_ _15436_/Q _15622_/Q _12910_/S vssd1 vssd1 vccd1 vccd1 _15436_/D sky130_fd_sc_hd__mux2_1
XFILLER_35_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13888_ _15331_/CLK _13888_/D vssd1 vssd1 vccd1 vccd1 _13888_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_179_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15627_ _15632_/CLK _15627_/D vssd1 vssd1 vccd1 vccd1 _15627_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12839_ _14717_/Q _12839_/B _10099_/C vssd1 vssd1 vccd1 vccd1 _12839_/X sky130_fd_sc_hd__or3b_4
XTAP_2091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15558_ _15558_/CLK _15558_/D vssd1 vssd1 vccd1 vccd1 _15558_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_483 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14509_ _14510_/CLK _14509_/D vssd1 vssd1 vccd1 vccd1 _14509_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_147_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15489_ _15489_/CLK _15489_/D vssd1 vssd1 vccd1 vccd1 _15489_/Q sky130_fd_sc_hd__dfxtp_1
X_08030_ _12647_/B _12763_/S vssd1 vssd1 vccd1 vccd1 _08030_/Y sky130_fd_sc_hd__nor2_8
Xinput30 ext_read_data[7] vssd1 vssd1 vccd1 vccd1 input30/X sky130_fd_sc_hd__buf_4
XFILLER_162_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09981_ _11868_/A1 _14340_/Q _09991_/S vssd1 vssd1 vccd1 vccd1 _14340_/D sky130_fd_sc_hd__mux2_1
XFILLER_107_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08932_ _14230_/Q _14262_/Q _14294_/Q _14326_/Q _09484_/S _08519_/A vssd1 vssd1 vccd1
+ vccd1 _08932_/X sky130_fd_sc_hd__mux4_1
XFILLER_88_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08863_ _13884_/Q _13328_/A0 _08880_/S vssd1 vssd1 vccd1 vccd1 _13884_/D sky130_fd_sc_hd__mux2_1
XFILLER_69_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07814_ _13516_/Q _13515_/Q _07813_/D _13517_/Q vssd1 vssd1 vccd1 vccd1 _07815_/B
+ sky130_fd_sc_hd__a31o_1
XTAP_3709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08794_ _11861_/A1 _13820_/Q _08811_/S vssd1 vssd1 vccd1 vccd1 _13820_/D sky130_fd_sc_hd__mux2_1
XFILLER_85_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07745_ _13499_/Q _07746_/C _13500_/Q vssd1 vssd1 vccd1 vccd1 _07745_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_42_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07676_ _07676_/A _07676_/B vssd1 vssd1 vccd1 vccd1 _07676_/Y sky130_fd_sc_hd__nand2_1
XFILLER_73_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09415_ _15298_/Q _15266_/Q _15234_/Q _15165_/Q _09444_/S _09446_/A1 vssd1 vssd1
+ vccd1 vccd1 _09415_/X sky130_fd_sc_hd__mux4_1
XFILLER_52_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09346_ _13134_/A _09346_/B _09346_/C vssd1 vssd1 vccd1 vccd1 _09346_/X sky130_fd_sc_hd__and3_1
XFILLER_21_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09277_ _15667_/Q _13401_/Q _09557_/S vssd1 vssd1 vccd1 vccd1 _09277_/X sky130_fd_sc_hd__mux2_1
XFILLER_166_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08228_ _07339_/X _10457_/A2 _08226_/X vssd1 vssd1 vccd1 vccd1 _08228_/X sky130_fd_sc_hd__a21o_2
XFILLER_20_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08159_ _08185_/A _08159_/B vssd1 vssd1 vccd1 vccd1 _08159_/X sky130_fd_sc_hd__and2_1
XFILLER_10_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11170_ _13251_/A _11380_/A _13251_/B _10984_/Y vssd1 vssd1 vccd1 vccd1 _11170_/X
+ sky130_fd_sc_hd__a31o_4
XFILLER_134_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10121_ _14507_/Q _14755_/Q _10124_/S vssd1 vssd1 vccd1 vccd1 _14507_/D sky130_fd_sc_hd__mux2_1
XFILLER_106_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10052_ _14409_/Q _13338_/A0 _10064_/S vssd1 vssd1 vccd1 vccd1 _14409_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14860_ _15500_/CLK _14860_/D vssd1 vssd1 vccd1 vccd1 _14860_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13811_ _15209_/CLK _13811_/D vssd1 vssd1 vccd1 vccd1 _13811_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_180_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14791_ _15606_/CLK _14791_/D vssd1 vssd1 vccd1 vccd1 _14791_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_28_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13742_ _14863_/CLK _13742_/D vssd1 vssd1 vccd1 vccd1 _14927_/D sky130_fd_sc_hd__dfxtp_4
X_10954_ _11023_/A wire360/X _11317_/A vssd1 vssd1 vccd1 vccd1 _10955_/B sky130_fd_sc_hd__o21bai_1
XFILLER_71_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_75 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13673_ _15606_/CLK _13673_/D vssd1 vssd1 vccd1 vccd1 _13673_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_43_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_191_clk clkbuf_5_20_0_clk/X vssd1 vssd1 vccd1 vccd1 _15292_/CLK sky130_fd_sc_hd__clkbuf_16
X_10885_ _14917_/Q _15548_/Q _13134_/A vssd1 vssd1 vccd1 vccd1 _14917_/D sky130_fd_sc_hd__mux2_1
X_15412_ _15632_/CLK _15412_/D vssd1 vssd1 vccd1 vccd1 _15412_/Q sky130_fd_sc_hd__dfxtp_2
X_12624_ _15045_/Q _12834_/B _12785_/B _12623_/Y vssd1 vssd1 vccd1 vccd1 _12624_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_106_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15343_ _15647_/CLK _15343_/D vssd1 vssd1 vccd1 vccd1 _15343_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_12_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12555_ _15137_/Q _15105_/Q _15678_/Q _13412_/Q _12568_/S _12567_/A vssd1 vssd1 vccd1
+ vccd1 _12555_/X sky130_fd_sc_hd__mux4_1
XFILLER_185_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11506_ _11464_/B _11464_/C _11505_/X vssd1 vssd1 vccd1 vccd1 _11507_/B sky130_fd_sc_hd__o21a_1
X_15274_ _15676_/CLK _15274_/D vssd1 vssd1 vccd1 vccd1 _15274_/Q sky130_fd_sc_hd__dfxtp_1
X_12486_ _15134_/Q _15102_/Q _15675_/Q _13409_/Q _12499_/S _12486_/S1 vssd1 vssd1
+ vccd1 vccd1 _12486_/X sky130_fd_sc_hd__mux4_1
XFILLER_138_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_892 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14225_ _14225_/CLK _14225_/D vssd1 vssd1 vccd1 vccd1 _14225_/Q sky130_fd_sc_hd__dfxtp_1
X_11437_ _11437_/A _11437_/B _11437_/C vssd1 vssd1 vccd1 vccd1 _11476_/C sky130_fd_sc_hd__and3_2
XFILLER_138_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14156_ _15674_/CLK _14156_/D vssd1 vssd1 vccd1 vccd1 _14156_/Q sky130_fd_sc_hd__dfxtp_1
X_11368_ _11368_/A _11368_/B vssd1 vssd1 vccd1 vccd1 _11369_/C sky130_fd_sc_hd__and2_1
XFILLER_98_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13107_ _15521_/Q _13129_/A _13042_/A _13106_/X vssd1 vssd1 vccd1 vccd1 _15521_/D
+ sky130_fd_sc_hd__a22o_1
X_10319_ _14704_/Q _14889_/Q _10715_/S vssd1 vssd1 vccd1 vccd1 _14704_/D sky130_fd_sc_hd__mux2_1
XTAP_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14087_ _15292_/CLK _14087_/D vssd1 vssd1 vccd1 vccd1 _14087_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11299_ _11371_/A _11347_/B _11414_/A vssd1 vssd1 vccd1 vccd1 _11299_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_26_1022 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13038_ _10734_/X _14893_/Q _13038_/S vssd1 vssd1 vccd1 vccd1 _13038_/X sky130_fd_sc_hd__mux2_2
XFILLER_140_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_1055 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14989_ _15021_/CLK _14989_/D vssd1 vssd1 vccd1 vccd1 _14989_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07530_ _14760_/Q _13439_/Q _07535_/S vssd1 vssd1 vccd1 vccd1 _13439_/D sky130_fd_sc_hd__mux2_1
XFILLER_47_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07461_ _13340_/A0 _13404_/Q _07501_/S vssd1 vssd1 vccd1 vccd1 _13404_/D sky130_fd_sc_hd__mux2_1
XFILLER_179_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_182_clk clkbuf_5_20_0_clk/X vssd1 vssd1 vccd1 vccd1 _15677_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_50_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09200_ _14371_/Q _15187_/Q _13826_/Q _14565_/Q _09438_/S0 _09448_/S1 vssd1 vssd1
+ vccd1 vccd1 _09201_/B sky130_fd_sc_hd__mux4_1
XFILLER_34_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07392_ _14738_/Q _07391_/X _07500_/S vssd1 vssd1 vccd1 vccd1 _07392_/X sky130_fd_sc_hd__mux2_8
XFILLER_188_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09131_ _14529_/Q _14142_/Q _14174_/Q _14110_/Q _09225_/S0 _09225_/S1 vssd1 vssd1
+ vccd1 vccd1 _09131_/X sky130_fd_sc_hd__mux4_1
XFILLER_175_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09062_ _09405_/A _09062_/B _09062_/C vssd1 vssd1 vccd1 vccd1 _09062_/X sky130_fd_sc_hd__and3_1
XFILLER_163_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08013_ _13570_/Q _13569_/Q _08017_/D vssd1 vssd1 vccd1 vccd1 _08018_/B sky130_fd_sc_hd__and3_1
XFILLER_135_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09964_ _11710_/A _09964_/B vssd1 vssd1 vccd1 vccd1 _09964_/Y sky130_fd_sc_hd__nand2b_4
XFILLER_44_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08915_ _13876_/Q _13123_/B _08508_/Y _14391_/Q _13123_/A vssd1 vssd1 vccd1 vccd1
+ _08915_/X sky130_fd_sc_hd__a221o_1
XFILLER_58_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09895_ _13110_/B2 _14257_/Q _09897_/S vssd1 vssd1 vccd1 vccd1 _14257_/D sky130_fd_sc_hd__mux2_1
XFILLER_58_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08846_ _13869_/Q _13345_/A0 _08846_/S vssd1 vssd1 vccd1 vccd1 _13869_/D sky130_fd_sc_hd__mux2_1
XTAP_3506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08777_ _08777_/A _08777_/B vssd1 vssd1 vccd1 vccd1 _08779_/B sky130_fd_sc_hd__nand2_1
XTAP_2805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07728_ _07750_/A _07728_/B vssd1 vssd1 vccd1 vccd1 _07728_/Y sky130_fd_sc_hd__nand2_1
XTAP_2838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_173_clk clkbuf_5_23_0_clk/X vssd1 vssd1 vccd1 vccd1 _15304_/CLK sky130_fd_sc_hd__clkbuf_16
X_07659_ _14722_/Q _14721_/Q _14723_/Q _10098_/B vssd1 vssd1 vccd1 vccd1 _07907_/A
+ sky130_fd_sc_hd__nor4_4
XFILLER_129_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10670_ _14752_/Q _10669_/X _10715_/S vssd1 vssd1 vccd1 vccd1 _14752_/D sky130_fd_sc_hd__mux2_1
XFILLER_185_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09329_ _14249_/Q _14281_/Q _14313_/Q _14345_/Q _09469_/S _09546_/S1 vssd1 vssd1
+ vccd1 vccd1 _09329_/X sky130_fd_sc_hd__mux4_1
XFILLER_178_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_89 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12340_ _12333_/X _12335_/X _12337_/X _12339_/X _12616_/C1 vssd1 vssd1 vccd1 vccd1
+ _12340_/X sky130_fd_sc_hd__o221a_1
XFILLER_21_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_412 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12271_ _12264_/X _12266_/X _12268_/X _12270_/X _12455_/C1 vssd1 vssd1 vccd1 vccd1
+ _12271_/X sky130_fd_sc_hd__o221a_1
XFILLER_107_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14010_ _15276_/CLK _14010_/D vssd1 vssd1 vccd1 vccd1 _14010_/Q sky130_fd_sc_hd__dfxtp_1
X_11222_ _10528_/B _15010_/Q _11232_/S vssd1 vssd1 vccd1 vccd1 _15010_/D sky130_fd_sc_hd__mux2_1
XFILLER_153_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11153_ _11344_/A _11152_/X _11151_/Y _11202_/A vssd1 vssd1 vccd1 vccd1 _11153_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_108_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10104_ _14490_/Q _14738_/Q _10131_/S vssd1 vssd1 vccd1 vccd1 _14490_/D sky130_fd_sc_hd__mux2_1
XFILLER_95_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11084_ _11020_/Y _11038_/Y _11318_/S vssd1 vssd1 vccd1 vccd1 _11084_/X sky130_fd_sc_hd__mux2_1
XFILLER_150_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10035_ _14392_/Q _11854_/A1 _10064_/S vssd1 vssd1 vccd1 vccd1 _14392_/D sky130_fd_sc_hd__mux2_1
X_14912_ _15542_/CLK _14912_/D vssd1 vssd1 vccd1 vccd1 _14912_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14843_ _15587_/CLK _14843_/D vssd1 vssd1 vccd1 vccd1 _14843_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_84_52 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14774_ _14774_/CLK _14774_/D vssd1 vssd1 vccd1 vccd1 _14774_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_112_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11986_ _12273_/A1 _11981_/X _11984_/X _11985_/X _08449_/A vssd1 vssd1 vccd1 vccd1
+ _11998_/B sky130_fd_sc_hd__a221o_1
XFILLER_1_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13725_ _15006_/CLK _13725_/D vssd1 vssd1 vccd1 vccd1 _13725_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10937_ _11589_/B _10951_/B vssd1 vssd1 vccd1 vccd1 _10937_/Y sky130_fd_sc_hd__nand2_1
XFILLER_56_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_164_clk clkbuf_5_22_0_clk/X vssd1 vssd1 vccd1 vccd1 _15077_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_108_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13656_ _14851_/CLK _13656_/D vssd1 vssd1 vccd1 vccd1 _13656_/Q sky130_fd_sc_hd__dfxtp_1
X_10868_ _14900_/Q _15528_/Q _10868_/S vssd1 vssd1 vccd1 vccd1 _14900_/D sky130_fd_sc_hd__mux2_1
XFILLER_9_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12607_ _12618_/A1 _12602_/X _12605_/X _12606_/X _08405_/D vssd1 vssd1 vccd1 vccd1
+ _12619_/B sky130_fd_sc_hd__a221o_1
XPHY_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13587_ _15647_/CLK _13587_/D vssd1 vssd1 vccd1 vccd1 _13587_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10799_ _14831_/Q _07327_/A _10868_/S vssd1 vssd1 vccd1 vccd1 _14831_/D sky130_fd_sc_hd__mux2_1
X_15326_ _15326_/CLK _15326_/D vssd1 vssd1 vccd1 vccd1 _15326_/Q sky130_fd_sc_hd__dfxtp_4
X_12538_ _12595_/A1 _12533_/X _12536_/X _12537_/X _08405_/D vssd1 vssd1 vccd1 vccd1
+ _12550_/B sky130_fd_sc_hd__a221o_1
XFILLER_158_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15257_ _15289_/CLK _15257_/D vssd1 vssd1 vccd1 vccd1 _15257_/Q sky130_fd_sc_hd__dfxtp_1
X_12469_ _12503_/A1 _12464_/X _12467_/X _12468_/X _12515_/C1 vssd1 vssd1 vccd1 vccd1
+ _12481_/B sky130_fd_sc_hd__a221o_1
XFILLER_67_1100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14208_ _14530_/CLK _14208_/D vssd1 vssd1 vccd1 vccd1 _14208_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_126_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_172_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15188_ _15289_/CLK _15188_/D vssd1 vssd1 vccd1 vccd1 _15188_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_153_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_523 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14139_ _15657_/CLK _14139_/D vssd1 vssd1 vccd1 vccd1 _14139_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout409 _11354_/X vssd1 vssd1 vccd1 vccd1 _11641_/S sky130_fd_sc_hd__buf_12
XFILLER_101_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06961_ _14490_/Q _06746_/Y _14489_/Q _06748_/Y _06960_/Y vssd1 vssd1 vccd1 vccd1
+ _06961_/X sky130_fd_sc_hd__a221o_1
X_08700_ _13619_/Q _08750_/B1 _08538_/Y _15375_/Q _08697_/X vssd1 vssd1 vccd1 vccd1
+ _08700_/X sky130_fd_sc_hd__a221o_1
XFILLER_79_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09680_ _14051_/Q _13335_/A0 _09690_/S vssd1 vssd1 vccd1 vccd1 _14051_/D sky130_fd_sc_hd__mux2_1
XFILLER_67_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06892_ _15399_/Q _06688_/Y _06883_/X _06891_/X vssd1 vssd1 vccd1 vccd1 _06892_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_94_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08631_ _14503_/Q _08693_/A2 _08629_/X _08630_/X vssd1 vssd1 vccd1 vccd1 _08632_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_39_378 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08562_ _13472_/Q _08746_/A2 _08750_/A2 _13536_/Q _08561_/X vssd1 vssd1 vccd1 vccd1
+ _08566_/B sky130_fd_sc_hd__a221o_1
XFILLER_74_1104 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07513_ _14743_/Q _13422_/Q _07529_/S vssd1 vssd1 vccd1 vccd1 _13422_/D sky130_fd_sc_hd__mux2_1
XFILLER_23_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08493_ _09532_/A _09524_/A vssd1 vssd1 vccd1 vccd1 _08497_/A sky130_fd_sc_hd__nor2_8
XFILLER_63_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_155_clk clkbuf_5_18_0_clk/X vssd1 vssd1 vccd1 vccd1 _15525_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_161_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07444_ _14751_/Q _07443_/X _07480_/S vssd1 vssd1 vccd1 vccd1 _07444_/X sky130_fd_sc_hd__mux2_8
XFILLER_50_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07375_ _13649_/Q _07499_/A2 _07499_/B1 _14677_/Q _07371_/X vssd1 vssd1 vccd1 vccd1
+ _07375_/X sky130_fd_sc_hd__a221o_1
XFILLER_149_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09114_ _09405_/A _09107_/X _09110_/X _09450_/B1 vssd1 vssd1 vccd1 vccd1 _09114_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_129_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09045_ _14074_/Q _09445_/A2 _09522_/B1 _14042_/Q _09391_/A vssd1 vssd1 vccd1 vccd1
+ _09045_/X sky130_fd_sc_hd__a221o_1
XFILLER_159_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_887 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09947_ _13334_/A0 _14307_/Q _09958_/S vssd1 vssd1 vccd1 vccd1 _14307_/D sky130_fd_sc_hd__mux2_1
XFILLER_104_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09878_ _13331_/A0 _14240_/Q _09892_/S vssd1 vssd1 vccd1 vccd1 _14240_/D sky130_fd_sc_hd__mux2_1
XTAP_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08829_ _13852_/Q _11861_/A1 _08846_/S vssd1 vssd1 vccd1 vccd1 _13852_/D sky130_fd_sc_hd__mux2_1
XFILLER_73_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11840_ _15262_/Q _11873_/A1 _11850_/S vssd1 vssd1 vccd1 vccd1 _15262_/D sky130_fd_sc_hd__mux2_1
XTAP_2624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11771_ _11879_/A1 _15199_/Q _11775_/S vssd1 vssd1 vccd1 vccd1 _15199_/D sky130_fd_sc_hd__mux2_1
XTAP_2679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_146_clk clkbuf_5_25_0_clk/X vssd1 vssd1 vccd1 vccd1 _15461_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_26_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13510_ _15372_/CLK _13510_/D vssd1 vssd1 vccd1 vccd1 _13510_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10722_ _15582_/Q _10706_/B _10722_/B1 _14959_/Q vssd1 vssd1 vccd1 vccd1 _10722_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_159_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14490_ _15399_/CLK _14490_/D vssd1 vssd1 vccd1 vccd1 _14490_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_1989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13441_ _14493_/CLK _13441_/D vssd1 vssd1 vccd1 vccd1 _13441_/Q sky130_fd_sc_hd__dfxtp_1
X_10653_ _15568_/Q _10731_/B _10718_/A2 _14977_/Q vssd1 vssd1 vccd1 vccd1 _10653_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_110_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13372_ _14475_/Q vssd1 vssd1 vccd1 vccd1 _14475_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_6_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10584_ _07104_/C _10734_/A2 _10580_/X _10583_/X vssd1 vssd1 vccd1 vccd1 _10584_/X
+ sky130_fd_sc_hd__o22a_4
XFILLER_166_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_103 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15111_ _15303_/CLK _15111_/D vssd1 vssd1 vccd1 vccd1 _15111_/Q sky130_fd_sc_hd__dfxtp_1
X_12323_ _14473_/Q _14441_/Q _13862_/Q _14215_/Q _12543_/S _12544_/A vssd1 vssd1 vccd1
+ vccd1 _12323_/X sky130_fd_sc_hd__mux4_1
XFILLER_127_659 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_979 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15042_ _15042_/CLK _15042_/D vssd1 vssd1 vccd1 vccd1 _15042_/Q sky130_fd_sc_hd__dfxtp_1
X_12254_ _14470_/Q _14438_/Q _13859_/Q _14212_/Q _11993_/S _11992_/A vssd1 vssd1 vccd1
+ vccd1 _12254_/X sky130_fd_sc_hd__mux4_1
XFILLER_107_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11205_ _10555_/C _14994_/Q _11237_/S vssd1 vssd1 vccd1 vccd1 _14994_/D sky130_fd_sc_hd__mux2_1
XFILLER_135_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12185_ _14467_/Q _14435_/Q _13856_/Q _14209_/Q _12489_/S0 _12489_/S1 vssd1 vssd1
+ vccd1 vccd1 _12185_/X sky130_fd_sc_hd__mux4_1
XFILLER_69_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11136_ _11347_/A _11136_/B vssd1 vssd1 vccd1 vccd1 _11136_/X sky130_fd_sc_hd__or2_1
XFILLER_49_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11067_ _11065_/X _11066_/X _11252_/A vssd1 vssd1 vccd1 vccd1 _11067_/X sky130_fd_sc_hd__mux2_2
XFILLER_95_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_985 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10018_ _13339_/A0 _14376_/Q _10029_/S vssd1 vssd1 vccd1 vccd1 _14376_/D sky130_fd_sc_hd__mux2_1
XFILLER_92_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14826_ _15644_/CLK _14826_/D vssd1 vssd1 vccd1 vccd1 _14826_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14757_ _15438_/CLK _14757_/D vssd1 vssd1 vccd1 vccd1 _14757_/Q sky130_fd_sc_hd__dfxtp_4
X_11969_ _12080_/A _11969_/B vssd1 vssd1 vccd1 vccd1 _11969_/X sky130_fd_sc_hd__and2_1
XFILLER_63_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_137_clk clkbuf_5_29_0_clk/X vssd1 vssd1 vccd1 vccd1 _14517_/CLK sky130_fd_sc_hd__clkbuf_16
X_13708_ _15334_/CLK _13708_/D vssd1 vssd1 vccd1 vccd1 _13708_/Q sky130_fd_sc_hd__dfxtp_1
X_14688_ _14703_/CLK _14688_/D vssd1 vssd1 vccd1 vccd1 _14688_/Q sky130_fd_sc_hd__dfxtp_1
X_13639_ _15375_/CLK _13639_/D vssd1 vssd1 vccd1 vccd1 _13639_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07160_ _14860_/Q _14852_/Q _14844_/Q _14836_/Q _08094_/S _07104_/C vssd1 vssd1 vccd1
+ vccd1 _07161_/B sky130_fd_sc_hd__mux4_1
XFILLER_118_615 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_271 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15309_ _15510_/CLK _15309_/D vssd1 vssd1 vccd1 vccd1 _15309_/Q sky130_fd_sc_hd__dfxtp_1
X_07091_ _07090_/X _13609_/Q _12662_/S vssd1 vssd1 vccd1 vccd1 _07091_/X sky130_fd_sc_hd__mux2_1
XFILLER_146_968 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout206 _09696_/X vssd1 vssd1 vccd1 vccd1 _09728_/S sky130_fd_sc_hd__buf_12
XFILLER_119_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09801_ _14167_/Q _13323_/A0 _09823_/S vssd1 vssd1 vccd1 vccd1 _14167_/D sky130_fd_sc_hd__mux2_1
Xfanout217 _08819_/Y vssd1 vssd1 vccd1 vccd1 _08846_/S sky130_fd_sc_hd__buf_12
XFILLER_141_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout228 _07736_/A vssd1 vssd1 vccd1 vccd1 _07676_/A sky130_fd_sc_hd__buf_6
X_07993_ _07971_/A _07992_/X input35/X vssd1 vssd1 vccd1 vccd1 _07993_/Y sky130_fd_sc_hd__a21oi_1
Xfanout239 _13024_/B2 vssd1 vssd1 vccd1 vccd1 _12944_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_140_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09732_ _14100_/Q _13320_/A0 _09762_/S vssd1 vssd1 vccd1 vccd1 _14100_/D sky130_fd_sc_hd__mux2_1
XFILLER_86_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06944_ _06944_/A _06944_/B _06944_/C _06944_/D vssd1 vssd1 vccd1 vccd1 _06945_/A
+ sky130_fd_sc_hd__nor4_4
XFILLER_101_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09663_ _09696_/B _11818_/A vssd1 vssd1 vccd1 vccd1 _09663_/Y sky130_fd_sc_hd__nor2_8
XFILLER_27_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06875_ _06697_/Y _13504_/Q _06882_/B _06871_/Y _06873_/Y vssd1 vssd1 vccd1 vccd1
+ _06875_/X sky130_fd_sc_hd__o221a_1
XFILLER_27_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08614_ _13528_/Q _08683_/A2 _08691_/A2 _13599_/Q vssd1 vssd1 vccd1 vccd1 _08614_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_82_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09594_ _13970_/Q _13350_/A0 _09594_/S vssd1 vssd1 vccd1 vccd1 _13970_/D sky130_fd_sc_hd__mux2_1
XTAP_1208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08545_ _13571_/Q _08747_/A2 _08544_/X _08722_/A vssd1 vssd1 vccd1 vccd1 _08545_/X
+ sky130_fd_sc_hd__a211o_1
Xclkbuf_leaf_128_clk clkbuf_5_31_0_clk/X vssd1 vssd1 vccd1 vccd1 _14511_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_36_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08476_ _13769_/Q _13120_/S _08470_/X _14608_/Q vssd1 vssd1 vccd1 vccd1 _13769_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_126_1024 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_1098 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07427_ _13662_/Q _07483_/A2 _07483_/B1 _14690_/Q _07426_/X vssd1 vssd1 vccd1 vccd1
+ _07427_/X sky130_fd_sc_hd__a221o_1
XFILLER_50_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07358_ _07230_/C _07357_/X _07227_/Y vssd1 vssd1 vccd1 vccd1 _07358_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_109_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_570 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07289_ _07339_/S _13919_/Q _07288_/Y vssd1 vssd1 vccd1 vccd1 _07289_/X sky130_fd_sc_hd__o21a_4
X_09028_ _13945_/Q _13687_/Q _09521_/S vssd1 vssd1 vccd1 vccd1 _09028_/X sky130_fd_sc_hd__mux2_1
XFILLER_123_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_1039 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13990_ _15127_/CLK _13990_/D vssd1 vssd1 vccd1 vccd1 _13990_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12941_ _08405_/D _13318_/C _08817_/Y _06670_/A _12940_/X vssd1 vssd1 vccd1 vccd1
+ _12941_/Y sky130_fd_sc_hd__o221ai_2
XTAP_3111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15660_ _15660_/CLK _15660_/D vssd1 vssd1 vccd1 vccd1 _15660_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12872_ _15400_/Q _15585_/Q _12904_/S vssd1 vssd1 vccd1 vccd1 _15400_/D sky130_fd_sc_hd__mux2_1
XTAP_2410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_100 _15050_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_111 input8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_122 _07105_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14611_ _15648_/CLK _14611_/D vssd1 vssd1 vccd1 vccd1 _14611_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_2443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11823_ _15245_/Q _13323_/A0 _11849_/S vssd1 vssd1 vccd1 vccd1 _15245_/D sky130_fd_sc_hd__mux2_1
XANTENNA_133 input24/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_119_clk clkbuf_5_30_0_clk/X vssd1 vssd1 vccd1 vccd1 _14495_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_3199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15591_ _15591_/CLK _15591_/D vssd1 vssd1 vccd1 vccd1 _15591_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_802 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14542_ _14542_/CLK _14542_/D vssd1 vssd1 vccd1 vccd1 _14542_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11754_ _13329_/A0 _15182_/Q _11774_/S vssd1 vssd1 vccd1 vccd1 _15182_/D sky130_fd_sc_hd__mux2_1
XFILLER_186_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_576 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10705_ _14759_/Q _10704_/X _10710_/S vssd1 vssd1 vccd1 vccd1 _14759_/D sky130_fd_sc_hd__mux2_1
XTAP_1797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14473_ _14537_/CLK _14473_/D vssd1 vssd1 vccd1 vccd1 _14473_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11685_ _13327_/A0 _15116_/Q _11703_/S vssd1 vssd1 vccd1 vccd1 _15116_/D sky130_fd_sc_hd__mux2_1
XFILLER_81_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13424_ _15379_/CLK _13424_/D vssd1 vssd1 vccd1 vccd1 _13424_/Q sky130_fd_sc_hd__dfxtp_4
X_10636_ _15565_/Q _10706_/B vssd1 vssd1 vccd1 vccd1 _10636_/X sky130_fd_sc_hd__and2_1
XFILLER_155_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_220 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13355_ _14458_/Q vssd1 vssd1 vccd1 vccd1 _14458_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_6_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10567_ _14928_/Q _14927_/Q vssd1 vssd1 vccd1 vccd1 _10567_/Y sky130_fd_sc_hd__nor2_2
XFILLER_182_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12306_ _12536_/A _12306_/B vssd1 vssd1 vccd1 vccd1 _12306_/X sky130_fd_sc_hd__or2_1
X_13286_ _06658_/Y _15618_/Q _13291_/S vssd1 vssd1 vccd1 vccd1 _15618_/D sky130_fd_sc_hd__mux2_1
X_10498_ _07242_/X _08225_/Y _10497_/X vssd1 vssd1 vccd1 vccd1 _11569_/B sky130_fd_sc_hd__a21oi_4
XFILLER_6_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15025_ _15581_/CLK _15025_/D vssd1 vssd1 vccd1 vccd1 _15025_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12237_ _12502_/S _12237_/B vssd1 vssd1 vccd1 vccd1 _12237_/X sky130_fd_sc_hd__or2_1
XFILLER_107_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12168_ _12168_/A _12168_/B vssd1 vssd1 vccd1 vccd1 _12168_/X sky130_fd_sc_hd__or2_1
XFILLER_2_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11119_ _14968_/Q _10984_/Y _11118_/X vssd1 vssd1 vccd1 vccd1 _14968_/D sky130_fd_sc_hd__a21o_1
XFILLER_110_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12099_ _12260_/A _12099_/B vssd1 vssd1 vccd1 vccd1 _12099_/X sky130_fd_sc_hd__or2_1
XFILLER_7_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput6 ext_read_data[14] vssd1 vssd1 vccd1 vccd1 input6/X sky130_fd_sc_hd__clkbuf_4
XFILLER_77_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06660_ _07096_/S vssd1 vssd1 vccd1 vccd1 _07787_/A sky130_fd_sc_hd__inv_2
XFILLER_24_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_178 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14809_ _15628_/CLK _14809_/D vssd1 vssd1 vccd1 vccd1 _14809_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08330_ _08289_/X _08329_/X _11047_/B vssd1 vssd1 vccd1 vccd1 _08330_/X sky130_fd_sc_hd__mux2_2
XFILLER_33_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08261_ _11356_/B _10551_/A vssd1 vssd1 vccd1 vccd1 _08261_/X sky130_fd_sc_hd__and2_2
X_07212_ _07206_/X _07208_/Y _07210_/Y _07211_/X vssd1 vssd1 vccd1 vccd1 _07356_/A
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_137_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08192_ _13683_/Q _11854_/A1 _08221_/S vssd1 vssd1 vccd1 vccd1 _13683_/D sky130_fd_sc_hd__mux2_1
XFILLER_119_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07143_ _14835_/Q _07104_/X _07142_/X _07131_/A vssd1 vssd1 vccd1 vccd1 _07143_/X
+ sky130_fd_sc_hd__a22o_4
XFILLER_146_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07074_ _07073_/X _14757_/Q _07077_/S vssd1 vssd1 vccd1 vccd1 _13603_/D sky130_fd_sc_hd__mux2_1
XFILLER_146_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07976_ _14752_/Q _07971_/A _07975_/Y _07987_/C1 vssd1 vssd1 vccd1 vccd1 _13559_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_142_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09715_ _13337_/A0 _14085_/Q _09728_/S vssd1 vssd1 vccd1 vccd1 _14085_/D sky130_fd_sc_hd__mux2_1
X_06927_ _15395_/Q _06699_/Y _15394_/Q _06701_/Y _06888_/A vssd1 vssd1 vccd1 vccd1
+ _06927_/X sky130_fd_sc_hd__o221a_1
XFILLER_56_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09646_ _14019_/Q _13335_/A0 _09660_/S vssd1 vssd1 vccd1 vccd1 _14019_/D sky130_fd_sc_hd__mux2_1
X_06858_ _12834_/B vssd1 vssd1 vccd1 vccd1 _12828_/A sky130_fd_sc_hd__inv_4
XFILLER_35_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09577_ _13953_/Q _13333_/A0 _09589_/S vssd1 vssd1 vccd1 vccd1 _13953_/D sky130_fd_sc_hd__mux2_1
XFILLER_35_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06789_ _14587_/Q _06789_/B vssd1 vssd1 vccd1 vccd1 _08465_/B sky130_fd_sc_hd__nor2_8
XTAP_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08528_ _14609_/Q _08536_/B _08528_/C vssd1 vssd1 vccd1 vccd1 _08531_/C sky130_fd_sc_hd__or3_4
XFILLER_11_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08459_ _14597_/Q _08773_/B vssd1 vssd1 vccd1 vccd1 _08459_/X sky130_fd_sc_hd__and2_1
X_11470_ _13195_/B _11470_/B vssd1 vssd1 vccd1 vccd1 _11471_/B sky130_fd_sc_hd__and2_1
XFILLER_183_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10421_ _10507_/A1 _13744_/Q _15428_/Q _10515_/B2 vssd1 vssd1 vccd1 vccd1 _10421_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_136_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13140_ _08754_/A hold3/A _13140_/S vssd1 vssd1 vccd1 vccd1 _15537_/D sky130_fd_sc_hd__mux2_1
X_10352_ _10520_/A1 _13792_/Q _13760_/Q _10520_/B2 vssd1 vssd1 vccd1 vccd1 _10352_/X
+ sky130_fd_sc_hd__a22o_2
XFILLER_151_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13071_ _15503_/Q _13081_/A2 _13105_/B1 _13070_/X vssd1 vssd1 vccd1 vccd1 _15503_/D
+ sky130_fd_sc_hd__a22o_1
X_10283_ _14668_/Q _14821_/Q _10630_/S vssd1 vssd1 vccd1 vccd1 _14668_/D sky130_fd_sc_hd__mux2_1
XFILLER_183_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12022_ _15311_/Q _10877_/S _12021_/X vssd1 vssd1 vccd1 vccd1 _15311_/D sky130_fd_sc_hd__a21o_1
XFILLER_105_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout570 _08451_/A vssd1 vssd1 vccd1 vccd1 _12501_/C1 sky130_fd_sc_hd__buf_12
Xfanout581 _14600_/Q vssd1 vssd1 vccd1 vccd1 _08405_/B sky130_fd_sc_hd__buf_12
Xfanout592 fanout600/X vssd1 vssd1 vccd1 vccd1 _12590_/A sky130_fd_sc_hd__buf_12
XFILLER_111_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13973_ _15142_/CLK _13973_/D vssd1 vssd1 vccd1 vccd1 _13973_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_76_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12924_ _15452_/Q _15638_/Q _12929_/S vssd1 vssd1 vccd1 vccd1 _15452_/D sky130_fd_sc_hd__mux2_1
XFILLER_20_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12855_ _14749_/Q _15383_/Q _12866_/S vssd1 vssd1 vccd1 vccd1 _15383_/D sky130_fd_sc_hd__mux2_1
X_15643_ _15643_/CLK _15643_/D vssd1 vssd1 vccd1 vccd1 _15643_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_852 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11806_ _15229_/Q _11872_/A1 _11817_/S vssd1 vssd1 vccd1 vccd1 _15229_/D sky130_fd_sc_hd__mux2_1
X_15574_ _15581_/CLK _15574_/D vssd1 vssd1 vccd1 vccd1 _15574_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12786_ _15067_/Q _12783_/X _12792_/B vssd1 vssd1 vccd1 vccd1 _12786_/X sky130_fd_sc_hd__mux2_1
XTAP_1550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_632 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14525_ _14525_/CLK _14525_/D vssd1 vssd1 vccd1 vccd1 _14525_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11737_ _15166_/Q _13104_/B2 _11741_/S vssd1 vssd1 vccd1 vccd1 _15166_/D sky130_fd_sc_hd__mux2_1
XFILLER_175_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14456_ _15668_/CLK _14456_/D vssd1 vssd1 vccd1 vccd1 _14456_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_175_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11668_ _13343_/A0 _15100_/Q _11670_/S vssd1 vssd1 vccd1 vccd1 _15100_/D sky130_fd_sc_hd__mux2_1
XFILLER_128_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_1028 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13407_ _15500_/CLK _13407_/D vssd1 vssd1 vccd1 vccd1 _13407_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10619_ _15051_/Q _10714_/A2 _10616_/X _10618_/X vssd1 vssd1 vccd1 vccd1 _10619_/X
+ sky130_fd_sc_hd__o22a_2
X_14387_ _15203_/CLK _14387_/D vssd1 vssd1 vccd1 vccd1 _14387_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11599_ _13236_/A _11599_/B vssd1 vssd1 vccd1 vccd1 _11600_/B sky130_fd_sc_hd__or2_1
XFILLER_128_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_404 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13338_ _13338_/A0 _15668_/Q _13350_/S vssd1 vssd1 vccd1 vccd1 _15668_/D sky130_fd_sc_hd__mux2_1
Xclkbuf_5_18_0_clk clkbuf_4_9_0_clk/X vssd1 vssd1 vccd1 vccd1 clkbuf_5_18_0_clk/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_115_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13269_ _15353_/Q _15600_/Q _13309_/A vssd1 vssd1 vccd1 vccd1 _15600_/D sky130_fd_sc_hd__mux2_1
XFILLER_44_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_1080 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15008_ _15020_/CLK _15008_/D vssd1 vssd1 vccd1 vccd1 _15008_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_97_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07830_ _07830_/A _07830_/B vssd1 vssd1 vccd1 vccd1 _07830_/Y sky130_fd_sc_hd__nand2_1
XFILLER_96_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_1067 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07761_ _13504_/Q _07765_/C vssd1 vssd1 vccd1 vccd1 _07764_/B sky130_fd_sc_hd__and2_1
XFILLER_2_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09500_ _13872_/Q _14225_/Q _09535_/S vssd1 vssd1 vccd1 vccd1 _09500_/X sky130_fd_sc_hd__mux2_1
XFILLER_110_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06712_ _15388_/Q vssd1 vssd1 vccd1 vccd1 _06712_/Y sky130_fd_sc_hd__inv_2
XFILLER_65_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07692_ _14742_/Q _07713_/A _07691_/Y _07949_/C1 vssd1 vssd1 vccd1 vccd1 _13485_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_64_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09431_ _09405_/A _09424_/X _09427_/X _09450_/B1 vssd1 vssd1 vccd1 vccd1 _09431_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_53_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09362_ _09523_/A1 _09360_/X _09361_/X vssd1 vssd1 vccd1 vccd1 _09362_/X sky130_fd_sc_hd__a21o_1
XFILLER_80_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08313_ _11419_/A vssd1 vssd1 vccd1 vccd1 _08313_/Y sky130_fd_sc_hd__inv_2
XFILLER_33_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09293_ _14086_/Q _09522_/A2 _08512_/B _14054_/Q _09532_/A vssd1 vssd1 vccd1 vccd1
+ _09293_/X sky130_fd_sc_hd__a221o_1
XFILLER_75_1095 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_11 _10634_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_22 _13784_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_33 _14754_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08244_ _08244_/A _08244_/B vssd1 vssd1 vccd1 vccd1 _08244_/Y sky130_fd_sc_hd__nor2_2
XFILLER_178_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_44 input21/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_55 _07193_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_66 _07129_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_77 _07159_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08175_ _08133_/S input19/X _08185_/A vssd1 vssd1 vccd1 vccd1 _08175_/X sky130_fd_sc_hd__and3b_1
XANTENNA_88 _12515_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_99 _15065_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07126_ _14843_/Q _14835_/Q _08150_/S vssd1 vssd1 vccd1 vccd1 _07127_/B sky130_fd_sc_hd__mux2_1
XFILLER_118_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07057_ _14631_/Q _14663_/Q _07078_/S vssd1 vssd1 vccd1 vccd1 _07057_/X sky130_fd_sc_hd__mux2_1
XFILLER_134_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07959_ _07964_/A _07959_/B vssd1 vssd1 vccd1 vccd1 _07959_/Y sky130_fd_sc_hd__nand2_1
XFILLER_28_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10970_ _11025_/A _11500_/A vssd1 vssd1 vccd1 vccd1 _11242_/A sky130_fd_sc_hd__and2_1
XFILLER_28_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09629_ _13318_/D _09696_/B vssd1 vssd1 vccd1 vccd1 _09629_/Y sky130_fd_sc_hd__nor2_8
XFILLER_43_435 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12640_ _13417_/Q _12639_/X _12640_/S vssd1 vssd1 vccd1 vccd1 _12641_/B sky130_fd_sc_hd__mux2_1
XFILLER_62_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12571_ _12554_/X _12555_/X _12594_/S vssd1 vssd1 vccd1 vccd1 _12571_/X sky130_fd_sc_hd__mux2_1
XFILLER_62_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_50_clk clkbuf_5_8_0_clk/X vssd1 vssd1 vccd1 vccd1 _14997_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_11_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14310_ _15301_/CLK _14310_/D vssd1 vssd1 vccd1 vccd1 _14310_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_184_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11522_ _11531_/A _11522_/B vssd1 vssd1 vccd1 vccd1 _11544_/A sky130_fd_sc_hd__nand2_1
XFILLER_184_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15290_ _15666_/CLK _15290_/D vssd1 vssd1 vccd1 vccd1 _15290_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14241_ _15267_/CLK _14241_/D vssd1 vssd1 vccd1 vccd1 _14241_/Q sky130_fd_sc_hd__dfxtp_1
X_11453_ _11452_/Y _15054_/Q _11474_/S vssd1 vssd1 vccd1 vccd1 _15054_/D sky130_fd_sc_hd__mux2_1
XFILLER_165_860 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10404_ _11362_/B _13162_/B _10403_/Y _08261_/X vssd1 vssd1 vccd1 vccd1 _10404_/X
+ sky130_fd_sc_hd__a211o_1
X_14172_ _15663_/CLK _14172_/D vssd1 vssd1 vccd1 vccd1 _14172_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_164_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11384_ _11384_/A _11384_/B vssd1 vssd1 vccd1 vccd1 _11401_/A sky130_fd_sc_hd__nor2_1
XFILLER_180_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13123_ _13123_/A _13123_/B vssd1 vssd1 vccd1 vccd1 _13123_/Y sky130_fd_sc_hd__nor2_1
X_10335_ _14720_/Q _14913_/Q _10343_/S vssd1 vssd1 vccd1 vccd1 _14720_/D sky130_fd_sc_hd__mux2_1
XFILLER_97_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13054_ _12948_/X _13118_/A2 _13114_/B1 _07380_/X vssd1 vssd1 vccd1 vccd1 _13054_/X
+ sky130_fd_sc_hd__a22o_1
X_10266_ _14651_/Q _14804_/Q _10610_/S vssd1 vssd1 vccd1 vccd1 _14651_/D sky130_fd_sc_hd__mux2_1
X_12005_ _14361_/Q _15177_/Q _13816_/Q _14555_/Q _12407_/S _12406_/A vssd1 vssd1 vccd1
+ vccd1 _12005_/X sky130_fd_sc_hd__mux4_1
XFILLER_79_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10197_ _13350_/A0 _14581_/Q _10197_/S vssd1 vssd1 vccd1 vccd1 _14581_/D sky130_fd_sc_hd__mux2_1
XFILLER_78_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13956_ _14373_/CLK _13956_/D vssd1 vssd1 vccd1 vccd1 _13956_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_46_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12907_ _15435_/Q _15621_/Q _12932_/S vssd1 vssd1 vccd1 vccd1 _15435_/D sky130_fd_sc_hd__mux2_1
X_13887_ _15233_/CLK _13887_/D vssd1 vssd1 vccd1 vccd1 _13887_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_185_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15626_ _15626_/CLK _15626_/D vssd1 vssd1 vccd1 vccd1 _15626_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12838_ _15367_/Q _12743_/A _12837_/X input35/X vssd1 vssd1 vccd1 vccd1 _15367_/D
+ sky130_fd_sc_hd__a211o_1
XTAP_2081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12769_ _12776_/B _12769_/B vssd1 vssd1 vccd1 vccd1 _12770_/B sky130_fd_sc_hd__nor2_1
XTAP_1380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15557_ _15558_/CLK _15557_/D vssd1 vssd1 vccd1 vccd1 _15557_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_41_clk clkbuf_5_9_0_clk/X vssd1 vssd1 vccd1 vccd1 _15613_/CLK sky130_fd_sc_hd__clkbuf_16
X_14508_ _14510_/CLK _14508_/D vssd1 vssd1 vccd1 vccd1 _14508_/Q sky130_fd_sc_hd__dfxtp_1
X_15488_ _15501_/CLK _15488_/D vssd1 vssd1 vccd1 vccd1 _15488_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_187_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_5_1_0_clk clkbuf_5_1_0_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_5_1_0_clk/X sky130_fd_sc_hd__clkbuf_8
XFILLER_159_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput20 ext_read_data[27] vssd1 vssd1 vccd1 vccd1 input20/X sky130_fd_sc_hd__buf_8
Xinput31 ext_read_data[8] vssd1 vssd1 vccd1 vccd1 input31/X sky130_fd_sc_hd__buf_8
X_14439_ _14439_/CLK _14439_/D vssd1 vssd1 vccd1 vccd1 _14439_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09980_ _13334_/A0 _14339_/Q _09991_/S vssd1 vssd1 vccd1 vccd1 _14339_/D sky130_fd_sc_hd__mux2_1
XFILLER_115_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08931_ _13123_/A _08930_/X _08929_/X _09554_/A vssd1 vssd1 vccd1 vccd1 _08931_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_130_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08862_ _13883_/Q _13327_/A0 _08880_/S vssd1 vssd1 vccd1 vccd1 _13883_/D sky130_fd_sc_hd__mux2_1
XFILLER_85_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07813_ _13517_/Q _13516_/Q _13515_/Q _07813_/D vssd1 vssd1 vccd1 vccd1 _07825_/D
+ sky130_fd_sc_hd__and4_4
XFILLER_57_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08793_ _11860_/A1 _13819_/Q _08811_/S vssd1 vssd1 vccd1 vccd1 _13819_/D sky130_fd_sc_hd__mux2_1
XFILLER_96_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07744_ _14756_/Q _07750_/A _07743_/Y _08002_/C1 vssd1 vssd1 vccd1 vccd1 _13499_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_26_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07675_ _13481_/Q _07679_/C vssd1 vssd1 vccd1 vccd1 _07676_/B sky130_fd_sc_hd__xnor2_1
XFILLER_25_435 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09414_ _09435_/A _09414_/B vssd1 vssd1 vccd1 vccd1 _09414_/X sky130_fd_sc_hd__or2_1
XFILLER_13_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09345_ _08510_/B _09341_/X _09344_/X _09340_/X vssd1 vssd1 vccd1 vccd1 _09346_/C
+ sky130_fd_sc_hd__a211o_1
Xclkbuf_leaf_32_clk clkbuf_5_7_0_clk/X vssd1 vssd1 vccd1 vccd1 _15529_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_139_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09276_ _14536_/Q _14149_/Q _14181_/Q _14117_/Q _09557_/S _09550_/A1 vssd1 vssd1
+ vccd1 vccd1 _09276_/X sky130_fd_sc_hd__mux4_1
XFILLER_148_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08227_ _07339_/X _10457_/A2 _08226_/X vssd1 vssd1 vccd1 vccd1 _08227_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_147_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08158_ _13666_/Q _10695_/S _08155_/X _08157_/X vssd1 vssd1 vccd1 vccd1 _13666_/D
+ sky130_fd_sc_hd__o22a_1
X_07109_ _14831_/Q _07115_/B _07163_/A vssd1 vssd1 vccd1 vccd1 _07109_/X sky130_fd_sc_hd__and3_4
X_08089_ _13648_/Q _08085_/S _08078_/B vssd1 vssd1 vccd1 vccd1 _08089_/Y sky130_fd_sc_hd__a21oi_1
X_10120_ _14506_/Q _14754_/Q _10124_/S vssd1 vssd1 vccd1 vccd1 _14506_/D sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_99_clk clkbuf_5_25_0_clk/X vssd1 vssd1 vccd1 vccd1 _15644_/CLK sky130_fd_sc_hd__clkbuf_16
X_10051_ _14408_/Q _13337_/A0 _10064_/S vssd1 vssd1 vccd1 vccd1 _14408_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13810_ _15208_/CLK _13810_/D vssd1 vssd1 vccd1 vccd1 _13810_/Q sky130_fd_sc_hd__dfxtp_1
X_14790_ _15422_/CLK _14790_/D vssd1 vssd1 vccd1 vccd1 _14790_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_169_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13741_ _15046_/CLK _13741_/D vssd1 vssd1 vccd1 vccd1 _14928_/D sky130_fd_sc_hd__dfxtp_4
XFILLER_113_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10953_ _11023_/A _13236_/B vssd1 vssd1 vccd1 vccd1 _11317_/A sky130_fd_sc_hd__and2_1
XFILLER_44_744 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13672_ _15612_/CLK _13672_/D vssd1 vssd1 vccd1 vccd1 _13672_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10884_ _14916_/Q _15547_/Q _13134_/A vssd1 vssd1 vccd1 vccd1 _14916_/D sky130_fd_sc_hd__mux2_1
XFILLER_73_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15411_ _15596_/CLK _15411_/D vssd1 vssd1 vccd1 vccd1 _15411_/Q sky130_fd_sc_hd__dfxtp_2
X_12623_ _15338_/Q _12834_/B vssd1 vssd1 vccd1 vccd1 _12623_/Y sky130_fd_sc_hd__nand2_1
XFILLER_31_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_23_clk clkbuf_5_3_0_clk/X vssd1 vssd1 vccd1 vccd1 _14093_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_145_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15342_ _15622_/CLK _15342_/D vssd1 vssd1 vccd1 vccd1 _15342_/Q sky130_fd_sc_hd__dfxtp_4
X_12554_ _14547_/Q _14160_/Q _14192_/Q _14128_/Q _12568_/S _12567_/A vssd1 vssd1 vccd1
+ vccd1 _12554_/X sky130_fd_sc_hd__mux4_1
XFILLER_129_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11505_ _11505_/A _11505_/B _11505_/C _11505_/D vssd1 vssd1 vccd1 vccd1 _11505_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_8_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15273_ _15273_/CLK _15273_/D vssd1 vssd1 vccd1 vccd1 _15273_/Q sky130_fd_sc_hd__dfxtp_1
X_12485_ _14544_/Q _14157_/Q _14189_/Q _14125_/Q _12499_/S _12486_/S1 vssd1 vssd1
+ vccd1 vccd1 _12485_/X sky130_fd_sc_hd__mux4_1
XFILLER_156_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_172_627 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14224_ _15200_/CLK _14224_/D vssd1 vssd1 vccd1 vccd1 _14224_/Q sky130_fd_sc_hd__dfxtp_1
X_11436_ _11436_/A _11436_/B vssd1 vssd1 vccd1 vccd1 _11437_/C sky130_fd_sc_hd__and2_1
XFILLER_153_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14155_ _15500_/CLK _14155_/D vssd1 vssd1 vccd1 vccd1 _14155_/Q sky130_fd_sc_hd__dfxtp_1
X_11367_ _11368_/A _11368_/B vssd1 vssd1 vccd1 vccd1 _11369_/B sky130_fd_sc_hd__nor2_1
XFILLER_152_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13106_ _13026_/X _13118_/A2 _13114_/B1 _07484_/X vssd1 vssd1 vccd1 vccd1 _13106_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_98_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10318_ _14703_/Q _14888_/Q _10710_/S vssd1 vssd1 vccd1 vccd1 _14703_/D sky130_fd_sc_hd__mux2_1
XTAP_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14086_ _14537_/CLK _14086_/D vssd1 vssd1 vccd1 vccd1 _14086_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11298_ _11298_/A _11298_/B vssd1 vssd1 vccd1 vccd1 _11298_/Y sky130_fd_sc_hd__nor2_1
XTAP_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13037_ _15492_/Q _13139_/S _13116_/C _13036_/X vssd1 vssd1 vccd1 vccd1 _15492_/D
+ sky130_fd_sc_hd__a22o_1
X_10249_ _14634_/Q _14787_/Q _10715_/S vssd1 vssd1 vccd1 vccd1 _14634_/D sky130_fd_sc_hd__mux2_1
XFILLER_26_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_1067 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14988_ _14988_/CLK _14988_/D vssd1 vssd1 vccd1 vccd1 _14988_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13939_ _15665_/CLK _13939_/D vssd1 vssd1 vccd1 vccd1 _13939_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07460_ _14755_/Q _07459_/X _07480_/S vssd1 vssd1 vccd1 vccd1 _07460_/X sky130_fd_sc_hd__mux2_8
XFILLER_23_939 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15609_ _15641_/CLK _15609_/D vssd1 vssd1 vccd1 vccd1 _15609_/Q sky130_fd_sc_hd__dfxtp_1
X_07391_ _13653_/Q _07499_/A2 _07499_/B1 _14681_/Q _07390_/X vssd1 vssd1 vccd1 vccd1
+ _07391_/X sky130_fd_sc_hd__a221o_1
Xclkbuf_leaf_14_clk clkbuf_5_2_0_clk/X vssd1 vssd1 vccd1 vccd1 _15298_/CLK sky130_fd_sc_hd__clkbuf_16
X_09130_ _09130_/A _09130_/B _09130_/C vssd1 vssd1 vccd1 vccd1 _09130_/X sky130_fd_sc_hd__and3_1
XFILLER_33_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09061_ _09234_/S1 _09059_/X _09060_/X vssd1 vssd1 vccd1 vccd1 _09062_/C sky130_fd_sc_hd__a21o_1
XFILLER_136_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08012_ _14762_/Q _08012_/A2 _08011_/Y _08012_/C1 vssd1 vssd1 vccd1 vccd1 _13569_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_131_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_896 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09963_ _13350_/A0 _14323_/Q _09963_/S vssd1 vssd1 vccd1 vccd1 _14323_/D sky130_fd_sc_hd__mux2_1
XFILLER_89_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08914_ _13940_/Q _13682_/Q _09469_/S vssd1 vssd1 vccd1 vccd1 _08914_/X sky130_fd_sc_hd__mux2_1
XTAP_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09894_ _11847_/A1 _14256_/Q _09897_/S vssd1 vssd1 vccd1 vccd1 _14256_/D sky130_fd_sc_hd__mux2_1
XFILLER_131_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08845_ _13868_/Q _11877_/A1 _08846_/S vssd1 vssd1 vccd1 vccd1 _13868_/D sky130_fd_sc_hd__mux2_1
XTAP_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08776_ _13807_/Q _10892_/B _08775_/X vssd1 vssd1 vccd1 vccd1 _13807_/D sky130_fd_sc_hd__a21o_1
XFILLER_57_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_327 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07727_ _13495_/Q _07727_/B vssd1 vssd1 vccd1 vccd1 _07728_/B sky130_fd_sc_hd__xnor2_1
XTAP_2828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07658_ _14724_/Q _07658_/B vssd1 vssd1 vccd1 vccd1 _10098_/B sky130_fd_sc_hd__nand2_2
XFILLER_168_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07589_ _07587_/Y _07603_/C _07607_/A vssd1 vssd1 vccd1 vccd1 _07589_/Y sky130_fd_sc_hd__o21ai_1
Xclkbuf_4_8_0_clk clkbuf_4_9_0_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_8_0_clk/X sky130_fd_sc_hd__clkbuf_8
XFILLER_13_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_235 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09328_ _13123_/A _09327_/X _09326_/X _09382_/A vssd1 vssd1 vccd1 vccd1 _09328_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_159_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09259_ _13924_/Q _09258_/X _12573_/A vssd1 vssd1 vccd1 vccd1 _13924_/D sky130_fd_sc_hd__mux2_1
XFILLER_154_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12270_ _12500_/A1 _12269_/X _12468_/A1 vssd1 vssd1 vccd1 vccd1 _12270_/X sky130_fd_sc_hd__a21o_1
XFILLER_111_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11221_ _10366_/C _15009_/Q _11232_/S vssd1 vssd1 vccd1 vccd1 _15009_/D sky130_fd_sc_hd__mux2_1
XFILLER_153_148 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11152_ _11093_/X _11098_/X _11283_/A vssd1 vssd1 vccd1 vccd1 _11152_/X sky130_fd_sc_hd__mux2_1
XFILLER_150_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10103_ _14489_/Q _14737_/Q _10131_/S vssd1 vssd1 vccd1 vccd1 _14489_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11083_ _11077_/X _11082_/Y _11347_/A vssd1 vssd1 vccd1 vccd1 _11177_/B sky130_fd_sc_hd__mux2_1
XFILLER_49_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10034_ _14391_/Q _11853_/A1 _10064_/S vssd1 vssd1 vccd1 vccd1 _14391_/D sky130_fd_sc_hd__mux2_1
X_14911_ _15542_/CLK _14911_/D vssd1 vssd1 vccd1 vccd1 _14911_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14842_ _15508_/CLK _14842_/D vssd1 vssd1 vccd1 vccd1 _14842_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11985_ _12500_/B1 _11982_/X _12501_/C1 vssd1 vssd1 vccd1 vccd1 _11985_/X sky130_fd_sc_hd__o21a_1
X_14773_ _15646_/CLK _14773_/D vssd1 vssd1 vccd1 vccd1 _14773_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13724_ _15006_/CLK _13724_/D vssd1 vssd1 vccd1 vccd1 _13724_/Q sky130_fd_sc_hd__dfxtp_1
X_10936_ _14952_/Q _10491_/A _10948_/B vssd1 vssd1 vccd1 vccd1 _14952_/D sky130_fd_sc_hd__mux2_1
XFILLER_95_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10867_ _14899_/Q _15536_/Q _13138_/S vssd1 vssd1 vccd1 vccd1 _14899_/D sky130_fd_sc_hd__mux2_1
X_13655_ _14892_/CLK _13655_/D vssd1 vssd1 vccd1 vccd1 _13655_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_158_911 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12606_ _12615_/B1 _12603_/X _12616_/C1 vssd1 vssd1 vccd1 vccd1 _12606_/X sky130_fd_sc_hd__o21a_1
X_13586_ _15622_/CLK _13586_/D vssd1 vssd1 vccd1 vccd1 _13586_/Q sky130_fd_sc_hd__dfxtp_2
XPHY_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10798_ _14830_/Q _07331_/A _12504_/A vssd1 vssd1 vccd1 vccd1 _14830_/D sky130_fd_sc_hd__mux2_1
XFILLER_185_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12537_ _12615_/B1 _12534_/X _12616_/C1 vssd1 vssd1 vccd1 vccd1 _12537_/X sky130_fd_sc_hd__o21a_1
X_15325_ _15676_/CLK _15325_/D vssd1 vssd1 vccd1 vccd1 _15325_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_487 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12468_ _12468_/A1 _12465_/X _12501_/C1 vssd1 vssd1 vccd1 vccd1 _12468_/X sky130_fd_sc_hd__o21a_1
X_15256_ _15332_/CLK _15256_/D vssd1 vssd1 vccd1 vccd1 _15256_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11419_ _11419_/A _11419_/B vssd1 vssd1 vccd1 vccd1 _11420_/B sky130_fd_sc_hd__nand2_1
X_14207_ _15663_/CLK _14207_/D vssd1 vssd1 vccd1 vccd1 _14207_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15187_ _15306_/CLK _15187_/D vssd1 vssd1 vccd1 vccd1 _15187_/Q sky130_fd_sc_hd__dfxtp_1
X_12399_ _06670_/A _12396_/X _06671_/A vssd1 vssd1 vccd1 vccd1 _12399_/X sky130_fd_sc_hd__o21a_1
XFILLER_113_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14138_ _14525_/CLK _14138_/D vssd1 vssd1 vccd1 vccd1 _14138_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_152_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14069_ _15142_/CLK _14069_/D vssd1 vssd1 vccd1 vccd1 _14069_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06960_ _06960_/A _06960_/B vssd1 vssd1 vccd1 vccd1 _06960_/Y sky130_fd_sc_hd__nor2_1
XFILLER_140_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_3_clk clkbuf_5_0_0_clk/X vssd1 vssd1 vccd1 vccd1 _15181_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_140_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06891_ _15398_/Q _06691_/Y _15397_/Q _06694_/Y _06890_/X vssd1 vssd1 vccd1 vccd1
+ _06891_/X sky130_fd_sc_hd__a221o_1
XFILLER_95_964 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08630_ _13494_/Q _08691_/B1 _08693_/B1 _13629_/Q vssd1 vssd1 vccd1 vccd1 _08630_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_55_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08561_ _13607_/Q _08749_/A2 _08750_/B1 _13639_/Q vssd1 vssd1 vccd1 vccd1 _08561_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_81_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07512_ _14742_/Q _13421_/Q _07529_/S vssd1 vssd1 vccd1 vccd1 _13421_/D sky130_fd_sc_hd__mux2_1
XFILLER_23_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08492_ _13774_/Q _12900_/S _08491_/X vssd1 vssd1 vccd1 vccd1 _13774_/D sky130_fd_sc_hd__o21a_1
XFILLER_63_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07443_ _13666_/Q _07483_/A2 _07483_/B1 _14694_/Q _07442_/X vssd1 vssd1 vccd1 vccd1
+ _07443_/X sky130_fd_sc_hd__a221o_1
XFILLER_50_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07374_ _07474_/B _07498_/C vssd1 vssd1 vccd1 vccd1 _07374_/X sky130_fd_sc_hd__and2b_1
XFILLER_10_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09113_ _09449_/A1 _09111_/X _09112_/X _09449_/B2 vssd1 vssd1 vccd1 vccd1 _09113_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_164_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09044_ _14010_/Q _13978_/Q _09047_/S vssd1 vssd1 vccd1 vccd1 _09044_/X sky130_fd_sc_hd__mux2_1
XFILLER_135_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09946_ _13080_/B2 _14306_/Q _09958_/S vssd1 vssd1 vccd1 vccd1 _14306_/D sky130_fd_sc_hd__mux2_1
XFILLER_38_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09877_ _13330_/A0 _14239_/Q _09892_/S vssd1 vssd1 vccd1 vccd1 _14239_/D sky130_fd_sc_hd__mux2_1
XTAP_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08828_ _13851_/Q _11860_/A1 _08846_/S vssd1 vssd1 vccd1 vccd1 _13851_/D sky130_fd_sc_hd__mux2_1
XFILLER_161_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08759_ _14596_/Q _14595_/Q _14597_/Q vssd1 vssd1 vccd1 vccd1 _08759_/X sky130_fd_sc_hd__a21o_1
XTAP_2614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11770_ _13345_/A0 _15198_/Q _11774_/S vssd1 vssd1 vccd1 vccd1 _15198_/D sky130_fd_sc_hd__mux2_1
XTAP_1924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10721_ _15023_/Q _10569_/B _10733_/A2 _14991_/Q _10732_/C1 vssd1 vssd1 vccd1 vccd1
+ _10721_/X sky130_fd_sc_hd__a221o_1
XFILLER_53_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13440_ _15393_/CLK _13440_/D vssd1 vssd1 vccd1 vccd1 _13440_/Q sky130_fd_sc_hd__dfxtp_1
X_10652_ _13728_/Q _10652_/B vssd1 vssd1 vccd1 vccd1 _10652_/X sky130_fd_sc_hd__and2_1
XFILLER_70_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13371_ _14474_/Q vssd1 vssd1 vccd1 vccd1 _14474_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_166_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10583_ _13714_/Q _10602_/B _10582_/X vssd1 vssd1 vccd1 vccd1 _10583_/X sky130_fd_sc_hd__a21o_1
XFILLER_167_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15110_ _15651_/CLK _15110_/D vssd1 vssd1 vccd1 vccd1 _15110_/Q sky130_fd_sc_hd__dfxtp_1
X_12322_ _14247_/Q _14279_/Q _14311_/Q _14343_/Q _12543_/S _12544_/A vssd1 vssd1 vccd1
+ vccd1 _12322_/X sky130_fd_sc_hd__mux4_1
XFILLER_166_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_295 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15041_ _15041_/CLK _15041_/D vssd1 vssd1 vccd1 vccd1 _15041_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_6_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12253_ _14244_/Q _14276_/Q _14308_/Q _14340_/Q _12154_/S _12253_/S1 vssd1 vssd1
+ vccd1 vccd1 _12253_/X sky130_fd_sc_hd__mux4_1
XFILLER_108_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11204_ _14928_/D _14927_/D _14929_/D vssd1 vssd1 vccd1 vccd1 _11204_/X sky130_fd_sc_hd__or3b_2
X_12184_ _14241_/Q _14273_/Q _14305_/Q _14337_/Q _12489_/S0 _12489_/S1 vssd1 vssd1
+ vccd1 vccd1 _12184_/X sky130_fd_sc_hd__mux4_1
XFILLER_122_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11135_ _11129_/A _11016_/X _11129_/Y vssd1 vssd1 vccd1 vccd1 _11189_/B sky130_fd_sc_hd__a21oi_1
XFILLER_68_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11066_ _10971_/Y _10992_/B _11318_/S vssd1 vssd1 vccd1 vccd1 _11066_/X sky130_fd_sc_hd__mux2_1
XFILLER_77_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10017_ _11838_/A1 _14375_/Q _10029_/S vssd1 vssd1 vccd1 vccd1 _14375_/D sky130_fd_sc_hd__mux2_1
XFILLER_77_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14825_ _15643_/CLK _14825_/D vssd1 vssd1 vccd1 vccd1 _14825_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14756_ _15624_/CLK _14756_/D vssd1 vssd1 vccd1 vccd1 _14756_/Q sky130_fd_sc_hd__dfxtp_4
X_11968_ _14006_/Q _13974_/Q _12079_/S vssd1 vssd1 vccd1 vccd1 _11969_/B sky130_fd_sc_hd__mux2_1
XFILLER_32_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13707_ _15507_/CLK _13707_/D vssd1 vssd1 vccd1 vccd1 _13707_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_177_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10919_ _14942_/Q _10944_/B _10918_/Y _11475_/B vssd1 vssd1 vccd1 vccd1 _14942_/D
+ sky130_fd_sc_hd__o22a_1
X_14687_ _15422_/CLK _14687_/D vssd1 vssd1 vccd1 vccd1 _14687_/Q sky130_fd_sc_hd__dfxtp_1
X_11899_ _14003_/Q _13971_/Q _12269_/S vssd1 vssd1 vccd1 vccd1 _11900_/B sky130_fd_sc_hd__mux2_1
XFILLER_60_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13638_ _13798_/CLK _13638_/D vssd1 vssd1 vccd1 vccd1 _13638_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_121_1103 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13569_ _13569_/CLK _13569_/D vssd1 vssd1 vccd1 vccd1 _13569_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_173_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_627 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15308_ _15527_/CLK _15308_/D vssd1 vssd1 vccd1 vccd1 _15308_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07090_ _14642_/Q _14674_/Q _07096_/S vssd1 vssd1 vccd1 vccd1 _07090_/X sky130_fd_sc_hd__mux2_1
XFILLER_8_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15239_ _15303_/CLK _15239_/D vssd1 vssd1 vccd1 vccd1 _15239_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_630 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09800_ _14166_/Q _11680_/A0 _09823_/S vssd1 vssd1 vccd1 vccd1 _14166_/D sky130_fd_sc_hd__mux2_1
Xfanout207 _09663_/Y vssd1 vssd1 vccd1 vccd1 _09690_/S sky130_fd_sc_hd__buf_12
Xfanout218 _08819_/Y vssd1 vssd1 vccd1 vccd1 _08851_/S sky130_fd_sc_hd__buf_12
XFILLER_119_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07992_ _13564_/Q _07992_/B vssd1 vssd1 vccd1 vccd1 _07992_/X sky130_fd_sc_hd__xor2_1
Xfanout229 _07713_/A vssd1 vssd1 vccd1 vccd1 _07750_/A sky130_fd_sc_hd__buf_6
XFILLER_101_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06943_ _06943_/A _06943_/B vssd1 vssd1 vccd1 vccd1 _06944_/D sky130_fd_sc_hd__nand2_1
XFILLER_140_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09731_ _14099_/Q _13319_/A0 _09757_/S vssd1 vssd1 vccd1 vccd1 _14099_/D sky130_fd_sc_hd__mux2_1
XFILLER_39_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09662_ _14713_/Q _09662_/B vssd1 vssd1 vccd1 vccd1 _11818_/A sky130_fd_sc_hd__or2_4
X_06874_ _06874_/A _13507_/Q vssd1 vssd1 vccd1 vccd1 _06879_/C sky130_fd_sc_hd__or2_1
XFILLER_95_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08613_ _13786_/Q _08626_/S _08612_/X vssd1 vssd1 vccd1 vccd1 _13786_/D sky130_fd_sc_hd__o21a_1
XFILLER_39_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09593_ _13969_/Q _11816_/A1 _09594_/S vssd1 vssd1 vccd1 vccd1 _13969_/D sky130_fd_sc_hd__mux2_1
XFILLER_27_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08544_ _15398_/Q _08748_/A2 _08736_/A2 _13443_/Q _08543_/X vssd1 vssd1 vccd1 vccd1
+ _08544_/X sky130_fd_sc_hd__a221o_1
XFILLER_82_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1003 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08475_ _13768_/Q _10764_/S _08470_/X _14609_/Q vssd1 vssd1 vccd1 vccd1 _13768_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_39_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07426_ _14658_/Q _07474_/B _07482_/C vssd1 vssd1 vccd1 vccd1 _07426_/X sky130_fd_sc_hd__and3_1
XFILLER_50_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07357_ _07230_/B _07231_/B _07356_/Y _07205_/X vssd1 vssd1 vccd1 vccd1 _07357_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_149_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07288_ _15506_/Q _07339_/S vssd1 vssd1 vccd1 vccd1 _07288_/Y sky130_fd_sc_hd__nand2b_2
XFILLER_136_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09027_ _09523_/A1 _09025_/X _09026_/X vssd1 vssd1 vccd1 vccd1 _09027_/X sky130_fd_sc_hd__a21o_1
XFILLER_108_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_47 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09929_ _13349_/A0 _14290_/Q _09930_/S vssd1 vssd1 vccd1 vccd1 _14290_/D sky130_fd_sc_hd__mux2_1
XFILLER_59_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12940_ _12563_/A _08852_/B _11743_/C _08405_/C vssd1 vssd1 vccd1 vccd1 _12940_/X
+ sky130_fd_sc_hd__o2bb2a_1
XTAP_3112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12871_ _14765_/Q _15399_/Q _12871_/S vssd1 vssd1 vccd1 vccd1 _15399_/D sky130_fd_sc_hd__mux2_1
XANTENNA_101 _15051_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_112 input8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_123 _08885_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14610_ _15501_/CLK _14610_/D vssd1 vssd1 vccd1 vccd1 _14610_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_2433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_134 _15344_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11822_ _15244_/Q _13322_/A0 _11849_/S vssd1 vssd1 vccd1 vccd1 _15244_/D sky130_fd_sc_hd__mux2_1
XTAP_2444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15590_ _15646_/CLK _15590_/D vssd1 vssd1 vccd1 vccd1 _15590_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11753_ _11861_/A1 _15181_/Q _11774_/S vssd1 vssd1 vccd1 vccd1 _15181_/D sky130_fd_sc_hd__mux2_1
X_14541_ _15672_/CLK _14541_/D vssd1 vssd1 vccd1 vccd1 _14541_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_516 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10704_ _15068_/Q _10714_/A2 _10701_/X _10703_/X vssd1 vssd1 vccd1 vccd1 _10704_/X
+ sky130_fd_sc_hd__o22a_1
XTAP_1787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11684_ _13326_/A0 _15115_/Q _11703_/S vssd1 vssd1 vccd1 vccd1 _15115_/D sky130_fd_sc_hd__mux2_1
X_14472_ _15301_/CLK _14472_/D vssd1 vssd1 vccd1 vccd1 _14472_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10635_ _14745_/Q _10634_/X _10650_/S vssd1 vssd1 vccd1 vccd1 _14745_/D sky130_fd_sc_hd__mux2_1
X_13423_ _15379_/CLK _13423_/D vssd1 vssd1 vccd1 vccd1 _13423_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_128_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13354_ _14457_/Q vssd1 vssd1 vccd1 vccd1 _14457_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_182_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10566_ _15075_/Q _10566_/B vssd1 vssd1 vccd1 vccd1 _14733_/D sky130_fd_sc_hd__or2_1
XFILLER_154_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_917 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12305_ _15291_/Q _15259_/Q _15227_/Q _15158_/Q _12541_/S _12544_/A vssd1 vssd1 vccd1
+ vccd1 _12306_/B sky130_fd_sc_hd__mux4_1
X_13285_ _14389_/Q _15617_/Q _13291_/S vssd1 vssd1 vccd1 vccd1 _15617_/D sky130_fd_sc_hd__mux2_1
XFILLER_127_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10497_ _10520_/A1 _13785_/Q _13753_/Q _10520_/B2 vssd1 vssd1 vccd1 vccd1 _10497_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_108_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12236_ _15288_/Q _15256_/Q _15224_/Q _15155_/Q _12499_/S _12486_/S1 vssd1 vssd1
+ vccd1 vccd1 _12237_/B sky130_fd_sc_hd__mux4_1
X_15024_ _15581_/CLK _15024_/D vssd1 vssd1 vccd1 vccd1 _15024_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12167_ _15285_/Q _15253_/Q _15221_/Q _15152_/Q _12154_/S _11992_/A vssd1 vssd1 vccd1
+ vccd1 _12168_/B sky130_fd_sc_hd__mux4_1
XFILLER_96_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11118_ _08233_/B _11114_/X _11117_/Y _11202_/A vssd1 vssd1 vccd1 vccd1 _11118_/X
+ sky130_fd_sc_hd__o211a_1
X_12098_ _15282_/Q _15250_/Q _15218_/Q _15149_/Q _12472_/S _12465_/S1 vssd1 vssd1
+ vccd1 vccd1 _12099_/B sky130_fd_sc_hd__mux4_1
XFILLER_68_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11049_ _11298_/A _11136_/B _11046_/X _11048_/Y _11043_/X vssd1 vssd1 vccd1 vccd1
+ _11050_/B sky130_fd_sc_hd__o221a_1
Xinput7 ext_read_data[15] vssd1 vssd1 vccd1 vccd1 input7/X sky130_fd_sc_hd__clkbuf_4
XFILLER_37_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14808_ _15626_/CLK _14808_/D vssd1 vssd1 vccd1 vccd1 _14808_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14739_ _15620_/CLK _14739_/D vssd1 vssd1 vccd1 vccd1 _14739_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_71_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08260_ _11351_/C1 _08249_/Y _08259_/Y _08232_/A _13714_/Q vssd1 vssd1 vccd1 vccd1
+ _13714_/D sky130_fd_sc_hd__a32o_1
XFILLER_178_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07211_ _15332_/Q _15488_/Q _07340_/S vssd1 vssd1 vccd1 vccd1 _07211_/X sky130_fd_sc_hd__mux2_4
X_08191_ _13682_/Q _11853_/A1 _08221_/S vssd1 vssd1 vccd1 vccd1 _13682_/D sky130_fd_sc_hd__mux2_1
XFILLER_186_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_733 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07142_ _14851_/Q _14843_/Q _08150_/S vssd1 vssd1 vccd1 vccd1 _07142_/X sky130_fd_sc_hd__mux2_1
XFILLER_119_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07073_ _07072_/X _13603_/Q _12764_/S vssd1 vssd1 vccd1 vccd1 _07073_/X sky130_fd_sc_hd__mux2_1
XFILLER_156_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07975_ _07984_/D _07974_/Y _07971_/A vssd1 vssd1 vccd1 vccd1 _07975_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_102_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06926_ _06920_/A _06918_/X _06922_/B _06925_/Y vssd1 vssd1 vccd1 vccd1 _06926_/X
+ sky130_fd_sc_hd__o2bb2a_1
X_09714_ _11761_/A0 _14084_/Q _09728_/S vssd1 vssd1 vccd1 vccd1 _14084_/D sky130_fd_sc_hd__mux2_1
XFILLER_132_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09645_ _14018_/Q _13082_/B2 _09660_/S vssd1 vssd1 vccd1 vccd1 _14018_/D sky130_fd_sc_hd__mux2_1
X_06857_ _07104_/C _08094_/S _06857_/C _14923_/Q vssd1 vssd1 vccd1 vccd1 _06857_/X
+ sky130_fd_sc_hd__or4b_4
XFILLER_16_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09576_ _13952_/Q _13078_/B2 _09589_/S vssd1 vssd1 vccd1 vccd1 _13952_/D sky130_fd_sc_hd__mux2_1
XTAP_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06788_ _06789_/B vssd1 vssd1 vccd1 vccd1 _06798_/C sky130_fd_sc_hd__inv_2
XTAP_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08527_ _15399_/Q _08748_/A2 _08514_/X _08526_/X vssd1 vssd1 vccd1 vccd1 _08527_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_150_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08458_ _13759_/Q _12900_/S _08426_/X _08457_/X vssd1 vssd1 vccd1 vccd1 _13759_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_50_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07409_ _13327_/A0 _13391_/Q _07481_/S vssd1 vssd1 vccd1 vccd1 _13391_/D sky130_fd_sc_hd__mux2_1
XFILLER_11_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08389_ _08388_/X _11327_/A _11346_/A2 _13728_/Q vssd1 vssd1 vccd1 vccd1 _13728_/D
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_51_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xwire438 wire438/A vssd1 vssd1 vccd1 vccd1 wire438/X sky130_fd_sc_hd__buf_4
X_10420_ _10420_/A _10420_/B vssd1 vssd1 vccd1 vccd1 _11639_/A sky130_fd_sc_hd__nand2_2
XFILLER_167_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10351_ _13252_/A _13251_/B vssd1 vssd1 vccd1 vccd1 _10420_/A sky130_fd_sc_hd__or2_2
X_13070_ _12972_/X _13104_/A2 _13104_/B1 _13328_/A0 vssd1 vssd1 vccd1 vccd1 _13070_/X
+ sky130_fd_sc_hd__a22o_1
X_10282_ _14667_/Q _14820_/Q _10715_/S vssd1 vssd1 vccd1 vccd1 _14667_/D sky130_fd_sc_hd__mux2_1
XFILLER_124_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12021_ _12573_/A _12021_/B _12021_/C vssd1 vssd1 vccd1 vccd1 _12021_/X sky130_fd_sc_hd__and3_2
XFILLER_151_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout560 _09551_/S vssd1 vssd1 vccd1 vccd1 _09481_/S sky130_fd_sc_hd__buf_8
Xfanout571 _08451_/A vssd1 vssd1 vccd1 vccd1 _12455_/C1 sky130_fd_sc_hd__clkbuf_16
XFILLER_93_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout582 _12061_/A vssd1 vssd1 vccd1 vccd1 _12253_/S1 sky130_fd_sc_hd__buf_12
XFILLER_120_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout593 fanout600/X vssd1 vssd1 vccd1 vccd1 _12406_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_58_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13972_ _15125_/CLK _13972_/D vssd1 vssd1 vccd1 vccd1 _13972_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12923_ _15451_/Q _15637_/Q _12929_/S vssd1 vssd1 vccd1 vccd1 _15451_/D sky130_fd_sc_hd__mux2_1
XFILLER_46_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15642_ _15643_/CLK _15642_/D vssd1 vssd1 vccd1 vccd1 _15642_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12854_ _14748_/Q _15382_/Q _12866_/S vssd1 vssd1 vccd1 vccd1 _15382_/D sky130_fd_sc_hd__mux2_1
XTAP_2241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11805_ _15228_/Q _11838_/A1 _11817_/S vssd1 vssd1 vccd1 vccd1 _15228_/D sky130_fd_sc_hd__mux2_1
XTAP_2274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15573_ _15591_/CLK _15573_/D vssd1 vssd1 vccd1 vccd1 _15573_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12785_ _13604_/Q _12785_/B vssd1 vssd1 vccd1 vccd1 _12785_/X sky130_fd_sc_hd__or2_1
XFILLER_15_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14524_ _15655_/CLK _14524_/D vssd1 vssd1 vccd1 vccd1 _14524_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_644 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11736_ _15165_/Q _11877_/A1 _11741_/S vssd1 vssd1 vccd1 vccd1 _15165_/D sky130_fd_sc_hd__mux2_1
XFILLER_41_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14455_ _14606_/CLK _14455_/D vssd1 vssd1 vccd1 vccd1 _14455_/Q sky130_fd_sc_hd__dfxtp_1
X_11667_ _13342_/A0 _15099_/Q _11675_/S vssd1 vssd1 vccd1 vccd1 _15099_/D sky130_fd_sc_hd__mux2_1
X_13406_ _15672_/CLK _13406_/D vssd1 vssd1 vccd1 vccd1 _13406_/Q sky130_fd_sc_hd__dfxtp_1
X_10618_ _14970_/Q _10718_/A2 _10722_/B1 _14938_/Q _10617_/X vssd1 vssd1 vccd1 vccd1
+ _10618_/X sky130_fd_sc_hd__a221o_1
X_11598_ _11598_/A _11598_/B vssd1 vssd1 vccd1 vccd1 _11599_/B sky130_fd_sc_hd__nor2_1
X_14386_ _14420_/CLK _14386_/D vssd1 vssd1 vccd1 vccd1 _14386_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_183_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13337_ _13337_/A0 _15667_/Q _13350_/S vssd1 vssd1 vccd1 vccd1 _15667_/D sky130_fd_sc_hd__mux2_1
X_10549_ _11371_/A _13165_/B vssd1 vssd1 vccd1 vccd1 _10556_/B sky130_fd_sc_hd__xnor2_1
XFILLER_115_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13268_ _15352_/Q _15599_/Q _13288_/S vssd1 vssd1 vccd1 vccd1 _15599_/D sky130_fd_sc_hd__mux2_1
XFILLER_29_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15007_ _15577_/CLK _15007_/D vssd1 vssd1 vccd1 vccd1 _15007_/Q sky130_fd_sc_hd__dfxtp_1
X_12219_ _13889_/Q _14404_/Q _12476_/S vssd1 vssd1 vccd1 vccd1 _12219_/X sky130_fd_sc_hd__mux2_1
X_13199_ _13217_/A _13199_/B vssd1 vssd1 vccd1 vccd1 _13199_/X sky130_fd_sc_hd__or2_1
XFILLER_111_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_1079 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_1_1_0_clk clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 clkbuf_1_1_1_clk/A sky130_fd_sc_hd__clkbuf_8
X_07760_ _13504_/Q _07765_/C vssd1 vssd1 vccd1 vccd1 _07760_/Y sky130_fd_sc_hd__nor2_1
XFILLER_110_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06711_ _13466_/Q vssd1 vssd1 vccd1 vccd1 _06711_/Y sky130_fd_sc_hd__inv_2
XFILLER_37_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07691_ _07713_/A _07691_/B vssd1 vssd1 vccd1 vccd1 _07691_/Y sky130_fd_sc_hd__nand2_1
XFILLER_53_915 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_200_clk clkbuf_5_17_0_clk/X vssd1 vssd1 vccd1 vccd1 _15142_/CLK sky130_fd_sc_hd__clkbuf_16
X_09430_ _09449_/A1 _09428_/X _09429_/X _09449_/B2 vssd1 vssd1 vccd1 vccd1 _09430_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_80_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09361_ _13897_/Q _09522_/A2 _09519_/B1 _14412_/Q _08507_/A vssd1 vssd1 vccd1 vccd1
+ _09361_/X sky130_fd_sc_hd__a221o_1
XFILLER_24_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_1052 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08312_ _07307_/X _10523_/A2 _08311_/X vssd1 vssd1 vccd1 vccd1 _11419_/A sky130_fd_sc_hd__a21oi_4
X_09292_ _14022_/Q _13990_/Q _09484_/S vssd1 vssd1 vccd1 vccd1 _09292_/X sky130_fd_sc_hd__mux2_1
XFILLER_32_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_12 _10684_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_23 _13779_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08243_ _11356_/B _11349_/B vssd1 vssd1 vccd1 vccd1 _11362_/C sky130_fd_sc_hd__nor2_2
XFILLER_166_828 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_34 _14760_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_45 input23/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_56 _07193_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_67 _07131_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_78 _07159_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08174_ _13674_/Q _10285_/S _08155_/X _08173_/X vssd1 vssd1 vccd1 vccd1 _13674_/D
+ sky130_fd_sc_hd__o22a_1
XANTENNA_89 _07042_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07125_ _07131_/A _07125_/B vssd1 vssd1 vccd1 vccd1 _07125_/X sky130_fd_sc_hd__and2_4
XFILLER_107_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07056_ _07055_/X _14751_/Q _07077_/S vssd1 vssd1 vccd1 vccd1 _13597_/D sky130_fd_sc_hd__mux2_1
XFILLER_173_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07958_ _13555_/Q _07958_/B vssd1 vssd1 vccd1 vccd1 _07959_/B sky130_fd_sc_hd__xor2_1
XFILLER_28_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06909_ _06906_/X _06907_/X _06908_/X vssd1 vssd1 vccd1 vccd1 _06909_/X sky130_fd_sc_hd__a21o_1
XFILLER_28_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07889_ _13537_/Q _07900_/C vssd1 vssd1 vccd1 vccd1 _07890_/B sky130_fd_sc_hd__xnor2_1
XFILLER_44_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09628_ _14002_/Q _11883_/A1 _09628_/S vssd1 vssd1 vccd1 vccd1 _14002_/D sky130_fd_sc_hd__mux2_1
XFILLER_44_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xcore_648 vssd1 vssd1 vccd1 vccd1 core_648/HI ext_address[0] sky130_fd_sc_hd__conb_1
XFILLER_43_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09559_ _08507_/Y _09555_/X _09556_/X _09558_/X vssd1 vssd1 vccd1 vccd1 _09559_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_71_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12570_ _12563_/X _12565_/X _12567_/X _12569_/X _06671_/A vssd1 vssd1 vccd1 vccd1
+ _12570_/X sky130_fd_sc_hd__o221a_1
XFILLER_52_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11521_ _11521_/A _11521_/B vssd1 vssd1 vccd1 vccd1 _11522_/B sky130_fd_sc_hd__or2_1
XFILLER_12_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11452_ _11459_/B _11452_/B vssd1 vssd1 vccd1 vccd1 _11452_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_156_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14240_ _15285_/CLK _14240_/D vssd1 vssd1 vccd1 vccd1 _14240_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10403_ _10403_/A _13159_/B vssd1 vssd1 vccd1 vccd1 _10403_/Y sky130_fd_sc_hd__nor2_1
XFILLER_165_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14171_ _15212_/CLK _14171_/D vssd1 vssd1 vccd1 vccd1 _14171_/Q sky130_fd_sc_hd__dfxtp_1
X_11383_ _11383_/A _11383_/B vssd1 vssd1 vccd1 vccd1 _11384_/B sky130_fd_sc_hd__and2_1
XFILLER_139_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_596 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13122_ hold1/A _10871_/S _09829_/B _08402_/X vssd1 vssd1 vccd1 vccd1 _15531_/D sky130_fd_sc_hd__o22a_1
X_10334_ _14719_/Q _14912_/Q _10343_/S vssd1 vssd1 vccd1 vccd1 _14719_/D sky130_fd_sc_hd__mux2_1
XFILLER_125_758 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13053_ _15494_/Q _13105_/A2 _13105_/B1 _13052_/X vssd1 vssd1 vccd1 vccd1 _15494_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_97_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10265_ _14650_/Q _14803_/Q _10730_/S vssd1 vssd1 vccd1 vccd1 _14650_/D sky130_fd_sc_hd__mux2_1
XFILLER_127_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_599 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12004_ _12000_/X _12001_/X _12594_/S vssd1 vssd1 vccd1 vccd1 _12004_/X sky130_fd_sc_hd__mux2_1
XFILLER_78_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10196_ _11816_/A1 _14580_/Q _10197_/S vssd1 vssd1 vccd1 vccd1 _14580_/D sky130_fd_sc_hd__mux2_1
XFILLER_121_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout390 _11380_/A vssd1 vssd1 vccd1 vccd1 _11199_/A sky130_fd_sc_hd__buf_6
X_13955_ _15657_/CLK _13955_/D vssd1 vssd1 vccd1 vccd1 _13955_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12906_ _15434_/Q _15620_/Q _12906_/S vssd1 vssd1 vccd1 vccd1 _15434_/D sky130_fd_sc_hd__mux2_1
XFILLER_61_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13886_ _15285_/CLK _13886_/D vssd1 vssd1 vccd1 vccd1 _13886_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_46_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15625_ _15626_/CLK _15625_/D vssd1 vssd1 vccd1 vccd1 _15625_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12837_ _13444_/Q _12640_/S _12835_/X _12836_/X _12759_/B vssd1 vssd1 vccd1 vccd1
+ _12837_/X sky130_fd_sc_hd__o221a_1
XTAP_2071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15556_ _15556_/CLK _15556_/D vssd1 vssd1 vccd1 vccd1 _15556_/Q sky130_fd_sc_hd__dfxtp_1
X_12768_ _15357_/Q _12767_/C _15358_/Q vssd1 vssd1 vccd1 vccd1 _12769_/B sky130_fd_sc_hd__a21oi_1
XTAP_1381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14507_ _14510_/CLK _14507_/D vssd1 vssd1 vccd1 vccd1 _14507_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_175_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11719_ _15148_/Q _13327_/A0 _11741_/S vssd1 vssd1 vccd1 vccd1 _15148_/D sky130_fd_sc_hd__mux2_1
XFILLER_175_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15487_ _15519_/CLK _15487_/D vssd1 vssd1 vccd1 vccd1 _15487_/Q sky130_fd_sc_hd__dfxtp_1
X_12699_ _12737_/A _12699_/B vssd1 vssd1 vccd1 vccd1 _12699_/X sky130_fd_sc_hd__or2_1
XFILLER_30_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14438_ _15108_/CLK _14438_/D vssd1 vssd1 vccd1 vccd1 _14438_/Q sky130_fd_sc_hd__dfxtp_1
Xinput10 ext_read_data[18] vssd1 vssd1 vccd1 vccd1 input10/X sky130_fd_sc_hd__buf_6
XFILLER_174_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput21 ext_read_data[28] vssd1 vssd1 vccd1 vccd1 input21/X sky130_fd_sc_hd__buf_8
Xinput32 ext_read_data[9] vssd1 vssd1 vccd1 vccd1 input32/X sky130_fd_sc_hd__buf_4
Xclkbuf_leaf_249_clk clkbuf_5_1_0_clk/X vssd1 vssd1 vccd1 vccd1 _15253_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_122_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14369_ _15674_/CLK _14369_/D vssd1 vssd1 vccd1 vccd1 _14369_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_155_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_875 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08930_ _15275_/Q _15243_/Q _15211_/Q _15142_/Q _09484_/S _08519_/A vssd1 vssd1 vccd1
+ vccd1 _08930_/X sky130_fd_sc_hd__mux4_1
XFILLER_69_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08861_ _13882_/Q _13326_/A0 _08880_/S vssd1 vssd1 vccd1 vccd1 _13882_/D sky130_fd_sc_hd__mux2_1
XFILLER_123_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07812_ _14741_/Q _07816_/A _07811_/Y _07938_/C1 vssd1 vssd1 vccd1 vccd1 _13516_/D
+ sky130_fd_sc_hd__o211a_1
X_08792_ _12967_/A1 _13818_/Q _08811_/S vssd1 vssd1 vccd1 vccd1 _13818_/D sky130_fd_sc_hd__mux2_1
XFILLER_123_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07743_ _07750_/A _07743_/B vssd1 vssd1 vccd1 vccd1 _07743_/Y sky130_fd_sc_hd__nand2_1
XFILLER_38_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07674_ _14737_/Q _07676_/A _07673_/Y _08084_/C1 vssd1 vssd1 vccd1 vccd1 _13480_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_65_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09413_ _14381_/Q _15197_/Q _13836_/Q _14575_/Q _09190_/S _09446_/A1 vssd1 vssd1
+ vccd1 vccd1 _09414_/B sky130_fd_sc_hd__mux4_1
XFILLER_34_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09344_ _15097_/Q _08540_/B _09343_/X _08501_/A vssd1 vssd1 vccd1 vccd1 _09344_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_139_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09275_ _09554_/A _09275_/B _09275_/C vssd1 vssd1 vccd1 vccd1 _09275_/X sky130_fd_sc_hd__and3_1
XFILLER_166_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08226_ _08240_/A _13803_/Q _13771_/Q _08237_/A vssd1 vssd1 vccd1 vccd1 _08226_/X
+ sky130_fd_sc_hd__a22o_2
XFILLER_101_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08157_ _08185_/A _08157_/B vssd1 vssd1 vccd1 vccd1 _08157_/X sky130_fd_sc_hd__and2_1
XFILLER_146_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07108_ _14830_/Q _07115_/B _07163_/A vssd1 vssd1 vccd1 vccd1 _07108_/X sky130_fd_sc_hd__and3_4
XFILLER_134_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08088_ _14737_/Q _08083_/A _08087_/X vssd1 vssd1 vccd1 vccd1 _13647_/D sky130_fd_sc_hd__o21ba_1
XFILLER_134_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07039_ _14625_/Q _14657_/Q _07078_/S vssd1 vssd1 vccd1 vccd1 _07039_/X sky130_fd_sc_hd__mux2_1
XFILLER_122_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10050_ _14407_/Q _11761_/A0 _10064_/S vssd1 vssd1 vccd1 vccd1 _14407_/D sky130_fd_sc_hd__mux2_1
XFILLER_88_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_915 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13740_ _14863_/CLK _13740_/D vssd1 vssd1 vccd1 vccd1 _14929_/D sky130_fd_sc_hd__dfxtp_4
X_10952_ _14961_/Q _10894_/X _10951_/Y _13251_/B vssd1 vssd1 vccd1 vccd1 _14961_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_43_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_5_17_0_clk clkbuf_4_8_0_clk/X vssd1 vssd1 vccd1 vccd1 clkbuf_5_17_0_clk/X
+ sky130_fd_sc_hd__clkbuf_8
X_13671_ _15438_/CLK _13671_/D vssd1 vssd1 vccd1 vccd1 _13671_/Q sky130_fd_sc_hd__dfxtp_1
X_10883_ _14915_/Q _15546_/Q _13134_/A vssd1 vssd1 vccd1 vccd1 _14915_/D sky130_fd_sc_hd__mux2_1
X_15410_ _15599_/CLK _15410_/D vssd1 vssd1 vccd1 vccd1 _15410_/Q sky130_fd_sc_hd__dfxtp_2
X_12622_ _12622_/A _15615_/D vssd1 vssd1 vccd1 vccd1 _12622_/X sky130_fd_sc_hd__or2_2
XFILLER_106_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15341_ _15429_/CLK _15341_/D vssd1 vssd1 vccd1 vccd1 _15341_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_8_602 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12553_ _14483_/Q _14451_/Q _13872_/Q _14225_/Q _12430_/S _12567_/A vssd1 vssd1 vccd1
+ vccd1 _12553_/X sky130_fd_sc_hd__mux4_1
XFILLER_106_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11504_ _11492_/A _11502_/Y _11503_/X _11482_/X vssd1 vssd1 vccd1 vccd1 _11507_/A
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_12_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15272_ _15304_/CLK _15272_/D vssd1 vssd1 vccd1 vccd1 _15272_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12484_ _14480_/Q _14448_/Q _13869_/Q _14222_/Q _12489_/S0 _12489_/S1 vssd1 vssd1
+ vccd1 vccd1 _12484_/X sky130_fd_sc_hd__mux4_1
XFILLER_185_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14223_ _15300_/CLK _14223_/D vssd1 vssd1 vccd1 vccd1 _14223_/Q sky130_fd_sc_hd__dfxtp_1
X_11435_ _11434_/Y _15052_/Q _11474_/S vssd1 vssd1 vccd1 vccd1 _15052_/D sky130_fd_sc_hd__mux2_1
XFILLER_7_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14154_ _15672_/CLK _14154_/D vssd1 vssd1 vccd1 vccd1 _14154_/Q sky130_fd_sc_hd__dfxtp_1
X_11366_ _10551_/B _11360_/B _11359_/A vssd1 vssd1 vccd1 vccd1 _11368_/B sky130_fd_sc_hd__a21o_1
XFILLER_152_341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10317_ _14702_/Q _14887_/Q _10710_/S vssd1 vssd1 vccd1 vccd1 _14702_/D sky130_fd_sc_hd__mux2_1
X_13105_ _15520_/Q _13105_/A2 _13105_/B1 _13104_/X vssd1 vssd1 vccd1 vccd1 _15520_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_153_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14085_ _15668_/CLK _14085_/D vssd1 vssd1 vccd1 vccd1 _14085_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_112_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11297_ _11266_/X _11296_/Y _11297_/S vssd1 vssd1 vccd1 vccd1 _11347_/B sky130_fd_sc_hd__mux2_1
XFILLER_152_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10248_ _14633_/Q _14786_/Q _10665_/S vssd1 vssd1 vccd1 vccd1 _14633_/D sky130_fd_sc_hd__mux2_1
XTAP_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13036_ _07496_/X _13039_/A2 _13035_/X _12944_/A vssd1 vssd1 vccd1 vccd1 _13036_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_78_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10179_ _13332_/A0 _14563_/Q _10192_/S vssd1 vssd1 vccd1 vccd1 _14563_/D sky130_fd_sc_hd__mux2_1
XFILLER_26_1079 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_1098 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14987_ _14988_/CLK _14987_/D vssd1 vssd1 vccd1 vccd1 _14987_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13938_ _15650_/CLK _13938_/D vssd1 vssd1 vccd1 vccd1 _13938_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13869_ _15556_/CLK _13869_/D vssd1 vssd1 vccd1 vccd1 _13869_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15608_ _15608_/CLK _15608_/D vssd1 vssd1 vccd1 vccd1 _15608_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07390_ _14649_/Q _07498_/B _07498_/C vssd1 vssd1 vccd1 vccd1 _07390_/X sky130_fd_sc_hd__and3_1
XFILLER_148_603 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15539_ _15617_/CLK _15539_/D vssd1 vssd1 vccd1 vccd1 _15539_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_147_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09060_ _14075_/Q _09445_/A2 _09522_/B1 _14043_/Q _09391_/A vssd1 vssd1 vccd1 vccd1
+ _09060_/X sky130_fd_sc_hd__a221o_1
XFILLER_72_1099 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_850 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08011_ _08022_/B _08011_/B vssd1 vssd1 vccd1 vccd1 _08011_/Y sky130_fd_sc_hd__nand2_1
XFILLER_129_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09962_ _13349_/A0 _14322_/Q _09963_/S vssd1 vssd1 vccd1 vccd1 _14322_/D sky130_fd_sc_hd__mux2_1
XFILLER_104_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08913_ _08510_/B _08909_/X _08912_/X _08908_/X vssd1 vssd1 vccd1 vccd1 _08926_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_103_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09893_ _13346_/A0 _14255_/Q _09897_/S vssd1 vssd1 vccd1 vccd1 _14255_/D sky130_fd_sc_hd__mux2_1
XTAP_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08844_ _13867_/Q _13343_/A0 _08846_/S vssd1 vssd1 vccd1 vccd1 _13867_/D sky130_fd_sc_hd__mux2_1
XFILLER_84_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08775_ _08757_/Y _08766_/X _08774_/X _10871_/S vssd1 vssd1 vccd1 vccd1 _08775_/X
+ sky130_fd_sc_hd__o31a_2
XFILLER_26_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07726_ _14751_/Q _07750_/A _07725_/Y _07987_/C1 vssd1 vssd1 vccd1 vccd1 _13494_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_2818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07657_ _14765_/Q _07644_/A _07656_/Y _08016_/C1 vssd1 vssd1 vccd1 vccd1 _13476_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_25_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07588_ _13458_/Q _13457_/Q _13456_/Q _07588_/D vssd1 vssd1 vccd1 vccd1 _07603_/C
+ sky130_fd_sc_hd__and4_4
XFILLER_80_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09327_ _15294_/Q _15262_/Q _15230_/Q _15161_/Q _09469_/S _09546_/S1 vssd1 vssd1
+ vccd1 vccd1 _09327_/X sky130_fd_sc_hd__mux4_1
XFILLER_182_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09258_ _09242_/X _09245_/X _09252_/X _09257_/X vssd1 vssd1 vccd1 vccd1 _09258_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_127_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08209_ _13700_/Q _13338_/A0 _08221_/S vssd1 vssd1 vccd1 vccd1 _13700_/D sky130_fd_sc_hd__mux2_1
X_09189_ _09427_/A1 _09187_/X _09188_/X vssd1 vssd1 vccd1 vccd1 _09189_/X sky130_fd_sc_hd__a21o_1
XFILLER_147_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11220_ _10366_/A _15008_/Q _11232_/S vssd1 vssd1 vccd1 vccd1 _15008_/D sky130_fd_sc_hd__mux2_1
XFILLER_5_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11151_ _11199_/A _11195_/B vssd1 vssd1 vccd1 vccd1 _11151_/Y sky130_fd_sc_hd__nand2_1
XFILLER_135_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10102_ _14488_/Q _14736_/Q _10131_/S vssd1 vssd1 vccd1 vccd1 _14488_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11082_ _11082_/A vssd1 vssd1 vccd1 vccd1 _11082_/Y sky130_fd_sc_hd__inv_2
XFILLER_122_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10033_ _14390_/Q _13319_/A0 _10059_/S vssd1 vssd1 vccd1 vccd1 _14390_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14910_ _15199_/CLK _14910_/D vssd1 vssd1 vccd1 vccd1 _14910_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_5_0_0_clk clkbuf_5_1_0_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_5_0_0_clk/X sky130_fd_sc_hd__clkbuf_8
X_14841_ _15508_/CLK _14841_/D vssd1 vssd1 vccd1 vccd1 _14841_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14772_ _15589_/CLK _14772_/D vssd1 vssd1 vccd1 vccd1 _14772_/Q sky130_fd_sc_hd__dfxtp_1
X_11984_ _12260_/A _11984_/B vssd1 vssd1 vccd1 vccd1 _11984_/X sky130_fd_sc_hd__or2_1
XFILLER_112_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13723_ _15020_/CLK _13723_/D vssd1 vssd1 vccd1 vccd1 _13723_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_182_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10935_ _14951_/Q _10948_/B _10934_/Y _13220_/B vssd1 vssd1 vccd1 vccd1 _14951_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_31_203 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13654_ _15620_/CLK _13654_/D vssd1 vssd1 vccd1 vccd1 _13654_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_143_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10866_ _14898_/Q _15535_/Q _13138_/S vssd1 vssd1 vccd1 vccd1 _14898_/D sky130_fd_sc_hd__mux2_1
XFILLER_176_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12605_ _12617_/S _12605_/B vssd1 vssd1 vccd1 vccd1 _12605_/X sky130_fd_sc_hd__or2_1
XPHY_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13585_ _15429_/CLK _13585_/D vssd1 vssd1 vccd1 vccd1 _13585_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10797_ _14829_/Q _15461_/Q _12933_/S vssd1 vssd1 vccd1 vccd1 _14829_/D sky130_fd_sc_hd__mux2_1
XFILLER_129_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15324_ _15324_/CLK _15324_/D vssd1 vssd1 vccd1 vccd1 _15324_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_185_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12536_ _12536_/A _12536_/B vssd1 vssd1 vccd1 vccd1 _12536_/X sky130_fd_sc_hd__or2_1
XFILLER_129_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_1050 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15255_ _15287_/CLK _15255_/D vssd1 vssd1 vccd1 vccd1 _15255_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_157_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12467_ _12490_/A _12467_/B vssd1 vssd1 vccd1 vccd1 _12467_/X sky130_fd_sc_hd__or2_1
XFILLER_144_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14206_ _15556_/CLK _14206_/D vssd1 vssd1 vccd1 vccd1 _14206_/Q sky130_fd_sc_hd__dfxtp_1
X_11418_ _11419_/A _11419_/B vssd1 vssd1 vccd1 vccd1 _11418_/X sky130_fd_sc_hd__and2_1
XFILLER_172_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15186_ _15287_/CLK _15186_/D vssd1 vssd1 vccd1 vccd1 _15186_/Q sky130_fd_sc_hd__dfxtp_1
X_12398_ _12594_/S _12398_/B vssd1 vssd1 vccd1 vccd1 _12398_/X sky130_fd_sc_hd__or2_1
XFILLER_126_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14137_ _15655_/CLK _14137_/D vssd1 vssd1 vccd1 vccd1 _14137_/Q sky130_fd_sc_hd__dfxtp_1
X_11349_ _11349_/A _11349_/B _11349_/C vssd1 vssd1 vccd1 vccd1 _11349_/X sky130_fd_sc_hd__and3_1
XFILLER_125_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_682 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14068_ _15077_/CLK _14068_/D vssd1 vssd1 vccd1 vccd1 _14068_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13019_ _15486_/Q _13119_/S _13025_/B1 _13018_/X vssd1 vssd1 vccd1 vccd1 _15486_/D
+ sky130_fd_sc_hd__a22o_1
X_06890_ _06929_/A _06889_/X _06884_/X vssd1 vssd1 vccd1 vccd1 _06890_/X sky130_fd_sc_hd__o21a_1
XFILLER_95_976 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08560_ _13778_/Q _08573_/S _08559_/X vssd1 vssd1 vccd1 vccd1 _13778_/D sky130_fd_sc_hd__o21a_1
X_07511_ _14741_/Q _13420_/Q _07535_/S vssd1 vssd1 vccd1 vccd1 _13420_/D sky130_fd_sc_hd__mux2_1
X_08491_ _08457_/A _08477_/X _08490_/X _13120_/S vssd1 vssd1 vccd1 vccd1 _08491_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_81_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07442_ _14662_/Q _07474_/B _07482_/C vssd1 vssd1 vccd1 vccd1 _07442_/X sky130_fd_sc_hd__and3_1
XFILLER_22_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07373_ _07498_/B _07498_/C vssd1 vssd1 vccd1 vccd1 _07373_/X sky130_fd_sc_hd__or2_2
XFILLER_176_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_742 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09112_ _14528_/Q _14141_/Q _14173_/Q _14109_/Q _09190_/S _09429_/S1 vssd1 vssd1
+ vccd1 vccd1 _09112_/X sky130_fd_sc_hd__mux4_1
XFILLER_176_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09043_ _09449_/A1 _09041_/X _09042_/X _09449_/B2 _09040_/X vssd1 vssd1 vccd1 vccd1
+ _09043_/X sky130_fd_sc_hd__a221o_4
XFILLER_164_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_300 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09945_ _13078_/B2 _14305_/Q _09958_/S vssd1 vssd1 vccd1 vccd1 _14305_/D sky130_fd_sc_hd__mux2_1
XFILLER_86_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09876_ _13072_/B2 _14238_/Q _09892_/S vssd1 vssd1 vccd1 vccd1 _14238_/D sky130_fd_sc_hd__mux2_1
XFILLER_135_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08827_ _13850_/Q _12967_/A1 _08846_/S vssd1 vssd1 vccd1 vccd1 _13850_/D sky130_fd_sc_hd__mux2_1
XFILLER_18_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08758_ _14596_/Q _08400_/C _08465_/X vssd1 vssd1 vccd1 vccd1 _08758_/X sky130_fd_sc_hd__a21o_1
XTAP_2615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07709_ _13490_/Q _13489_/Q _07732_/A vssd1 vssd1 vccd1 vccd1 _07712_/B sky130_fd_sc_hd__and3_2
XTAP_1903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08689_ _13797_/Q _12927_/S _08688_/X vssd1 vssd1 vccd1 vccd1 _13797_/D sky130_fd_sc_hd__o21a_1
XTAP_1925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10720_ _14762_/Q _10719_/X _10735_/S vssd1 vssd1 vccd1 vccd1 _14762_/D sky130_fd_sc_hd__mux2_1
XFILLER_13_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10651_ _15009_/Q _10717_/A2 _10722_/B1 _14945_/Q _10732_/C1 vssd1 vssd1 vccd1 vccd1
+ _10651_/X sky130_fd_sc_hd__a221o_1
XFILLER_16_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_1083 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13370_ _14473_/Q vssd1 vssd1 vccd1 vccd1 _14473_/D sky130_fd_sc_hd__clkbuf_2
X_10582_ _15554_/Q _10731_/B _10733_/B1 _14931_/Q vssd1 vssd1 vccd1 vccd1 _10582_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_142_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12321_ _15324_/Q _13149_/S _12320_/X vssd1 vssd1 vccd1 vccd1 _15324_/D sky130_fd_sc_hd__a21o_1
XFILLER_155_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15040_ _15042_/CLK _15040_/D vssd1 vssd1 vccd1 vccd1 _15040_/Q sky130_fd_sc_hd__dfxtp_1
X_12252_ _15321_/Q _13105_/A2 _12251_/X vssd1 vssd1 vccd1 vccd1 _15321_/D sky130_fd_sc_hd__a21o_1
XFILLER_79_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11203_ _14993_/Q _10984_/Y _11202_/X _13251_/B vssd1 vssd1 vccd1 vccd1 _14993_/D
+ sky130_fd_sc_hd__a22o_1
X_12183_ _15318_/Q _13081_/A2 _12182_/X vssd1 vssd1 vccd1 vccd1 _15318_/D sky130_fd_sc_hd__a21o_1
XFILLER_123_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11134_ _14970_/Q _10984_/Y _11131_/Y _11133_/X vssd1 vssd1 vccd1 vccd1 _14970_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_77_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11065_ _10985_/Y _10991_/Y _11330_/A vssd1 vssd1 vccd1 vccd1 _11065_/X sky130_fd_sc_hd__mux2_1
XFILLER_77_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10016_ _11870_/A1 _14374_/Q _10029_/S vssd1 vssd1 vccd1 vccd1 _14374_/D sky130_fd_sc_hd__mux2_1
XFILLER_76_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14824_ _15643_/CLK _14824_/D vssd1 vssd1 vccd1 vccd1 _14824_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14755_ _15624_/CLK _14755_/D vssd1 vssd1 vccd1 vccd1 _14755_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_63_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11967_ _12500_/A1 _11966_/X _12582_/A vssd1 vssd1 vccd1 vccd1 _11967_/X sky130_fd_sc_hd__a21o_1
XFILLER_91_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13706_ _14405_/CLK _13706_/D vssd1 vssd1 vccd1 vccd1 _13706_/Q sky130_fd_sc_hd__dfxtp_1
X_10918_ _11457_/A _10944_/B vssd1 vssd1 vccd1 vccd1 _10918_/Y sky130_fd_sc_hd__nand2_1
X_14686_ _15607_/CLK _14686_/D vssd1 vssd1 vccd1 vccd1 _14686_/Q sky130_fd_sc_hd__dfxtp_1
X_11898_ _12500_/A1 _11897_/X _12260_/A vssd1 vssd1 vccd1 vccd1 _11898_/X sky130_fd_sc_hd__a21o_1
X_13637_ _14511_/CLK _13637_/D vssd1 vssd1 vccd1 vccd1 _13637_/Q sky130_fd_sc_hd__dfxtp_1
X_10849_ _14881_/Q _13787_/Q _12929_/S vssd1 vssd1 vccd1 vccd1 _14881_/D sky130_fd_sc_hd__mux2_1
XFILLER_60_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13568_ _13569_/CLK _13568_/D vssd1 vssd1 vccd1 vccd1 _13568_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_185_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15307_ _15536_/CLK _15307_/D vssd1 vssd1 vccd1 vccd1 _15307_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_185_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12519_ _12615_/A1 _12518_/X _12617_/S vssd1 vssd1 vccd1 vccd1 _12519_/X sky130_fd_sc_hd__a21o_1
XFILLER_118_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13499_ _13565_/CLK _13499_/D vssd1 vssd1 vccd1 vccd1 _13499_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_67_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15238_ _15335_/CLK _15238_/D vssd1 vssd1 vccd1 vccd1 _15238_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_173_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_661 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15169_ _15335_/CLK _15169_/D vssd1 vssd1 vccd1 vccd1 _15169_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_158_1071 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout208 _09663_/Y vssd1 vssd1 vccd1 vccd1 _09695_/S sky130_fd_sc_hd__buf_12
XFILLER_141_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout219 _08784_/X vssd1 vssd1 vccd1 vccd1 _08811_/S sky130_fd_sc_hd__buf_12
XFILLER_113_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07991_ _14756_/Q _07971_/A _07990_/X _08002_/C1 vssd1 vssd1 vccd1 vccd1 _13563_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_140_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_4_7_0_clk clkbuf_4_7_0_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_7_0_clk/X sky130_fd_sc_hd__clkbuf_8
X_09730_ _11710_/A _10132_/B vssd1 vssd1 vccd1 vccd1 _09730_/Y sky130_fd_sc_hd__nor2_8
X_06942_ _06728_/Y _13489_/Q _06730_/Y _13488_/Q _06934_/X vssd1 vssd1 vccd1 vccd1
+ _06943_/B sky130_fd_sc_hd__o221a_1
XFILLER_41_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09661_ _14034_/Q _11883_/A1 _09661_/S vssd1 vssd1 vccd1 vccd1 _14034_/D sky130_fd_sc_hd__mux2_1
XFILLER_67_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06873_ _14514_/Q _06873_/B vssd1 vssd1 vccd1 vccd1 _06873_/Y sky130_fd_sc_hd__nand2_1
XFILLER_55_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08612_ _08722_/A _08612_/B _08612_/C vssd1 vssd1 vccd1 vccd1 _08612_/X sky130_fd_sc_hd__or3_2
XFILLER_94_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09592_ _13968_/Q _11881_/A1 _09594_/S vssd1 vssd1 vccd1 vccd1 _13968_/D sky130_fd_sc_hd__mux2_1
XFILLER_131_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08543_ _14516_/Q _08748_/B1 _08750_/B1 _13642_/Q vssd1 vssd1 vccd1 vccd1 _08543_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_42_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08474_ _13767_/Q _13120_/S _08470_/X _14610_/Q vssd1 vssd1 vccd1 vccd1 _13767_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_24_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07425_ _13331_/A0 _13395_/Q _07481_/S vssd1 vssd1 vccd1 vccd1 _13395_/D sky130_fd_sc_hd__mux2_1
XFILLER_126_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07356_ _07356_/A _07356_/B vssd1 vssd1 vccd1 vccd1 _07356_/Y sky130_fd_sc_hd__nand2_1
XFILLER_164_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07287_ _07287_/A _07287_/B vssd1 vssd1 vccd1 vccd1 _07287_/X sky130_fd_sc_hd__or2_1
XFILLER_163_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09026_ _14073_/Q _09231_/A2 _09403_/B1 _14041_/Q _09532_/A vssd1 vssd1 vccd1 vccd1
+ _09026_/X sky130_fd_sc_hd__a221o_1
XFILLER_164_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09928_ _13110_/B2 _14289_/Q _09930_/S vssd1 vssd1 vccd1 vccd1 _14289_/D sky130_fd_sc_hd__mux2_1
XFILLER_92_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09859_ _14223_/Q _11879_/A1 _09863_/S vssd1 vssd1 vccd1 vccd1 _14223_/D sky130_fd_sc_hd__mux2_1
XFILLER_105_63 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12870_ _14764_/Q _15398_/Q _12871_/S vssd1 vssd1 vccd1 vccd1 _15398_/D sky130_fd_sc_hd__mux2_1
XFILLER_171_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_102 _13444_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11821_ _15243_/Q _11854_/A1 _11850_/S vssd1 vssd1 vccd1 vccd1 _15243_/D sky130_fd_sc_hd__mux2_1
XTAP_2434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_113 input14/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_124 _10192_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1003 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14540_ _15081_/CLK _14540_/D vssd1 vssd1 vccd1 vccd1 _14540_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_42_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11752_ _11860_/A1 _15180_/Q _11774_/S vssd1 vssd1 vccd1 vccd1 _15180_/D sky130_fd_sc_hd__mux2_1
XTAP_1744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_1047 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10703_ _14987_/Q _10733_/A2 _10733_/B1 _14955_/Q _10702_/X vssd1 vssd1 vccd1 vccd1
+ _10703_/X sky130_fd_sc_hd__a221o_2
XTAP_1777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14471_ _15094_/CLK _14471_/D vssd1 vssd1 vccd1 vccd1 _14471_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11683_ _13325_/A0 _15114_/Q _11708_/S vssd1 vssd1 vccd1 vccd1 _15114_/D sky130_fd_sc_hd__mux2_1
XFILLER_14_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13422_ _15379_/CLK _13422_/D vssd1 vssd1 vccd1 vccd1 _13422_/Q sky130_fd_sc_hd__dfxtp_2
X_10634_ _10631_/X _10632_/X _10633_/X _10714_/A2 _15054_/Q vssd1 vssd1 vccd1 vccd1
+ _10634_/X sky130_fd_sc_hd__o32a_4
XFILLER_167_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13353_ _14456_/Q vssd1 vssd1 vccd1 vccd1 _14456_/D sky130_fd_sc_hd__clkbuf_2
X_10565_ _14732_/Q _10735_/S _10564_/Y _14924_/Q vssd1 vssd1 vccd1 vccd1 _14732_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_127_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12304_ _14374_/Q _15190_/Q _13829_/Q _14568_/Q _12541_/S _12544_/A vssd1 vssd1 vccd1
+ vccd1 _12304_/X sky130_fd_sc_hd__mux4_1
XFILLER_6_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_929 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13284_ _14388_/Q _15616_/Q _13284_/S vssd1 vssd1 vccd1 vccd1 _15616_/D sky130_fd_sc_hd__mux2_1
X_10496_ _11536_/B _11500_/A vssd1 vssd1 vccd1 vccd1 _10528_/B sky130_fd_sc_hd__xnor2_1
XFILLER_6_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15023_ _15582_/CLK _15023_/D vssd1 vssd1 vccd1 vccd1 _15023_/Q sky130_fd_sc_hd__dfxtp_1
X_12235_ _14371_/Q _15187_/Q _13826_/Q _14565_/Q _12499_/S _12486_/S1 vssd1 vssd1
+ vccd1 vccd1 _12235_/X sky130_fd_sc_hd__mux4_1
XFILLER_154_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_940 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_962 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12166_ _14368_/Q _15184_/Q _13823_/Q _14562_/Q _12476_/S _12498_/A vssd1 vssd1 vccd1
+ vccd1 _12166_/X sky130_fd_sc_hd__mux4_1
XFILLER_69_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_995 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11117_ _11129_/A _11161_/B _11116_/X vssd1 vssd1 vccd1 vccd1 _11117_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_1_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12097_ _14365_/Q _15181_/Q _13820_/Q _14559_/Q _12472_/S _12465_/S1 vssd1 vssd1
+ vccd1 vccd1 _12097_/X sky130_fd_sc_hd__mux4_1
XFILLER_7_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11048_ _11298_/A _11362_/B vssd1 vssd1 vccd1 vccd1 _11048_/Y sky130_fd_sc_hd__nand2_8
Xinput8 ext_read_data[16] vssd1 vssd1 vccd1 vccd1 input8/X sky130_fd_sc_hd__buf_4
XFILLER_37_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14807_ _15626_/CLK _14807_/D vssd1 vssd1 vccd1 vccd1 _14807_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12999_ _10669_/X _14880_/Q _13029_/S vssd1 vssd1 vccd1 vccd1 _12999_/X sky130_fd_sc_hd__mux2_4
XFILLER_92_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14738_ _15587_/CLK _14738_/D vssd1 vssd1 vccd1 vccd1 _14738_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_44_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14669_ _15606_/CLK _14669_/D vssd1 vssd1 vccd1 vccd1 _14669_/Q sky130_fd_sc_hd__dfxtp_1
X_07210_ _07210_/A vssd1 vssd1 vccd1 vccd1 _07210_/Y sky130_fd_sc_hd__inv_2
X_08190_ _13681_/Q _13319_/A0 _08216_/S vssd1 vssd1 vccd1 vccd1 _13681_/D sky130_fd_sc_hd__mux2_1
XFILLER_146_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07141_ _14834_/Q _07104_/X _07140_/X _07131_/A vssd1 vssd1 vccd1 vccd1 _07141_/X
+ sky130_fd_sc_hd__a22o_4
XFILLER_125_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_1092 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07072_ _14636_/Q _14668_/Q _07078_/S vssd1 vssd1 vccd1 vccd1 _07072_/X sky130_fd_sc_hd__mux2_2
XFILLER_69_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_995 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07974_ _13558_/Q _13557_/Q _07973_/D _13559_/Q vssd1 vssd1 vccd1 vccd1 _07974_/Y
+ sky130_fd_sc_hd__a31oi_1
X_09713_ _13335_/A0 _14083_/Q _09723_/S vssd1 vssd1 vccd1 vccd1 _14083_/D sky130_fd_sc_hd__mux2_1
XFILLER_56_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06925_ _06916_/X _06924_/X _06921_/B vssd1 vssd1 vccd1 vccd1 _06925_/Y sky130_fd_sc_hd__a21oi_1
X_09644_ _14017_/Q _13333_/A0 _09660_/S vssd1 vssd1 vccd1 vccd1 _14017_/D sky130_fd_sc_hd__mux2_1
XFILLER_132_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06856_ _07104_/C _08094_/S vssd1 vssd1 vccd1 vccd1 _07115_/B sky130_fd_sc_hd__nor2_8
XFILLER_167_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09575_ _13951_/Q _11689_/A0 _09589_/S vssd1 vssd1 vccd1 vccd1 _13951_/D sky130_fd_sc_hd__mux2_1
XFILLER_70_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06787_ _08392_/A _06791_/B vssd1 vssd1 vccd1 vccd1 _06789_/B sky130_fd_sc_hd__or2_4
XTAP_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_670 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08526_ _13476_/Q _08746_/A2 _08750_/A2 _13540_/Q _08525_/X vssd1 vssd1 vccd1 vccd1
+ _08526_/X sky130_fd_sc_hd__a221o_1
XFILLER_35_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08457_ _08457_/A _08773_/B vssd1 vssd1 vccd1 vccd1 _08457_/X sky130_fd_sc_hd__and2_1
XFILLER_52_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07408_ _14742_/Q _07407_/X _07480_/S vssd1 vssd1 vccd1 vccd1 _07408_/X sky130_fd_sc_hd__mux2_8
XFILLER_23_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08388_ _08309_/B _11298_/B _11298_/A vssd1 vssd1 vccd1 vccd1 _08388_/X sky130_fd_sc_hd__mux2_2
XFILLER_183_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07339_ _13910_/Q _15497_/Q _07339_/S vssd1 vssd1 vccd1 vccd1 _07339_/X sky130_fd_sc_hd__mux2_8
XFILLER_136_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10350_ _13251_/B vssd1 vssd1 vccd1 vccd1 _10350_/Y sky130_fd_sc_hd__inv_2
XFILLER_125_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09009_ _14523_/Q _14136_/Q _14168_/Q _14104_/Q _09005_/S _09511_/S1 vssd1 vssd1
+ vccd1 vccd1 _09009_/X sky130_fd_sc_hd__mux4_1
XFILLER_151_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10281_ _14666_/Q _14819_/Q _10715_/S vssd1 vssd1 vccd1 vccd1 _14666_/D sky130_fd_sc_hd__mux2_1
XFILLER_2_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12020_ _12595_/A1 _12019_/X _12018_/X _12618_/C1 vssd1 vssd1 vccd1 vccd1 _12021_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_183_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout550 _09047_/S vssd1 vssd1 vccd1 vccd1 _09407_/S sky130_fd_sc_hd__buf_12
XFILLER_120_656 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout561 _09551_/S vssd1 vssd1 vccd1 vccd1 _09557_/S sky130_fd_sc_hd__buf_12
Xfanout572 _14601_/Q vssd1 vssd1 vccd1 vccd1 _08451_/A sky130_fd_sc_hd__buf_12
Xfanout583 _12061_/A vssd1 vssd1 vccd1 vccd1 _11992_/A sky130_fd_sc_hd__buf_6
X_13971_ _14470_/CLK _13971_/D vssd1 vssd1 vccd1 vccd1 _13971_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout594 fanout600/X vssd1 vssd1 vccd1 vccd1 _12563_/A sky130_fd_sc_hd__buf_12
X_12922_ _15450_/Q _15636_/Q _12929_/S vssd1 vssd1 vccd1 vccd1 _15450_/D sky130_fd_sc_hd__mux2_1
XFILLER_18_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15641_ _15641_/CLK _15641_/D vssd1 vssd1 vccd1 vccd1 _15641_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_74_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12853_ _14747_/Q _15381_/Q _12866_/S vssd1 vssd1 vccd1 vccd1 _15381_/D sky130_fd_sc_hd__mux2_1
XTAP_2220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11804_ _15227_/Q _11870_/A1 _11817_/S vssd1 vssd1 vccd1 vccd1 _15227_/D sky130_fd_sc_hd__mux2_1
XTAP_2264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15572_ _15572_/CLK _15572_/D vssd1 vssd1 vccd1 vccd1 _15572_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12784_ _13437_/Q _12647_/B _12737_/A vssd1 vssd1 vccd1 vccd1 _12784_/X sky130_fd_sc_hd__a21o_1
XTAP_2275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14523_ _15081_/CLK _14523_/D vssd1 vssd1 vccd1 vccd1 _14523_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11735_ _15164_/Q _11876_/A1 _11741_/S vssd1 vssd1 vccd1 vccd1 _15164_/D sky130_fd_sc_hd__mux2_1
XTAP_1574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_656 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14454_ _15172_/CLK _14454_/D vssd1 vssd1 vccd1 vccd1 _14454_/Q sky130_fd_sc_hd__dfxtp_1
X_11666_ _13341_/A0 _15098_/Q _11670_/S vssd1 vssd1 vccd1 vccd1 _15098_/D sky130_fd_sc_hd__mux2_1
XFILLER_128_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13405_ _15130_/CLK _13405_/D vssd1 vssd1 vccd1 vccd1 _13405_/Q sky130_fd_sc_hd__dfxtp_1
X_10617_ _15002_/Q _10717_/A2 _10652_/B _13721_/Q _10717_/C1 vssd1 vssd1 vccd1 vccd1
+ _10617_/X sky130_fd_sc_hd__a221o_1
X_14385_ _15666_/CLK _14385_/D vssd1 vssd1 vccd1 vccd1 _14385_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_167_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11597_ _11596_/Y _15068_/Q _11614_/S vssd1 vssd1 vccd1 vccd1 _15068_/D sky130_fd_sc_hd__mux2_1
XFILLER_155_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_183_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13336_ _13336_/A0 _15666_/Q _13350_/S vssd1 vssd1 vccd1 vccd1 _15666_/D sky130_fd_sc_hd__mux2_1
X_10548_ _10548_/A _10548_/B _10548_/C vssd1 vssd1 vccd1 vccd1 _11239_/B sky130_fd_sc_hd__and3_1
XFILLER_143_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13267_ _15351_/Q _15598_/Q _13300_/S vssd1 vssd1 vccd1 vccd1 _15598_/D sky130_fd_sc_hd__mux2_1
X_10479_ _10520_/A1 _13789_/Q _13757_/Q _10520_/B2 vssd1 vssd1 vccd1 vccd1 _10479_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_142_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15006_ _15006_/CLK _15006_/D vssd1 vssd1 vccd1 vccd1 _15006_/Q sky130_fd_sc_hd__dfxtp_1
X_12218_ _12498_/A _12218_/B vssd1 vssd1 vccd1 vccd1 _12218_/X sky130_fd_sc_hd__and2_1
XFILLER_29_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13198_ _15567_/Q _13214_/B vssd1 vssd1 vccd1 vccd1 _13198_/X sky130_fd_sc_hd__and2_1
XFILLER_155_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12149_ _12268_/A _12149_/B vssd1 vssd1 vccd1 vccd1 _12149_/X sky130_fd_sc_hd__and2_1
XFILLER_111_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06710_ _14507_/Q vssd1 vssd1 vccd1 vccd1 _06710_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07690_ _13485_/Q _07717_/A vssd1 vssd1 vccd1 vccd1 _07691_/B sky130_fd_sc_hd__xnor2_1
XFILLER_92_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_467 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09360_ _13961_/Q _13703_/Q _09521_/S vssd1 vssd1 vccd1 vccd1 _09360_/X sky130_fd_sc_hd__mux2_1
XFILLER_80_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08311_ _08244_/A _13766_/Q _15406_/Q _08244_/B vssd1 vssd1 vccd1 vccd1 _08311_/X
+ sky130_fd_sc_hd__a22o_2
XFILLER_177_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09291_ _08510_/B _09287_/X _09290_/X _09286_/X vssd1 vssd1 vccd1 vccd1 _09291_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_178_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_13 _10734_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08242_ _13774_/Q _08237_/A _07331_/A _10457_/A2 _08240_/X vssd1 vssd1 vccd1 vccd1
+ _08242_/X sky130_fd_sc_hd__a221o_2
XANTENNA_24 _15418_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_35 _14743_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_46 input24/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_57 _07165_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08173_ _08133_/S input18/X _08185_/A vssd1 vssd1 vccd1 vccd1 _08173_/X sky130_fd_sc_hd__and3b_1
XANTENNA_68 _07133_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_79 _07110_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07124_ _14842_/Q _14834_/Q _08094_/S vssd1 vssd1 vccd1 vccd1 _07125_/B sky130_fd_sc_hd__mux2_1
XFILLER_180_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07055_ _07054_/X _13597_/Q _12764_/S vssd1 vssd1 vccd1 vccd1 _07055_/X sky130_fd_sc_hd__mux2_1
XFILLER_133_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_910 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07957_ _14747_/Q _07964_/A _07956_/X _07965_/C1 vssd1 vssd1 vccd1 vccd1 _13554_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_96_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06908_ _15382_/Q _07595_/B _15381_/Q _06727_/Y _06894_/X vssd1 vssd1 vccd1 vccd1
+ _06908_/X sky130_fd_sc_hd__a221o_1
X_07888_ _14761_/Q _07903_/A _07887_/Y _08012_/C1 vssd1 vssd1 vccd1 vccd1 _13536_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_56_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09627_ _14001_/Q _11816_/A1 _09627_/S vssd1 vssd1 vccd1 vccd1 _14001_/D sky130_fd_sc_hd__mux2_1
XFILLER_56_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06839_ _08668_/C _14905_/Q _06837_/X _06838_/X vssd1 vssd1 vccd1 vccd1 _06839_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_43_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xcore_649 vssd1 vssd1 vccd1 vccd1 core_649/HI ext_address[1] sky130_fd_sc_hd__conb_1
X_09558_ _15139_/Q _09558_/A2 _13130_/C1 _09557_/X vssd1 vssd1 vccd1 vccd1 _09558_/X
+ sky130_fd_sc_hd__a22o_1
X_08509_ _08668_/D _08512_/B vssd1 vssd1 vccd1 vccd1 _08769_/B sky130_fd_sc_hd__nand2_1
XFILLER_12_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09489_ _15104_/Q _08497_/A _09519_/B1 _08501_/A vssd1 vssd1 vccd1 vccd1 _09489_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_52_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11520_ _11521_/A _11521_/B vssd1 vssd1 vccd1 vccd1 _11531_/A sky130_fd_sc_hd__nand2_1
XFILLER_62_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11451_ _11440_/A _11440_/B _11443_/Y vssd1 vssd1 vccd1 vccd1 _11452_/B sky130_fd_sc_hd__a21oi_1
X_10402_ _13171_/B _11414_/D vssd1 vssd1 vccd1 vccd1 _10410_/A sky130_fd_sc_hd__or2_1
XFILLER_183_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14170_ _15212_/CLK _14170_/D vssd1 vssd1 vccd1 vccd1 _14170_/Q sky130_fd_sc_hd__dfxtp_1
X_11382_ _11384_/A vssd1 vssd1 vccd1 vccd1 _11382_/Y sky130_fd_sc_hd__inv_2
XFILLER_180_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13121_ _15530_/Q _10871_/S _08402_/X vssd1 vssd1 vccd1 vccd1 _15530_/D sky130_fd_sc_hd__o21a_1
XFILLER_164_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10333_ _14718_/Q _14911_/Q _10343_/S vssd1 vssd1 vccd1 vccd1 _14718_/D sky130_fd_sc_hd__mux2_1
XFILLER_139_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13052_ _12937_/X _13104_/A2 _13104_/B1 _07376_/X vssd1 vssd1 vccd1 vccd1 _13052_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_152_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10264_ _14649_/Q _14802_/Q _10615_/S vssd1 vssd1 vccd1 vccd1 _14649_/D sky130_fd_sc_hd__mux2_1
X_12003_ _15113_/Q _15081_/Q _15654_/Q _13388_/Q _12407_/S _12590_/A vssd1 vssd1 vccd1
+ vccd1 _12003_/X sky130_fd_sc_hd__mux4_1
X_10195_ _11881_/A1 _14579_/Q _10197_/S vssd1 vssd1 vccd1 vccd1 _14579_/D sky130_fd_sc_hd__mux2_1
Xfanout380 _11349_/A vssd1 vssd1 vccd1 vccd1 _11088_/S sky130_fd_sc_hd__buf_12
XFILLER_16_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout391 _08231_/X vssd1 vssd1 vccd1 vccd1 _11380_/A sky130_fd_sc_hd__buf_12
XFILLER_93_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13954_ _15497_/CLK _13954_/D vssd1 vssd1 vccd1 vccd1 _13954_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12905_ _15433_/Q _15619_/Q _12932_/S vssd1 vssd1 vccd1 vccd1 _15433_/D sky130_fd_sc_hd__mux2_1
XFILLER_35_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_194_clk clkbuf_5_20_0_clk/X vssd1 vssd1 vccd1 vccd1 _15127_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_19_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13885_ _14415_/CLK _13885_/D vssd1 vssd1 vccd1 vccd1 _13885_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_74_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15624_ _15624_/CLK _15624_/D vssd1 vssd1 vccd1 vccd1 _15624_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12836_ _13611_/Q _12647_/B _06863_/B vssd1 vssd1 vccd1 vccd1 _12836_/X sky130_fd_sc_hd__o21a_1
XTAP_2061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15555_ _15556_/CLK _15555_/D vssd1 vssd1 vccd1 vccd1 _15555_/Q sky130_fd_sc_hd__dfxtp_1
X_12767_ _15358_/Q _15357_/Q _12767_/C vssd1 vssd1 vccd1 vccd1 _12776_/B sky130_fd_sc_hd__and3_1
XTAP_1360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14506_ _14506_/CLK _14506_/D vssd1 vssd1 vccd1 vccd1 _14506_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_148_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11718_ _15147_/Q _12967_/A1 _11741_/S vssd1 vssd1 vccd1 vccd1 _15147_/D sky130_fd_sc_hd__mux2_1
X_15486_ _15536_/CLK _15486_/D vssd1 vssd1 vccd1 vccd1 _15486_/Q sky130_fd_sc_hd__dfxtp_1
X_12698_ _13425_/Q _12697_/X _12728_/S vssd1 vssd1 vccd1 vccd1 _12699_/B sky130_fd_sc_hd__mux2_1
XFILLER_174_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14437_ _15332_/CLK _14437_/D vssd1 vssd1 vccd1 vccd1 _14437_/Q sky130_fd_sc_hd__dfxtp_1
Xinput11 ext_read_data[19] vssd1 vssd1 vccd1 vccd1 input11/X sky130_fd_sc_hd__buf_4
X_11649_ _11649_/A0 _15081_/Q _11675_/S vssd1 vssd1 vccd1 vccd1 _15081_/D sky130_fd_sc_hd__mux2_1
Xinput22 ext_read_data[29] vssd1 vssd1 vccd1 vccd1 input22/X sky130_fd_sc_hd__buf_6
Xinput33 ext_ready vssd1 vssd1 vccd1 vccd1 input33/X sky130_fd_sc_hd__buf_4
XFILLER_162_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14368_ _15184_/CLK _14368_/D vssd1 vssd1 vccd1 vccd1 _14368_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_183_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_1103 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13319_ _13319_/A0 _15649_/Q _13345_/S vssd1 vssd1 vccd1 vccd1 _15649_/D sky130_fd_sc_hd__mux2_1
XFILLER_115_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14299_ _15660_/CLK _14299_/D vssd1 vssd1 vccd1 vccd1 _14299_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_171_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08860_ _13881_/Q _11858_/A1 _08885_/S vssd1 vssd1 vccd1 vccd1 _13881_/D sky130_fd_sc_hd__mux2_1
XFILLER_69_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07811_ _07816_/A _07811_/B vssd1 vssd1 vccd1 vccd1 _07811_/Y sky130_fd_sc_hd__nand2_1
XFILLER_57_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08791_ _11858_/A1 _13817_/Q _08811_/S vssd1 vssd1 vccd1 vccd1 _13817_/D sky130_fd_sc_hd__mux2_1
XFILLER_96_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07742_ _13499_/Q _07746_/C vssd1 vssd1 vccd1 vccd1 _07743_/B sky130_fd_sc_hd__xnor2_1
XFILLER_38_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07673_ _07671_/Y _07679_/C _07676_/A vssd1 vssd1 vccd1 vccd1 _07673_/Y sky130_fd_sc_hd__o21ai_1
Xclkbuf_leaf_185_clk clkbuf_5_21_0_clk/X vssd1 vssd1 vccd1 vccd1 _14482_/CLK sky130_fd_sc_hd__clkbuf_16
X_09412_ _13931_/Q _13119_/S _09411_/X vssd1 vssd1 vccd1 vccd1 _13931_/D sky130_fd_sc_hd__a21o_1
X_09343_ _15129_/Q _09536_/A2 _13130_/C1 _09342_/X vssd1 vssd1 vccd1 vccd1 _09343_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_21_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09274_ _09550_/A1 _09272_/X _09273_/X vssd1 vssd1 vccd1 vccd1 _09275_/C sky130_fd_sc_hd__a21o_1
XFILLER_166_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08225_ _08237_/A _08240_/A vssd1 vssd1 vccd1 vccd1 _08225_/Y sky130_fd_sc_hd__nor2_8
XFILLER_165_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08156_ _13665_/Q _10285_/S _08154_/X _08155_/X vssd1 vssd1 vccd1 vccd1 _13665_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_162_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07107_ _14900_/Q _08151_/S _07163_/A _07103_/B _08121_/B vssd1 vssd1 vccd1 vccd1
+ _07107_/X sky130_fd_sc_hd__o2111a_4
XFILLER_180_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08087_ _06825_/C _08083_/A _08086_/Y input35/X vssd1 vssd1 vccd1 vccd1 _08087_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_164_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07038_ _07037_/X _14745_/Q _07077_/S vssd1 vssd1 vccd1 vccd1 _13591_/D sky130_fd_sc_hd__mux2_1
XFILLER_79_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08989_ _15112_/Q _09536_/A2 _13130_/B1 _15080_/Q _08988_/X vssd1 vssd1 vccd1 vccd1
+ _08989_/X sky130_fd_sc_hd__a221o_1
XFILLER_57_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10951_ _13252_/A _10951_/B vssd1 vssd1 vccd1 vccd1 _10951_/Y sky130_fd_sc_hd__nand2_1
XFILLER_16_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_176_clk clkbuf_5_23_0_clk/X vssd1 vssd1 vccd1 vccd1 _15326_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_17_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13670_ _15645_/CLK _13670_/D vssd1 vssd1 vccd1 vccd1 _13670_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10882_ _14914_/Q _15545_/Q _13134_/A vssd1 vssd1 vccd1 vccd1 _14914_/D sky130_fd_sc_hd__mux2_1
X_12621_ _12622_/A _15615_/D vssd1 vssd1 vccd1 vccd1 _12621_/Y sky130_fd_sc_hd__nor2_4
XFILLER_188_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15340_ _15620_/CLK _15340_/D vssd1 vssd1 vccd1 vccd1 _15340_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_19_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12552_ _14257_/Q _14289_/Q _14321_/Q _14353_/Q _12430_/S _12567_/A vssd1 vssd1 vccd1
+ vccd1 _12552_/X sky130_fd_sc_hd__mux4_1
XFILLER_184_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11503_ _11505_/C _11505_/D vssd1 vssd1 vccd1 vccd1 _11503_/X sky130_fd_sc_hd__and2_1
X_15271_ _15303_/CLK _15271_/D vssd1 vssd1 vccd1 vccd1 _15271_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_157_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12483_ _14254_/Q _14286_/Q _14318_/Q _14350_/Q _12489_/S0 _12489_/S1 vssd1 vssd1
+ vccd1 vccd1 _12483_/X sky130_fd_sc_hd__mux4_1
Xclkbuf_1_0_0_clk clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 clkbuf_1_0_1_clk/A sky130_fd_sc_hd__clkbuf_8
XFILLER_7_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14222_ _15556_/CLK _14222_/D vssd1 vssd1 vccd1 vccd1 _14222_/Q sky130_fd_sc_hd__dfxtp_1
X_11434_ _11460_/B _11441_/B vssd1 vssd1 vccd1 vccd1 _11434_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_144_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14153_ _15679_/CLK _14153_/D vssd1 vssd1 vccd1 vccd1 _14153_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_100_clk _15447_/CLK vssd1 vssd1 vccd1 vccd1 _15375_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_138_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11365_ _11363_/X _11365_/B vssd1 vssd1 vccd1 vccd1 _11368_/A sky130_fd_sc_hd__and2b_1
XFILLER_164_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13104_ _13023_/X _13104_/A2 _13104_/B1 _13104_/B2 vssd1 vssd1 vccd1 vccd1 _13104_/X
+ sky130_fd_sc_hd__a22o_1
X_10316_ _14701_/Q _14886_/Q _10695_/S vssd1 vssd1 vccd1 vccd1 _14701_/D sky130_fd_sc_hd__mux2_1
XFILLER_4_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14084_ _15651_/CLK _14084_/D vssd1 vssd1 vccd1 vccd1 _14084_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_112_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11296_ _11296_/A vssd1 vssd1 vccd1 vccd1 _11296_/Y sky130_fd_sc_hd__inv_2
XTAP_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13035_ _10729_/X _14892_/Q _13038_/S vssd1 vssd1 vccd1 vccd1 _13035_/X sky130_fd_sc_hd__mux2_4
X_10247_ _14632_/Q _14785_/Q _10630_/S vssd1 vssd1 vccd1 vccd1 _14632_/D sky130_fd_sc_hd__mux2_1
XFILLER_152_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10178_ _13331_/A0 _14562_/Q _10192_/S vssd1 vssd1 vccd1 vccd1 _14562_/D sky130_fd_sc_hd__mux2_1
XFILLER_94_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14986_ _14988_/CLK _14986_/D vssd1 vssd1 vccd1 vccd1 _14986_/Q sky130_fd_sc_hd__dfxtp_1
X_13937_ _15673_/CLK _13937_/D vssd1 vssd1 vccd1 vccd1 _13937_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_167_clk clkbuf_5_22_0_clk/X vssd1 vssd1 vccd1 vccd1 _15552_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_62_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13868_ _15662_/CLK _13868_/D vssd1 vssd1 vccd1 vccd1 _13868_/Q sky130_fd_sc_hd__dfxtp_1
X_15607_ _15607_/CLK _15607_/D vssd1 vssd1 vccd1 vccd1 _15607_/Q sky130_fd_sc_hd__dfxtp_1
X_12819_ _15365_/Q _12819_/B vssd1 vssd1 vccd1 vccd1 _12820_/B sky130_fd_sc_hd__nor2_1
X_13799_ _15461_/CLK _13799_/D vssd1 vssd1 vccd1 vccd1 _13799_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_43_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15538_ _15617_/CLK _15538_/D vssd1 vssd1 vccd1 vccd1 _15538_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_187_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_935 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15469_ _15501_/CLK _15469_/D vssd1 vssd1 vccd1 vccd1 _15469_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_176_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_495 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08010_ _13569_/Q _08017_/D vssd1 vssd1 vccd1 vccd1 _08011_/B sky130_fd_sc_hd__xnor2_1
XFILLER_147_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09961_ _13110_/B2 _14321_/Q _09963_/S vssd1 vssd1 vccd1 vccd1 _14321_/D sky130_fd_sc_hd__mux2_1
XFILLER_116_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08912_ _14455_/Q _09536_/A2 _08540_/B _14423_/Q _08911_/X vssd1 vssd1 vccd1 vccd1
+ _08912_/X sky130_fd_sc_hd__a221o_1
XFILLER_98_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09892_ _13345_/A0 _14254_/Q _09892_/S vssd1 vssd1 vccd1 vccd1 _14254_/D sky130_fd_sc_hd__mux2_1
XTAP_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08843_ _13866_/Q _13098_/B2 _08851_/S vssd1 vssd1 vccd1 vccd1 _13866_/D sky130_fd_sc_hd__mux2_1
XTAP_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08774_ _06796_/B _08477_/C _08772_/X _08773_/Y vssd1 vssd1 vccd1 vccd1 _08774_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_38_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07725_ _07723_/Y _07727_/B _07750_/A vssd1 vssd1 vccd1 vccd1 _07725_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_26_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_158_clk clkbuf_5_19_0_clk/X vssd1 vssd1 vccd1 vccd1 _15648_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_81_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07656_ _07653_/Y _07665_/C _07644_/A vssd1 vssd1 vccd1 vccd1 _07656_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_129_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07587_ _13458_/Q _07587_/B vssd1 vssd1 vccd1 vccd1 _07587_/Y sky130_fd_sc_hd__nor2_1
XFILLER_179_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_902 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09326_ _09466_/A _09326_/B vssd1 vssd1 vccd1 vccd1 _09326_/X sky130_fd_sc_hd__or2_1
XFILLER_40_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09257_ _08510_/B _09253_/X _09256_/X vssd1 vssd1 vccd1 vccd1 _09257_/X sky130_fd_sc_hd__a21o_1
XFILLER_167_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08208_ _13699_/Q _13337_/A0 _08221_/S vssd1 vssd1 vccd1 vccd1 _13699_/D sky130_fd_sc_hd__mux2_1
XFILLER_126_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09188_ _14081_/Q _09231_/A2 _09403_/B1 _14049_/Q _09221_/A vssd1 vssd1 vccd1 vccd1
+ _09188_/X sky130_fd_sc_hd__a221o_1
X_08139_ _08151_/S _08137_/X _08138_/Y _08121_/X vssd1 vssd1 vccd1 vccd1 _08139_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_134_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11150_ _11129_/A _11096_/B _11129_/Y vssd1 vssd1 vccd1 vccd1 _11195_/B sky130_fd_sc_hd__a21oi_1
XFILLER_175_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10101_ _14487_/Q _14735_/Q _10131_/S vssd1 vssd1 vccd1 vccd1 _14487_/D sky130_fd_sc_hd__mux2_1
XFILLER_108_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_96 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11081_ _10350_/Y _11363_/B _11080_/X _11362_/B vssd1 vssd1 vccd1 vccd1 _11082_/A
+ sky130_fd_sc_hd__o22ai_4
XFILLER_103_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10032_ _10032_/A _11818_/A vssd1 vssd1 vccd1 vccd1 _10032_/Y sky130_fd_sc_hd__nor2_8
XFILLER_103_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14840_ _15507_/CLK _14840_/D vssd1 vssd1 vccd1 vccd1 _14840_/Q sky130_fd_sc_hd__dfxtp_1
X_14771_ _15588_/CLK _14771_/D vssd1 vssd1 vccd1 vccd1 _14771_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_112_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11983_ _15277_/Q _15245_/Q _15213_/Q _15144_/Q _12154_/S _12253_/S1 vssd1 vssd1
+ vccd1 vccd1 _11984_/B sky130_fd_sc_hd__mux4_1
XFILLER_17_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_149_clk clkbuf_5_25_0_clk/X vssd1 vssd1 vccd1 vccd1 _15615_/CLK sky130_fd_sc_hd__clkbuf_16
X_13722_ _15006_/CLK _13722_/D vssd1 vssd1 vccd1 vccd1 _13722_/Q sky130_fd_sc_hd__dfxtp_1
X_10934_ _11569_/B _10948_/B vssd1 vssd1 vccd1 vccd1 _10934_/Y sky130_fd_sc_hd__nand2_1
XFILLER_56_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_351 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13653_ _14892_/CLK _13653_/D vssd1 vssd1 vccd1 vccd1 _13653_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10865_ _14897_/Q _15534_/Q _12904_/S vssd1 vssd1 vccd1 vccd1 _14897_/D sky130_fd_sc_hd__mux2_1
X_12604_ _15304_/Q _15272_/Q _15240_/Q _15171_/Q _12518_/S _12613_/A vssd1 vssd1 vccd1
+ vccd1 _12605_/B sky130_fd_sc_hd__mux4_1
XPHY_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_250 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13584_ _15620_/CLK _13584_/D vssd1 vssd1 vccd1 vccd1 _13584_/Q sky130_fd_sc_hd__dfxtp_2
X_10796_ _14828_/Q _15460_/Q _12932_/S vssd1 vssd1 vccd1 vccd1 _14828_/D sky130_fd_sc_hd__mux2_1
XPHY_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15323_ _15666_/CLK _15323_/D vssd1 vssd1 vccd1 vccd1 _15323_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_158_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12535_ _15301_/Q _15269_/Q _15237_/Q _15168_/Q _12612_/S _12613_/A vssd1 vssd1 vccd1
+ vccd1 _12536_/B sky130_fd_sc_hd__mux4_1
XFILLER_185_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_927 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15254_ _15286_/CLK _15254_/D vssd1 vssd1 vccd1 vccd1 _15254_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_92 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12466_ _15298_/Q _15266_/Q _15234_/Q _15165_/Q _12489_/S0 _12489_/S1 vssd1 vssd1
+ vccd1 vccd1 _12467_/B sky130_fd_sc_hd__mux4_1
XFILLER_173_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_1062 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14205_ _15181_/CLK _14205_/D vssd1 vssd1 vccd1 vccd1 _14205_/Q sky130_fd_sc_hd__dfxtp_1
X_11417_ _11419_/A _11419_/B vssd1 vssd1 vccd1 vccd1 _11420_/A sky130_fd_sc_hd__or2_1
X_15185_ _15218_/CLK _15185_/D vssd1 vssd1 vccd1 vccd1 _15185_/Q sky130_fd_sc_hd__dfxtp_1
X_12397_ _15295_/Q _15263_/Q _15231_/Q _15162_/Q _12591_/S _12590_/A vssd1 vssd1 vccd1
+ vccd1 _12398_/B sky130_fd_sc_hd__mux4_1
XFILLER_153_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14136_ _15081_/CLK _14136_/D vssd1 vssd1 vccd1 vccd1 _14136_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_126_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11348_ _11007_/B _11013_/X _11259_/S vssd1 vssd1 vccd1 vccd1 _11348_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_4_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14067_ _14470_/CLK _14067_/D vssd1 vssd1 vccd1 vccd1 _14067_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11279_ _11025_/A _13217_/B _11027_/A vssd1 vssd1 vccd1 vccd1 _11280_/B sky130_fd_sc_hd__o21ai_1
X_13018_ _13343_/A0 _13024_/A2 _13017_/X _13024_/B2 vssd1 vssd1 vccd1 vccd1 _13018_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_39_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14969_ _15584_/CLK _14969_/D vssd1 vssd1 vccd1 vccd1 _14969_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07510_ _14740_/Q _13419_/Q _07535_/S vssd1 vssd1 vccd1 vccd1 _13419_/D sky130_fd_sc_hd__mux2_1
X_08490_ _08490_/A1 _08421_/Y _08465_/X hold5/A vssd1 vssd1 vccd1 vccd1 _08490_/X
+ sky130_fd_sc_hd__a22o_1
X_07441_ _13335_/A0 _13399_/Q _07481_/S vssd1 vssd1 vccd1 vccd1 _13399_/D sky130_fd_sc_hd__mux2_1
X_07372_ _07482_/C _07474_/B vssd1 vssd1 vccd1 vccd1 _07372_/X sky130_fd_sc_hd__and2b_2
X_09111_ _15118_/Q _15086_/Q _15659_/Q _13393_/Q _09190_/S _09429_/S1 vssd1 vssd1
+ vccd1 vccd1 _09111_/X sky130_fd_sc_hd__mux4_1
XFILLER_31_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09042_ _14235_/Q _14267_/Q _14299_/Q _14331_/Q _09225_/S0 _09225_/S1 vssd1 vssd1
+ vccd1 vccd1 _09042_/X sky130_fd_sc_hd__mux4_2
XFILLER_108_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_5_16_0_clk clkbuf_4_8_0_clk/X vssd1 vssd1 vccd1 vccd1 clkbuf_5_16_0_clk/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_131_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09944_ _13331_/A0 _14304_/Q _09958_/S vssd1 vssd1 vccd1 vccd1 _14304_/D sky130_fd_sc_hd__mux2_1
XFILLER_86_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09875_ _11861_/A1 _14237_/Q _09892_/S vssd1 vssd1 vccd1 vccd1 _14237_/D sky130_fd_sc_hd__mux2_1
XFILLER_112_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08826_ _13849_/Q _11858_/A1 _08846_/S vssd1 vssd1 vccd1 vccd1 _13849_/D sky130_fd_sc_hd__mux2_1
XFILLER_57_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_178 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08757_ _08421_/A _08777_/B _08755_/X vssd1 vssd1 vccd1 vccd1 _08757_/Y sky130_fd_sc_hd__o21ai_1
XTAP_2605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07708_ _13489_/Q _07732_/A _13490_/Q vssd1 vssd1 vccd1 vccd1 _07708_/Y sky130_fd_sc_hd__a21oi_1
XTAP_2638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08688_ _10765_/S _08688_/B _08688_/C vssd1 vssd1 vccd1 vccd1 _08688_/X sky130_fd_sc_hd__or3_4
XFILLER_54_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07639_ _13472_/Q _13471_/Q _13470_/Q _13469_/Q vssd1 vssd1 vccd1 vccd1 _07655_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_41_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10650_ _14748_/Q _10649_/X _10650_/S vssd1 vssd1 vccd1 vccd1 _14748_/D sky130_fd_sc_hd__mux2_1
XFILLER_110_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09309_ _14474_/Q _14442_/Q _13863_/Q _14216_/Q _09481_/S _09553_/A1 vssd1 vssd1
+ vccd1 vccd1 _09309_/X sky130_fd_sc_hd__mux4_1
XFILLER_166_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_1095 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10581_ _10581_/A _10581_/B _14927_/Q vssd1 vssd1 vccd1 vccd1 _10581_/X sky130_fd_sc_hd__and3_1
XFILLER_70_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12320_ _12320_/A _12320_/B _12320_/C vssd1 vssd1 vccd1 vccd1 _12320_/X sky130_fd_sc_hd__and3_1
XFILLER_142_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12251_ _12504_/A _12251_/B _12251_/C vssd1 vssd1 vccd1 vccd1 _12251_/X sky130_fd_sc_hd__and3_1
XFILLER_5_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11202_ _11202_/A _11389_/B _11389_/C vssd1 vssd1 vccd1 vccd1 _11202_/X sky130_fd_sc_hd__and3_1
XFILLER_135_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12182_ _12596_/A _12182_/B _12182_/C vssd1 vssd1 vccd1 vccd1 _12182_/X sky130_fd_sc_hd__and3_1
XFILLER_79_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11133_ _11344_/A _11132_/X _11202_/A vssd1 vssd1 vccd1 vccd1 _11133_/X sky130_fd_sc_hd__o21a_1
XFILLER_134_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11064_ _11414_/A _11175_/B vssd1 vssd1 vccd1 vccd1 _11064_/Y sky130_fd_sc_hd__nor2_1
XFILLER_76_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10015_ _11761_/A0 _14373_/Q _10029_/S vssd1 vssd1 vccd1 vccd1 _14373_/D sky130_fd_sc_hd__mux2_1
XFILLER_49_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14823_ _15606_/CLK _14823_/D vssd1 vssd1 vccd1 vccd1 _14823_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_28_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14754_ _15452_/CLK _14754_/D vssd1 vssd1 vccd1 vccd1 _14754_/Q sky130_fd_sc_hd__dfxtp_4
X_11966_ _13878_/Q _14393_/Q _12079_/S vssd1 vssd1 vccd1 vccd1 _11966_/X sky130_fd_sc_hd__mux2_1
XFILLER_44_340 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10917_ _14941_/Q _10944_/B _10916_/Y _13189_/B vssd1 vssd1 vccd1 vccd1 _14941_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_17_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13705_ _14542_/CLK _13705_/D vssd1 vssd1 vccd1 vccd1 _13705_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14685_ _15607_/CLK _14685_/D vssd1 vssd1 vccd1 vccd1 _14685_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11897_ _13875_/Q _14390_/Q _12269_/S vssd1 vssd1 vccd1 vccd1 _11897_/X sky130_fd_sc_hd__mux2_1
X_13636_ _14510_/CLK _13636_/D vssd1 vssd1 vccd1 vccd1 _13636_/Q sky130_fd_sc_hd__dfxtp_1
X_10848_ _14880_/Q _13788_/Q _12929_/S vssd1 vssd1 vccd1 vccd1 _14880_/D sky130_fd_sc_hd__mux2_1
XFILLER_32_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13567_ _14511_/CLK _13567_/D vssd1 vssd1 vccd1 vccd1 _13567_/Q sky130_fd_sc_hd__dfxtp_2
X_10779_ _14811_/Q _15443_/Q _12918_/S vssd1 vssd1 vccd1 vccd1 _14811_/D sky130_fd_sc_hd__mux2_1
X_12518_ _13902_/Q _14417_/Q _12518_/S vssd1 vssd1 vccd1 vccd1 _12518_/X sky130_fd_sc_hd__mux2_1
X_15306_ _15306_/CLK _15306_/D vssd1 vssd1 vccd1 vccd1 _15306_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_173_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13498_ _13565_/CLK _13498_/D vssd1 vssd1 vccd1 vccd1 _13498_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_157_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15237_ _15326_/CLK _15237_/D vssd1 vssd1 vccd1 vccd1 _15237_/Q sky130_fd_sc_hd__dfxtp_1
X_12449_ _13899_/Q _14414_/Q _12453_/S vssd1 vssd1 vccd1 vccd1 _12449_/X sky130_fd_sc_hd__mux2_1
XFILLER_126_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_172_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15168_ _15326_/CLK _15168_/D vssd1 vssd1 vccd1 vccd1 _15168_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_992 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14119_ _15096_/CLK _14119_/D vssd1 vssd1 vccd1 vccd1 _14119_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07990_ _07992_/B _07989_/X _07971_/A vssd1 vssd1 vccd1 vccd1 _07990_/X sky130_fd_sc_hd__a21bo_1
Xfanout209 _09629_/Y vssd1 vssd1 vccd1 vccd1 _09660_/S sky130_fd_sc_hd__buf_12
X_15099_ _15328_/CLK _15099_/D vssd1 vssd1 vccd1 vccd1 _15099_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_141_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06941_ _06941_/A _06941_/B _06941_/C vssd1 vssd1 vccd1 vccd1 _06944_/C sky130_fd_sc_hd__nand3_2
XFILLER_68_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09660_ _14033_/Q _11816_/A1 _09660_/S vssd1 vssd1 vccd1 vccd1 _14033_/D sky130_fd_sc_hd__mux2_1
XFILLER_95_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06872_ _06872_/A _13508_/Q vssd1 vssd1 vccd1 vccd1 _06879_/B sky130_fd_sc_hd__or2_1
XFILLER_39_156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08611_ _14506_/Q _08748_/B1 _08609_/X _08610_/X vssd1 vssd1 vccd1 vccd1 _08612_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_95_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09591_ _13967_/Q _11847_/A1 _09594_/S vssd1 vssd1 vccd1 vccd1 _13967_/D sky130_fd_sc_hd__mux2_1
XFILLER_83_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08542_ _13475_/Q _08746_/A2 _08750_/A2 _13539_/Q _08541_/X vssd1 vssd1 vccd1 vccd1
+ _08542_/X sky130_fd_sc_hd__a221o_1
XFILLER_39_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08473_ _13766_/Q _10764_/S _08470_/X _14611_/Q vssd1 vssd1 vccd1 vccd1 _13766_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_50_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_518 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07424_ _14746_/Q _07423_/X _07480_/S vssd1 vssd1 vccd1 vccd1 _07424_/X sky130_fd_sc_hd__mux2_8
XFILLER_51_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07355_ _07355_/A _07355_/B vssd1 vssd1 vccd1 vccd1 _07355_/X sky130_fd_sc_hd__or2_1
XFILLER_148_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07286_ _07280_/Y _07281_/X _07287_/A _07287_/B vssd1 vssd1 vccd1 vccd1 _07348_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_164_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09025_ _14009_/Q _13977_/Q _09521_/S vssd1 vssd1 vccd1 vccd1 _09025_/X sky130_fd_sc_hd__mux2_1
XFILLER_40_49 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_1088 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09927_ _11847_/A1 _14288_/Q _09930_/S vssd1 vssd1 vccd1 vccd1 _14288_/D sky130_fd_sc_hd__mux2_1
XFILLER_77_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09858_ _14222_/Q _13345_/A0 _09858_/S vssd1 vssd1 vccd1 vccd1 _14222_/D sky130_fd_sc_hd__mux2_1
XTAP_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08809_ _11876_/A1 _13835_/Q _08811_/S vssd1 vssd1 vccd1 vccd1 _13835_/D sky130_fd_sc_hd__mux2_1
XTAP_3136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09789_ _14156_/Q _11877_/A1 _09790_/S vssd1 vssd1 vccd1 vccd1 _14156_/D sky130_fd_sc_hd__mux2_1
XTAP_3147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_103 _13789_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11820_ _15242_/Q _13320_/A0 _11850_/S vssd1 vssd1 vccd1 vccd1 _15242_/D sky130_fd_sc_hd__mux2_1
XTAP_3169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_114 input16/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_125 _09435_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11751_ _12967_/A1 _15179_/Q _11774_/S vssd1 vssd1 vccd1 vccd1 _15179_/D sky130_fd_sc_hd__mux2_1
XFILLER_14_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1015 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_80_clk clkbuf_5_15_0_clk/X vssd1 vssd1 vccd1 vccd1 _14774_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_1756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10702_ _15019_/Q _10717_/A2 _10652_/B _15036_/Q _10717_/C1 vssd1 vssd1 vccd1 vccd1
+ _10702_/X sky130_fd_sc_hd__a221o_1
XTAP_1767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14470_ _14470_/CLK _14470_/D vssd1 vssd1 vccd1 vccd1 _14470_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11682_ _13324_/A0 _15113_/Q _11708_/S vssd1 vssd1 vccd1 vccd1 _15113_/D sky130_fd_sc_hd__mux2_1
XTAP_1789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13421_ _15375_/CLK _13421_/D vssd1 vssd1 vccd1 vccd1 _13421_/Q sky130_fd_sc_hd__dfxtp_1
X_10633_ _15564_/Q _10706_/B _10718_/A2 _14973_/Q vssd1 vssd1 vccd1 vccd1 _10633_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_14_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13352_ _14455_/Q vssd1 vssd1 vccd1 vccd1 _14455_/D sky130_fd_sc_hd__clkbuf_2
X_10564_ _10564_/A vssd1 vssd1 vccd1 vccd1 _10564_/Y sky130_fd_sc_hd__inv_2
XFILLER_155_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12303_ _12299_/X _12300_/X _12617_/S vssd1 vssd1 vccd1 vccd1 _12303_/X sky130_fd_sc_hd__mux2_1
XFILLER_108_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13283_ _15367_/Q _15614_/Q _13291_/S vssd1 vssd1 vccd1 vccd1 _15614_/D sky130_fd_sc_hd__mux2_1
X_10495_ _07258_/A _10523_/A2 _10494_/X vssd1 vssd1 vccd1 vccd1 _11500_/A sky130_fd_sc_hd__a21o_4
X_15022_ _15041_/CLK _15022_/D vssd1 vssd1 vccd1 vccd1 _15022_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_142_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12234_ _12230_/X _12231_/X _12502_/S vssd1 vssd1 vccd1 vccd1 _12234_/X sky130_fd_sc_hd__mux2_1
XFILLER_154_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12165_ _12161_/X _12162_/X _12168_/A vssd1 vssd1 vccd1 vccd1 _12165_/X sky130_fd_sc_hd__mux2_1
XFILLER_151_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11116_ _11048_/Y _11065_/X _11070_/X _11307_/A _08233_/B vssd1 vssd1 vccd1 vccd1
+ _11116_/X sky130_fd_sc_hd__o221a_1
XFILLER_1_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12096_ _12092_/X _12093_/X _12168_/A vssd1 vssd1 vccd1 vccd1 _12096_/X sky130_fd_sc_hd__mux2_1
XFILLER_96_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11047_ _11371_/A _11047_/B vssd1 vssd1 vccd1 vccd1 _11047_/Y sky130_fd_sc_hd__nor2_4
XFILLER_7_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput9 ext_read_data[17] vssd1 vssd1 vccd1 vccd1 input9/X sky130_fd_sc_hd__clkbuf_4
XFILLER_65_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14806_ _15438_/CLK _14806_/D vssd1 vssd1 vccd1 vccd1 hold7/A sky130_fd_sc_hd__dfxtp_1
XTAP_3670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12998_ _15479_/Q _13093_/A2 _13116_/C _12997_/X vssd1 vssd1 vccd1 vccd1 _15479_/D
+ sky130_fd_sc_hd__a22o_1
XTAP_3692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14737_ _15589_/CLK _14737_/D vssd1 vssd1 vccd1 vccd1 _14737_/Q sky130_fd_sc_hd__dfxtp_4
X_11949_ _11942_/X _11944_/X _11946_/X _11948_/X _06671_/A vssd1 vssd1 vccd1 vccd1
+ _11949_/X sky130_fd_sc_hd__o221a_1
Xclkbuf_leaf_71_clk clkbuf_5_14_0_clk/X vssd1 vssd1 vccd1 vccd1 _15599_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_2980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14668_ _15641_/CLK _14668_/D vssd1 vssd1 vccd1 vccd1 _14668_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_177_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13619_ _14493_/CLK _13619_/D vssd1 vssd1 vccd1 vccd1 _13619_/Q sky130_fd_sc_hd__dfxtp_1
X_14599_ _15375_/CLK _14599_/D vssd1 vssd1 vccd1 vccd1 _14599_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_119_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07140_ _14850_/Q _14842_/Q _07146_/S vssd1 vssd1 vccd1 vccd1 _07140_/X sky130_fd_sc_hd__mux2_1
XFILLER_119_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07071_ _07070_/X _14756_/Q _07077_/S vssd1 vssd1 vccd1 vccd1 _13602_/D sky130_fd_sc_hd__mux2_1
XFILLER_156_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07973_ _13559_/Q _13558_/Q _13557_/Q _07973_/D vssd1 vssd1 vccd1 vccd1 _07984_/D
+ sky130_fd_sc_hd__and4_2
XFILLER_101_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09712_ _13082_/B2 _14082_/Q _09723_/S vssd1 vssd1 vccd1 vccd1 _14082_/D sky130_fd_sc_hd__mux2_1
XFILLER_68_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06924_ _06911_/X _06923_/B _06922_/A vssd1 vssd1 vccd1 vccd1 _06924_/X sky130_fd_sc_hd__a21o_1
XFILLER_45_1083 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09643_ _14016_/Q _13078_/B2 _09660_/S vssd1 vssd1 vccd1 vccd1 _14016_/D sky130_fd_sc_hd__mux2_1
X_06855_ _14894_/Q _06854_/X _14895_/Q vssd1 vssd1 vccd1 vccd1 _06857_/C sky130_fd_sc_hd__o21ai_2
XFILLER_55_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09574_ _13950_/Q _13074_/B2 _09589_/S vssd1 vssd1 vccd1 vccd1 _13950_/D sky130_fd_sc_hd__mux2_1
X_06786_ _14585_/Q _14586_/Q _14584_/Q _14583_/Q vssd1 vssd1 vccd1 vccd1 _06791_/B
+ sky130_fd_sc_hd__or4bb_2
XTAP_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_822 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_287 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08525_ _13648_/Q _08523_/Y _08749_/A2 _13611_/Q vssd1 vssd1 vccd1 vccd1 _08525_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_23_310 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_62_clk _15031_/CLK vssd1 vssd1 vccd1 vccd1 _15580_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_24_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08456_ _13758_/Q _12878_/S _08426_/X _08455_/X vssd1 vssd1 vccd1 vccd1 _13758_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_24_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07407_ _13657_/Q _07483_/A2 _07483_/B1 _14685_/Q _07406_/X vssd1 vssd1 vccd1 vccd1
+ _07407_/X sky130_fd_sc_hd__a221o_1
XFILLER_51_26 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08387_ _11252_/A _08386_/X _08381_/Y vssd1 vssd1 vccd1 vccd1 _11298_/B sky130_fd_sc_hd__o21a_1
XFILLER_167_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07338_ _07327_/Y _07329_/A _07333_/X _07337_/X vssd1 vssd1 vccd1 vccd1 _07362_/A
+ sky130_fd_sc_hd__o211a_1
X_07269_ _07235_/A _07235_/B _07237_/Y _07238_/X _07268_/Y vssd1 vssd1 vccd1 vccd1
+ _07269_/X sky130_fd_sc_hd__o221a_1
XFILLER_100_1019 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09008_ _09524_/A _09008_/B _09008_/C vssd1 vssd1 vccd1 vccd1 _09008_/X sky130_fd_sc_hd__and3_1
X_10280_ _14665_/Q _14818_/Q _10665_/S vssd1 vssd1 vccd1 vccd1 _14665_/D sky130_fd_sc_hd__mux2_1
XFILLER_3_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout540 _13144_/A0 vssd1 vssd1 vccd1 vccd1 _09546_/S1 sky130_fd_sc_hd__buf_12
XFILLER_104_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout551 _08490_/A1 vssd1 vssd1 vccd1 vccd1 _09047_/S sky130_fd_sc_hd__clkbuf_16
XFILLER_116_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout562 _08490_/A1 vssd1 vssd1 vccd1 vccd1 _09551_/S sky130_fd_sc_hd__buf_12
XFILLER_120_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13970_ _15301_/CLK _13970_/D vssd1 vssd1 vccd1 vccd1 _13970_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout573 _08405_/C vssd1 vssd1 vccd1 vccd1 _06671_/A sky130_fd_sc_hd__buf_12
Xfanout584 _12498_/A vssd1 vssd1 vccd1 vccd1 _12465_/S1 sky130_fd_sc_hd__buf_12
Xfanout595 fanout600/X vssd1 vssd1 vccd1 vccd1 _12567_/A sky130_fd_sc_hd__buf_6
XFILLER_86_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12921_ _15449_/Q _15635_/Q _12928_/S vssd1 vssd1 vccd1 vccd1 _15449_/D sky130_fd_sc_hd__mux2_1
XFILLER_58_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15640_ _15643_/CLK _15640_/D vssd1 vssd1 vccd1 vccd1 _15640_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12852_ _14746_/Q _15380_/Q _12866_/S vssd1 vssd1 vccd1 vccd1 _15380_/D sky130_fd_sc_hd__mux2_1
XTAP_2221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11803_ _15226_/Q _13086_/B2 _11817_/S vssd1 vssd1 vccd1 vccd1 _15226_/D sky130_fd_sc_hd__mux2_1
XTAP_2254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15571_ _15572_/CLK _15571_/D vssd1 vssd1 vccd1 vccd1 _15571_/Q sky130_fd_sc_hd__dfxtp_1
X_12783_ _15360_/Q _12789_/C vssd1 vssd1 vccd1 vccd1 _12783_/X sky130_fd_sc_hd__xor2_1
XTAP_1520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14522_ _15649_/CLK _14522_/D vssd1 vssd1 vccd1 vccd1 _14522_/Q sky130_fd_sc_hd__dfxtp_1
X_11734_ _15163_/Q _13342_/A0 _11742_/S vssd1 vssd1 vccd1 vccd1 _15163_/D sky130_fd_sc_hd__mux2_1
XTAP_2298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14453_ _14485_/CLK _14453_/D vssd1 vssd1 vccd1 vccd1 _14453_/Q sky130_fd_sc_hd__dfxtp_1
X_11665_ _11873_/A1 _15097_/Q _11675_/S vssd1 vssd1 vccd1 vccd1 _15097_/D sky130_fd_sc_hd__mux2_1
Xclkbuf_4_6_0_clk clkbuf_4_7_0_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_6_0_clk/X sky130_fd_sc_hd__clkbuf_8
XFILLER_30_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10616_ _15561_/Q _10706_/B vssd1 vssd1 vccd1 vccd1 _10616_/X sky130_fd_sc_hd__and2_1
X_13404_ _15670_/CLK _13404_/D vssd1 vssd1 vccd1 vccd1 _13404_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_186_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14384_ _15200_/CLK _14384_/D vssd1 vssd1 vccd1 vccd1 _14384_/Q sky130_fd_sc_hd__dfxtp_1
X_11596_ _11596_/A _11604_/B vssd1 vssd1 vccd1 vccd1 _11596_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_128_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13335_ _13335_/A0 _15665_/Q _13345_/S vssd1 vssd1 vccd1 vccd1 _15665_/D sky130_fd_sc_hd__mux2_1
X_10547_ _10478_/B _10545_/X _10546_/Y _10557_/B vssd1 vssd1 vccd1 vccd1 _10548_/C
+ sky130_fd_sc_hd__a31o_1
XFILLER_41_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_575 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13266_ _15350_/Q _15597_/Q _13300_/S vssd1 vssd1 vccd1 vccd1 _15597_/D sky130_fd_sc_hd__mux2_1
X_10478_ _10478_/A _10478_/B vssd1 vssd1 vccd1 vccd1 _10527_/A sky130_fd_sc_hd__nand2_1
X_15005_ _15580_/CLK _15005_/D vssd1 vssd1 vccd1 vccd1 _15005_/Q sky130_fd_sc_hd__dfxtp_1
X_12217_ _13953_/Q _13695_/Q _12476_/S vssd1 vssd1 vccd1 vccd1 _12218_/B sky130_fd_sc_hd__mux2_1
X_13197_ _15566_/Q _13241_/A2 _13195_/Y _13196_/X vssd1 vssd1 vccd1 vccd1 _15566_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_123_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12148_ _13950_/Q _13692_/Q _12269_/S vssd1 vssd1 vccd1 vccd1 _12149_/B sky130_fd_sc_hd__mux2_1
XFILLER_69_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12079_ _13947_/Q _13689_/Q _12079_/S vssd1 vssd1 vccd1 vccd1 _12080_/B sky130_fd_sc_hd__mux2_1
XFILLER_2_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_947 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_44_clk clkbuf_5_9_0_clk/X vssd1 vssd1 vccd1 vccd1 _15553_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_178_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08310_ _13720_/Q _08232_/A _11351_/C1 _08309_/Y vssd1 vssd1 vccd1 vccd1 _13720_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_178_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09290_ _14473_/Q _09558_/A2 _09289_/X _13049_/A1 vssd1 vssd1 vccd1 vccd1 _09290_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_75_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08241_ _13774_/Q _08237_/A _07331_/A _10457_/A2 _08240_/X vssd1 vssd1 vccd1 vccd1
+ _08241_/Y sky130_fd_sc_hd__a221oi_4
XANTENNA_14 _10734_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_25 _14863_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_36 _15030_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_47 input24/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08172_ _13673_/Q _10285_/S _08155_/X _08171_/X vssd1 vssd1 vccd1 vccd1 _13673_/D
+ sky130_fd_sc_hd__o22a_1
XANTENNA_58 _07168_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_69 _07135_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07123_ _07131_/A _07123_/B vssd1 vssd1 vccd1 vccd1 _07123_/X sky130_fd_sc_hd__and2_2
XFILLER_146_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07054_ _14630_/Q _14662_/Q _07078_/S vssd1 vssd1 vccd1 vccd1 _07054_/X sky130_fd_sc_hd__mux2_1
XFILLER_146_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_1071 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07956_ _07958_/B _07955_/X _07964_/A vssd1 vssd1 vccd1 vccd1 _07956_/X sky130_fd_sc_hd__a21bo_1
XFILLER_87_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_999 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06907_ _15381_/Q _06727_/Y _15380_/Q _06729_/Y vssd1 vssd1 vccd1 vccd1 _06907_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_68_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07887_ _07900_/C _07886_/Y _07903_/A vssd1 vssd1 vccd1 vccd1 _07887_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_95_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09626_ _14000_/Q _11881_/A1 _09628_/S vssd1 vssd1 vccd1 vccd1 _14000_/D sky130_fd_sc_hd__mux2_1
X_06838_ _08508_/B _06845_/B _06681_/Y _13125_/B vssd1 vssd1 vccd1 vccd1 _06838_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_55_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09557_ _15680_/Q _13414_/Q _09557_/S vssd1 vssd1 vccd1 vccd1 _09557_/X sky130_fd_sc_hd__mux2_1
XFILLER_70_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06769_ _13229_/A vssd1 vssd1 vccd1 vccd1 _06769_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_43_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_35_clk clkbuf_5_13_0_clk/X vssd1 vssd1 vccd1 vccd1 _14861_/CLK sky130_fd_sc_hd__clkbuf_16
X_08508_ _08668_/C _08508_/B vssd1 vssd1 vccd1 vccd1 _08508_/Y sky130_fd_sc_hd__nor2_8
XFILLER_54_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09488_ _14546_/Q _14159_/Q _14191_/Q _14127_/Q _09551_/S _09550_/A1 vssd1 vssd1
+ vccd1 vccd1 _09488_/X sky130_fd_sc_hd__mux4_1
XFILLER_23_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08439_ _06676_/A _08390_/C _08425_/X _10764_/S vssd1 vssd1 vccd1 vccd1 _08439_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_12_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11450_ _11450_/A _11450_/B vssd1 vssd1 vccd1 vccd1 _11459_/B sky130_fd_sc_hd__and2_1
XFILLER_177_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10401_ _07319_/X _10457_/A2 _10400_/X vssd1 vssd1 vccd1 vccd1 _11414_/D sky130_fd_sc_hd__a21oi_4
X_11381_ _11383_/A _11383_/B vssd1 vssd1 vccd1 vccd1 _11384_/A sky130_fd_sc_hd__nor2_2
XFILLER_137_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13120_ _14597_/Q _15529_/Q _13120_/S vssd1 vssd1 vccd1 vccd1 _15529_/D sky130_fd_sc_hd__mux2_1
XFILLER_109_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10332_ _14717_/Q _14910_/Q _10343_/S vssd1 vssd1 vccd1 vccd1 _14717_/D sky130_fd_sc_hd__mux2_1
XFILLER_109_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13051_ _13118_/A2 _13051_/B vssd1 vssd1 vccd1 vccd1 _13051_/X sky130_fd_sc_hd__and2b_4
XFILLER_105_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10263_ _14648_/Q _14801_/Q _10735_/S vssd1 vssd1 vccd1 vccd1 _14648_/D sky130_fd_sc_hd__mux2_1
X_12002_ _14523_/Q _14136_/Q _14168_/Q _14104_/Q _12545_/S _12406_/A vssd1 vssd1 vccd1
+ vccd1 _12002_/X sky130_fd_sc_hd__mux4_1
XFILLER_133_771 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10194_ _11847_/A1 _14578_/Q _10197_/S vssd1 vssd1 vccd1 vccd1 _14578_/D sky130_fd_sc_hd__mux2_1
XFILLER_120_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout370 _08507_/Y vssd1 vssd1 vccd1 vccd1 _08668_/D sky130_fd_sc_hd__buf_12
XFILLER_47_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout381 _11259_/S vssd1 vssd1 vccd1 vccd1 _11318_/S sky130_fd_sc_hd__clkbuf_16
Xfanout392 _11414_/A vssd1 vssd1 vccd1 vccd1 _08233_/B sky130_fd_sc_hd__buf_8
XFILLER_87_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13953_ _15658_/CLK _13953_/D vssd1 vssd1 vccd1 vccd1 _13953_/Q sky130_fd_sc_hd__dfxtp_1
X_12904_ _15432_/Q _15618_/Q _12904_/S vssd1 vssd1 vccd1 vccd1 _15432_/D sky130_fd_sc_hd__mux2_1
X_13884_ _15088_/CLK _13884_/D vssd1 vssd1 vccd1 vccd1 _13884_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15623_ _15623_/CLK _15623_/D vssd1 vssd1 vccd1 vccd1 _15623_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12835_ _12828_/A _12833_/Y _12834_/X _12785_/B vssd1 vssd1 vccd1 vccd1 _12835_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_27_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_26_clk clkbuf_5_6_0_clk/X vssd1 vssd1 vccd1 vccd1 _15497_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_2062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15554_ _15556_/CLK _15554_/D vssd1 vssd1 vccd1 vccd1 _15554_/Q sky130_fd_sc_hd__dfxtp_1
X_12766_ _12737_/A _12764_/X _12765_/X _12788_/C1 vssd1 vssd1 vccd1 vccd1 _15357_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_1361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14505_ _15389_/CLK _14505_/D vssd1 vssd1 vccd1 vccd1 _14505_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11717_ _15146_/Q _11858_/A1 _11742_/S vssd1 vssd1 vccd1 vccd1 _15146_/D sky130_fd_sc_hd__mux2_1
XTAP_1394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12697_ _13592_/Q _12696_/X _12763_/S vssd1 vssd1 vccd1 vccd1 _12697_/X sky130_fd_sc_hd__mux2_1
XFILLER_14_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15485_ _15517_/CLK _15485_/D vssd1 vssd1 vccd1 vccd1 _15485_/Q sky130_fd_sc_hd__dfxtp_1
X_11648_ _11681_/A0 _15080_/Q _11670_/S vssd1 vssd1 vccd1 vccd1 _15080_/D sky130_fd_sc_hd__mux2_1
X_14436_ _15556_/CLK _14436_/D vssd1 vssd1 vccd1 vccd1 _14436_/Q sky130_fd_sc_hd__dfxtp_1
Xinput12 ext_read_data[1] vssd1 vssd1 vccd1 vccd1 input12/X sky130_fd_sc_hd__buf_6
Xinput23 ext_read_data[2] vssd1 vssd1 vccd1 vccd1 input23/X sky130_fd_sc_hd__clkbuf_4
Xinput34 meip vssd1 vssd1 vccd1 vccd1 input34/X sky130_fd_sc_hd__buf_6
X_11579_ _11542_/A _11556_/A _11554_/X _11576_/C _11576_/D vssd1 vssd1 vccd1 vccd1
+ _11579_/Y sky130_fd_sc_hd__a2111oi_1
X_14367_ _15220_/CLK _14367_/D vssd1 vssd1 vccd1 vccd1 _14367_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_183_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13318_ _14714_/Q _14715_/Q _13318_/C _13318_/D vssd1 vssd1 vccd1 vccd1 _13318_/X
+ sky130_fd_sc_hd__or4_4
X_14298_ _14462_/CLK _14298_/D vssd1 vssd1 vccd1 vccd1 _14298_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13249_ _13242_/A _11349_/C _13219_/S vssd1 vssd1 vccd1 vccd1 _13249_/X sky130_fd_sc_hd__o21a_1
XFILLER_112_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07810_ _13516_/Q _07810_/B vssd1 vssd1 vccd1 vccd1 _07811_/B sky130_fd_sc_hd__xor2_1
XFILLER_112_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08790_ _11857_/A1 _13816_/Q _08816_/S vssd1 vssd1 vccd1 vccd1 _13816_/D sky130_fd_sc_hd__mux2_1
XFILLER_112_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07741_ _14755_/Q _07736_/A _07740_/Y _08002_/C1 vssd1 vssd1 vccd1 vccd1 _13498_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_38_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_1075 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_243 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07672_ _13480_/Q _13479_/Q _07672_/C vssd1 vssd1 vccd1 vccd1 _07679_/C sky130_fd_sc_hd__and3_2
XFILLER_92_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09411_ _10868_/S _09411_/B _09411_/C vssd1 vssd1 vccd1 vccd1 _09411_/X sky130_fd_sc_hd__and3_1
XFILLER_93_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_17_clk clkbuf_5_2_0_clk/X vssd1 vssd1 vccd1 vccd1 _15267_/CLK sky130_fd_sc_hd__clkbuf_16
X_09342_ _15670_/Q _13404_/Q _09342_/S vssd1 vssd1 vccd1 vccd1 _09342_/X sky130_fd_sc_hd__mux2_1
XFILLER_178_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09273_ _14085_/Q _09522_/A2 _08512_/B _14053_/Q _09543_/A vssd1 vssd1 vccd1 vccd1
+ _09273_/X sky130_fd_sc_hd__a221o_1
XFILLER_139_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08224_ _13713_/Q _08232_/A vssd1 vssd1 vccd1 vccd1 _08224_/X sky130_fd_sc_hd__and2_1
XFILLER_166_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08155_ _06661_/Y _14899_/Q _14901_/Q _08151_/X _08119_/X vssd1 vssd1 vccd1 vccd1
+ _08155_/X sky130_fd_sc_hd__a41o_4
XFILLER_146_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07106_ _14900_/Q _14899_/Q vssd1 vssd1 vccd1 vccd1 _08121_/B sky130_fd_sc_hd__nand2_1
XFILLER_134_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08086_ _08086_/A _08086_/B vssd1 vssd1 vccd1 vccd1 _08086_/Y sky130_fd_sc_hd__nand2_1
X_07037_ _07036_/X _13591_/Q _12728_/S vssd1 vssd1 vccd1 vccd1 _07037_/X sky130_fd_sc_hd__mux2_1
XFILLER_164_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08988_ _08988_/A1 _09449_/A1 _08987_/X _09450_/B1 vssd1 vssd1 vccd1 vccd1 _08988_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_102_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07939_ _13550_/Q _07946_/D vssd1 vssd1 vccd1 vccd1 _07943_/B sky130_fd_sc_hd__nand2_1
XFILLER_21_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10950_ _14960_/Q _10429_/A _10951_/B vssd1 vssd1 vccd1 vccd1 _14960_/D sky130_fd_sc_hd__mux2_1
XFILLER_56_574 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09609_ _13983_/Q _11689_/A0 _09627_/S vssd1 vssd1 vccd1 vccd1 _13983_/D sky130_fd_sc_hd__mux2_1
XFILLER_83_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10881_ _14913_/Q _15544_/Q _13134_/A vssd1 vssd1 vccd1 vccd1 _14913_/D sky130_fd_sc_hd__mux2_1
XFILLER_73_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12620_ _15337_/Q _13149_/S _12619_/X vssd1 vssd1 vccd1 vccd1 _15337_/D sky130_fd_sc_hd__a21o_1
XFILLER_71_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12551_ _15334_/Q _13149_/S _12550_/X vssd1 vssd1 vccd1 vccd1 _15334_/D sky130_fd_sc_hd__a21o_1
XFILLER_145_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11502_ _11502_/A _11502_/B vssd1 vssd1 vccd1 vccd1 _11502_/Y sky130_fd_sc_hd__nor2_1
XFILLER_185_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15270_ _15335_/CLK _15270_/D vssd1 vssd1 vccd1 vccd1 _15270_/Q sky130_fd_sc_hd__dfxtp_1
X_12482_ _15331_/Q _13081_/A2 _12481_/X vssd1 vssd1 vccd1 vccd1 _15331_/D sky130_fd_sc_hd__a21o_1
XFILLER_11_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11433_ _11418_/X _11425_/B _11420_/A vssd1 vssd1 vccd1 vccd1 _11441_/B sky130_fd_sc_hd__o21a_1
XFILLER_172_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14221_ _15662_/CLK _14221_/D vssd1 vssd1 vccd1 vccd1 _14221_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_153_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14152_ _15161_/CLK _14152_/D vssd1 vssd1 vccd1 vccd1 _14152_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11364_ _11363_/B _11363_/C _13162_/B vssd1 vssd1 vccd1 vccd1 _11365_/B sky130_fd_sc_hd__a21bo_1
XFILLER_180_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10315_ _14700_/Q _14885_/Q _10695_/S vssd1 vssd1 vccd1 vccd1 _14700_/D sky130_fd_sc_hd__mux2_1
X_13103_ _15519_/Q _13119_/S _13105_/B1 _13102_/X vssd1 vssd1 vccd1 vccd1 _15519_/D
+ sky130_fd_sc_hd__a22o_1
X_14083_ _14083_/CLK _14083_/D vssd1 vssd1 vccd1 vccd1 _14083_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_579 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11295_ _11280_/B _11294_/Y _11318_/S vssd1 vssd1 vccd1 vccd1 _11296_/A sky130_fd_sc_hd__mux2_1
XFILLER_65_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13034_ _15491_/Q _10877_/S _13116_/C _13033_/X vssd1 vssd1 vccd1 vccd1 _15491_/D
+ sky130_fd_sc_hd__a22o_1
X_10246_ _14631_/Q _14784_/Q _10665_/S vssd1 vssd1 vccd1 vccd1 _14631_/D sky130_fd_sc_hd__mux2_1
XFILLER_112_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10177_ _13330_/A0 _14561_/Q _10192_/S vssd1 vssd1 vccd1 vccd1 _14561_/D sky130_fd_sc_hd__mux2_1
XFILLER_79_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14985_ _15582_/CLK _14985_/D vssd1 vssd1 vccd1 vccd1 _14985_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_93_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_80 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13936_ _15526_/CLK _13936_/D vssd1 vssd1 vccd1 vccd1 _13936_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13867_ _15510_/CLK _13867_/D vssd1 vssd1 vccd1 vccd1 _13867_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15606_ _15606_/CLK _15606_/D vssd1 vssd1 vccd1 vccd1 _15606_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_1100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12818_ _15365_/Q _12819_/B vssd1 vssd1 vccd1 vccd1 _12827_/B sky130_fd_sc_hd__and2_2
XFILLER_22_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13798_ _13798_/CLK _13798_/D vssd1 vssd1 vccd1 vccd1 _13798_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_16_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15537_ _15537_/CLK _15537_/D vssd1 vssd1 vccd1 vccd1 hold3/A sky130_fd_sc_hd__dfxtp_1
X_12749_ _13599_/Q _12748_/X _12785_/B vssd1 vssd1 vccd1 vccd1 _12749_/X sky130_fd_sc_hd__mux2_1
XFILLER_31_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15468_ _15500_/CLK _15468_/D vssd1 vssd1 vccd1 vccd1 _15468_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_175_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14419_ _15226_/CLK _14419_/D vssd1 vssd1 vccd1 vccd1 _14419_/Q sky130_fd_sc_hd__dfxtp_1
X_15399_ _15399_/CLK _15399_/D vssd1 vssd1 vccd1 vccd1 _15399_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_116_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09960_ _11847_/A1 _14320_/Q _09963_/S vssd1 vssd1 vccd1 vccd1 _14320_/D sky130_fd_sc_hd__mux2_1
XFILLER_104_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_6_clk clkbuf_5_1_0_clk/X vssd1 vssd1 vccd1 vccd1 _15658_/CLK sky130_fd_sc_hd__clkbuf_16
X_08911_ _08508_/B _08519_/B _08910_/X _13049_/A1 vssd1 vssd1 vccd1 vccd1 _08911_/X
+ sky130_fd_sc_hd__a31o_1
XTAP_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09891_ _11877_/A1 _14253_/Q _09892_/S vssd1 vssd1 vccd1 vccd1 _14253_/D sky130_fd_sc_hd__mux2_1
XTAP_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08842_ _13865_/Q _11874_/A1 _08851_/S vssd1 vssd1 vccd1 vccd1 _13865_/D sky130_fd_sc_hd__mux2_1
XFILLER_58_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08773_ _08773_/A _08773_/B _08753_/X vssd1 vssd1 vccd1 vccd1 _08773_/Y sky130_fd_sc_hd__nor3b_1
XFILLER_38_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07724_ _13494_/Q _13493_/Q _07724_/C vssd1 vssd1 vccd1 vccd1 _07727_/B sky130_fd_sc_hd__and3_2
XFILLER_150_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07655_ _07655_/A _07655_/B _07655_/C vssd1 vssd1 vccd1 vccd1 _07665_/C sky130_fd_sc_hd__and3_2
XFILLER_168_1063 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07586_ _14746_/Q _07607_/A _07585_/Y _12809_/C1 vssd1 vssd1 vccd1 vccd1 _13457_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_81_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09325_ _14377_/Q _15193_/Q _13832_/Q _14571_/Q _09342_/S _13144_/A0 vssd1 vssd1
+ vccd1 vccd1 _09326_/B sky130_fd_sc_hd__mux4_1
XFILLER_159_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_914 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_402 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09256_ _15125_/Q _09558_/A2 _08540_/B _15093_/Q _09255_/X vssd1 vssd1 vccd1 vccd1
+ _09256_/X sky130_fd_sc_hd__a221o_1
XFILLER_166_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08207_ _13698_/Q _11761_/A0 _08221_/S vssd1 vssd1 vccd1 vccd1 _13698_/D sky130_fd_sc_hd__mux2_1
XFILLER_5_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09187_ _14017_/Q _13985_/Q _09425_/S vssd1 vssd1 vccd1 vccd1 _09187_/X sky130_fd_sc_hd__mux2_1
XFILLER_135_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08138_ _08133_/S _06763_/Y _08151_/S vssd1 vssd1 vccd1 vccd1 _08138_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_181_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08069_ _14762_/Q _13640_/Q _08072_/S vssd1 vssd1 vccd1 vccd1 _13640_/D sky130_fd_sc_hd__mux2_1
XFILLER_135_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10100_ _14486_/Q _14734_/Q _10131_/S vssd1 vssd1 vccd1 vccd1 _14486_/D sky130_fd_sc_hd__mux2_1
XFILLER_122_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11080_ _11259_/S _11007_/B _11324_/A _11079_/Y vssd1 vssd1 vccd1 vccd1 _11080_/X
+ sky130_fd_sc_hd__a31o_2
XFILLER_89_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10031_ _12832_/C1 _13581_/Q _08030_/Y _06997_/B _14389_/Q vssd1 vssd1 vccd1 vccd1
+ _14389_/D sky130_fd_sc_hd__a32o_1
XFILLER_49_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14770_ _15587_/CLK _14770_/D vssd1 vssd1 vccd1 vccd1 _14770_/Q sky130_fd_sc_hd__dfxtp_1
X_11982_ _14360_/Q _15176_/Q _13815_/Q _14554_/Q _12154_/S _12253_/S1 vssd1 vssd1
+ vccd1 vccd1 _11982_/X sky130_fd_sc_hd__mux4_1
XFILLER_91_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13721_ _15020_/CLK _13721_/D vssd1 vssd1 vccd1 vccd1 _13721_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10933_ _14950_/Q _10511_/Y _10948_/B vssd1 vssd1 vccd1 vccd1 _14950_/D sky130_fd_sc_hd__mux2_1
XFILLER_147_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10864_ _13737_/Q _14896_/Q _13129_/A vssd1 vssd1 vccd1 vccd1 _14896_/D sky130_fd_sc_hd__mux2_1
X_13652_ _15620_/CLK _13652_/D vssd1 vssd1 vccd1 vccd1 _13652_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_182_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12603_ _14387_/Q _15203_/Q _13842_/Q _14581_/Q _12612_/S _12613_/A vssd1 vssd1 vccd1
+ vccd1 _12603_/X sky130_fd_sc_hd__mux4_1
XPHY_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13583_ _15619_/CLK _13583_/D vssd1 vssd1 vccd1 vccd1 _13583_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10795_ _14827_/Q _15459_/Q _12933_/S vssd1 vssd1 vccd1 vccd1 _14827_/D sky130_fd_sc_hd__mux2_1
XFILLER_169_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15322_ _15510_/CLK _15322_/D vssd1 vssd1 vccd1 vccd1 _15322_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12534_ _14384_/Q _15200_/Q _13839_/Q _14578_/Q _12612_/S _12613_/A vssd1 vssd1 vccd1
+ vccd1 _12534_/X sky130_fd_sc_hd__mux4_1
XFILLER_184_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15253_ _15253_/CLK _15253_/D vssd1 vssd1 vccd1 vccd1 _15253_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_184_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12465_ _14381_/Q _15197_/Q _13836_/Q _14575_/Q _12472_/S _12465_/S1 vssd1 vssd1
+ vccd1 vccd1 _12465_/X sky130_fd_sc_hd__mux4_1
XFILLER_173_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_1074 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14204_ _15281_/CLK _14204_/D vssd1 vssd1 vccd1 vccd1 _14204_/Q sky130_fd_sc_hd__dfxtp_1
X_11416_ _11436_/A _11416_/B vssd1 vssd1 vccd1 vccd1 _11419_/B sky130_fd_sc_hd__xnor2_1
X_12396_ _14378_/Q _15194_/Q _13833_/Q _14572_/Q _12591_/S _12590_/A vssd1 vssd1 vccd1
+ vccd1 _12396_/X sky130_fd_sc_hd__mux4_1
X_15184_ _15184_/CLK _15184_/D vssd1 vssd1 vccd1 vccd1 _15184_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_126_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14135_ _15273_/CLK _14135_/D vssd1 vssd1 vccd1 vccd1 _14135_/Q sky130_fd_sc_hd__dfxtp_1
X_11347_ _11347_/A _11347_/B vssd1 vssd1 vccd1 vccd1 _11347_/Y sky130_fd_sc_hd__nand2_1
XFILLER_113_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11278_ _15031_/Q wire438/X _11276_/X _11277_/X vssd1 vssd1 vccd1 vccd1 _15031_/D
+ sky130_fd_sc_hd__o22a_1
X_14066_ _15667_/CLK _14066_/D vssd1 vssd1 vccd1 vccd1 _14066_/Q sky130_fd_sc_hd__dfxtp_1
X_13017_ _10699_/X _14886_/Q _13029_/S vssd1 vssd1 vccd1 vccd1 _13017_/X sky130_fd_sc_hd__mux2_8
X_10229_ input25/X _14614_/Q _13282_/S vssd1 vssd1 vccd1 vccd1 _14614_/D sky130_fd_sc_hd__mux2_1
XFILLER_140_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1 hold1/A vssd1 vssd1 vccd1 vccd1 hold1/X sky130_fd_sc_hd__bufbuf_16
XFILLER_55_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14968_ _15000_/CLK _14968_/D vssd1 vssd1 vccd1 vccd1 _14968_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_894 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13919_ _15508_/CLK _13919_/D vssd1 vssd1 vccd1 vccd1 _13919_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_62_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14899_ _15536_/CLK _14899_/D vssd1 vssd1 vccd1 vccd1 _14899_/Q sky130_fd_sc_hd__dfxtp_2
X_07440_ _14750_/Q _07439_/X _07480_/S vssd1 vssd1 vccd1 vccd1 _07440_/X sky130_fd_sc_hd__mux2_8
XFILLER_63_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07371_ _14645_/Q _07498_/B _07498_/C vssd1 vssd1 vccd1 vccd1 _07371_/X sky130_fd_sc_hd__and3_1
XFILLER_50_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09110_ _09427_/A1 _09108_/X _09109_/X vssd1 vssd1 vccd1 vccd1 _09110_/X sky130_fd_sc_hd__a21o_1
XFILLER_128_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09041_ _14461_/Q _14429_/Q _13850_/Q _14203_/Q _09225_/S0 _09225_/S1 vssd1 vssd1
+ vccd1 vccd1 _09041_/X sky130_fd_sc_hd__mux4_2
XFILLER_148_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09943_ _13330_/A0 _14303_/Q _09958_/S vssd1 vssd1 vccd1 vccd1 _14303_/D sky130_fd_sc_hd__mux2_1
XFILLER_132_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09874_ _11860_/A1 _14236_/Q _09892_/S vssd1 vssd1 vccd1 vccd1 _14236_/D sky130_fd_sc_hd__mux2_1
XFILLER_97_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08825_ _13848_/Q _11649_/A0 _08851_/S vssd1 vssd1 vccd1 vccd1 _13848_/D sky130_fd_sc_hd__mux2_1
XTAP_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08756_ _14597_/Q _08756_/B vssd1 vssd1 vccd1 vccd1 _08777_/B sky130_fd_sc_hd__nor2_2
XFILLER_39_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07707_ _14746_/Q _07713_/A _07706_/Y _07949_/C1 vssd1 vssd1 vccd1 vccd1 _13489_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_26_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08687_ _14495_/Q _08693_/A2 _08685_/X _08686_/X vssd1 vssd1 vccd1 vccd1 _08688_/C
+ sky130_fd_sc_hd__a211o_1
XTAP_1905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07638_ _13471_/Q _07635_/B _13472_/Q vssd1 vssd1 vccd1 vccd1 _07638_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_13_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_547 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07569_ _14742_/Q _07629_/A _07568_/Y _07949_/C1 vssd1 vssd1 vccd1 vccd1 _13453_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_110_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09308_ _14248_/Q _14280_/Q _14312_/Q _14344_/Q _09481_/S _09553_/A1 vssd1 vssd1
+ vccd1 vccd1 _09308_/X sky130_fd_sc_hd__mux4_1
XFILLER_10_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10580_ _14995_/Q _10569_/B _10733_/A2 _14963_/Q _10732_/C1 vssd1 vssd1 vccd1 vccd1
+ _10580_/X sky130_fd_sc_hd__a221o_1
XFILLER_167_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09239_ _15290_/Q _15258_/Q _15226_/Q _15157_/Q _09535_/S _08494_/B vssd1 vssd1 vccd1
+ vccd1 _09239_/X sky130_fd_sc_hd__mux4_1
XFILLER_10_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12250_ _12503_/A1 _12249_/X _12248_/X _12503_/C1 vssd1 vssd1 vccd1 vccd1 _12251_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_108_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_459 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11201_ _13217_/A _11380_/A vssd1 vssd1 vccd1 vccd1 _11389_/C sky130_fd_sc_hd__nand2_1
XFILLER_119_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12181_ _12503_/A1 _12180_/X _12179_/X _12503_/C1 vssd1 vssd1 vccd1 vccd1 _12182_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_135_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11132_ _10981_/X _10994_/X _11283_/A vssd1 vssd1 vccd1 vccd1 _11132_/X sky130_fd_sc_hd__mux2_1
XFILLER_150_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_677 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11063_ _11058_/Y _11062_/X _11129_/A vssd1 vssd1 vccd1 vccd1 _11175_/B sky130_fd_sc_hd__mux2_2
XFILLER_135_62 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10014_ _11868_/A1 _14372_/Q _10028_/S vssd1 vssd1 vccd1 vccd1 _14372_/D sky130_fd_sc_hd__mux2_1
XFILLER_95_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14822_ _15606_/CLK _14822_/D vssd1 vssd1 vccd1 vccd1 _14822_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_76_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14753_ _15636_/CLK _14753_/D vssd1 vssd1 vccd1 vccd1 _14753_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_3874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11965_ _12080_/A _11965_/B vssd1 vssd1 vccd1 vccd1 _11965_/X sky130_fd_sc_hd__and2_1
XTAP_3885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13704_ _15328_/CLK _13704_/D vssd1 vssd1 vccd1 vccd1 _13704_/Q sky130_fd_sc_hd__dfxtp_1
X_10916_ _11476_/A _10944_/B vssd1 vssd1 vccd1 vccd1 _10916_/Y sky130_fd_sc_hd__nand2_1
XFILLER_45_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14684_ _15589_/CLK _14684_/D vssd1 vssd1 vccd1 vccd1 _14684_/Q sky130_fd_sc_hd__dfxtp_1
X_11896_ _12268_/A _11896_/B vssd1 vssd1 vccd1 vccd1 _11896_/X sky130_fd_sc_hd__and2_1
X_13635_ _14510_/CLK _13635_/D vssd1 vssd1 vccd1 vccd1 _13635_/Q sky130_fd_sc_hd__dfxtp_1
X_10847_ _14879_/Q _13789_/Q _12928_/S vssd1 vssd1 vccd1 vccd1 _14879_/D sky130_fd_sc_hd__mux2_1
XFILLER_158_744 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13566_ _14511_/CLK _13566_/D vssd1 vssd1 vccd1 vccd1 _13566_/Q sky130_fd_sc_hd__dfxtp_2
X_10778_ _14810_/Q _15442_/Q _12917_/S vssd1 vssd1 vccd1 vccd1 _14810_/D sky130_fd_sc_hd__mux2_1
XFILLER_8_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15305_ _15648_/CLK _15305_/D vssd1 vssd1 vccd1 vccd1 _15305_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_157_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12517_ _12521_/A _12517_/B vssd1 vssd1 vccd1 vccd1 _12517_/X sky130_fd_sc_hd__and2_1
XFILLER_8_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13497_ _13632_/CLK _13497_/D vssd1 vssd1 vccd1 vccd1 _13497_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_158_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15236_ _15544_/CLK _15236_/D vssd1 vssd1 vccd1 vccd1 _15236_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_161_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12448_ _12452_/A _12448_/B vssd1 vssd1 vccd1 vccd1 _12448_/X sky130_fd_sc_hd__and2_1
XFILLER_154_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15167_ _15544_/CLK _15167_/D vssd1 vssd1 vccd1 vccd1 _15167_/Q sky130_fd_sc_hd__dfxtp_1
X_12379_ _12379_/A _12379_/B vssd1 vssd1 vccd1 vccd1 _12379_/X sky130_fd_sc_hd__and2_1
X_14118_ _15668_/CLK _14118_/D vssd1 vssd1 vccd1 vccd1 _14118_/Q sky130_fd_sc_hd__dfxtp_1
X_15098_ _15130_/CLK _15098_/D vssd1 vssd1 vccd1 vccd1 _15098_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06940_ _14500_/Q _06724_/Y _14499_/Q _06726_/Y vssd1 vssd1 vccd1 vccd1 _06944_/B
+ sky130_fd_sc_hd__a22o_2
XFILLER_140_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14049_ _15133_/CLK _14049_/D vssd1 vssd1 vccd1 vccd1 _14049_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_140_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06871_ _06879_/A _06871_/B vssd1 vssd1 vccd1 vccd1 _06871_/Y sky130_fd_sc_hd__nor2_1
XFILLER_121_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08610_ _13497_/Q _08691_/B1 _08693_/B1 _13632_/Q vssd1 vssd1 vccd1 vccd1 _08610_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_55_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_230_clk clkbuf_5_6_0_clk/X vssd1 vssd1 vccd1 vccd1 _15661_/CLK sky130_fd_sc_hd__clkbuf_16
X_09590_ _13966_/Q _13346_/A0 _09594_/S vssd1 vssd1 vccd1 vccd1 _13966_/D sky130_fd_sc_hd__mux2_1
XFILLER_82_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08541_ _13610_/Q _08749_/A2 _08747_/B1 _13507_/Q _08540_/X vssd1 vssd1 vccd1 vccd1
+ _08541_/X sky130_fd_sc_hd__a221o_1
XFILLER_47_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08472_ _13765_/Q _10764_/S _08470_/X _14612_/Q vssd1 vssd1 vccd1 vccd1 _13765_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_51_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_1044 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07423_ _13661_/Q _07483_/A2 _07483_/B1 _14689_/Q _07422_/X vssd1 vssd1 vccd1 vccd1
+ _07423_/X sky130_fd_sc_hd__a221o_1
XFILLER_24_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07354_ _07235_/X _07269_/X _07363_/A _07353_/X vssd1 vssd1 vccd1 vccd1 _07355_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_149_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07285_ _15319_/Q _15475_/Q _07340_/S vssd1 vssd1 vccd1 vccd1 _07287_/B sky130_fd_sc_hd__mux2_4
XFILLER_164_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_118 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09024_ _09421_/A1 _09020_/X _09023_/X _09019_/X vssd1 vssd1 vccd1 vccd1 _09024_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_145_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09926_ _11879_/A1 _14287_/Q _09930_/S vssd1 vssd1 vccd1 vccd1 _14287_/D sky130_fd_sc_hd__mux2_1
XFILLER_120_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_444 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09857_ _14221_/Q _13344_/A0 _09858_/S vssd1 vssd1 vccd1 vccd1 _14221_/D sky130_fd_sc_hd__mux2_1
XFILLER_100_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_221_clk clkbuf_5_18_0_clk/X vssd1 vssd1 vccd1 vccd1 _15499_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_3115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08808_ _13098_/B2 _13834_/Q _08816_/S vssd1 vssd1 vccd1 vccd1 _13834_/D sky130_fd_sc_hd__mux2_1
XFILLER_58_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09788_ _14155_/Q _13343_/A0 _09790_/S vssd1 vssd1 vccd1 vccd1 _14155_/D sky130_fd_sc_hd__mux2_1
XFILLER_100_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08739_ _13804_/Q _08573_/S _08736_/X _08738_/X vssd1 vssd1 vccd1 vccd1 _13804_/D
+ sky130_fd_sc_hd__o22a_1
XANTENNA_104 _13799_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_115 input20/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_126 _12515_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11750_ _11858_/A1 _15178_/Q _11775_/S vssd1 vssd1 vccd1 vccd1 _15178_/D sky130_fd_sc_hd__mux2_1
XTAP_1724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_480 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10701_ _15578_/Q _10706_/B vssd1 vssd1 vccd1 vccd1 _10701_/X sky130_fd_sc_hd__and2_1
XFILLER_14_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11681_ _11681_/A0 _15112_/Q _11703_/S vssd1 vssd1 vccd1 vccd1 _15112_/D sky130_fd_sc_hd__mux2_1
XTAP_1779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13420_ _14493_/CLK _13420_/D vssd1 vssd1 vccd1 vccd1 _13420_/Q sky130_fd_sc_hd__dfxtp_1
X_10632_ _13724_/Q _10652_/B vssd1 vssd1 vccd1 vccd1 _10632_/X sky130_fd_sc_hd__and2_1
XFILLER_139_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13351_ _14454_/Q vssd1 vssd1 vccd1 vccd1 _14454_/D sky130_fd_sc_hd__clkbuf_2
X_10563_ _11777_/B _10563_/B vssd1 vssd1 vccd1 vccd1 _10564_/A sky130_fd_sc_hd__and2b_1
XFILLER_10_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12302_ _15126_/Q _15094_/Q _15667_/Q _13401_/Q _12614_/S _12383_/A vssd1 vssd1 vccd1
+ vccd1 _12302_/X sky130_fd_sc_hd__mux4_1
XFILLER_127_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10494_ _08244_/A _13758_/Q _15414_/Q _08244_/B vssd1 vssd1 vccd1 vccd1 _10494_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_5_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13282_ _15366_/Q _15613_/Q _13282_/S vssd1 vssd1 vccd1 vccd1 _15613_/D sky130_fd_sc_hd__mux2_1
XFILLER_6_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15021_ _15021_/CLK _15021_/D vssd1 vssd1 vccd1 vccd1 _15021_/Q sky130_fd_sc_hd__dfxtp_1
X_12233_ _15123_/Q _15091_/Q _15664_/Q _13398_/Q _12499_/S _12486_/S1 vssd1 vssd1
+ vccd1 vccd1 _12233_/X sky130_fd_sc_hd__mux4_1
X_12164_ _15120_/Q _15088_/Q _15661_/Q _13395_/Q _12246_/S _12452_/A vssd1 vssd1 vccd1
+ vccd1 _12164_/X sky130_fd_sc_hd__mux4_1
XFILLER_151_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11115_ _11059_/X _11066_/X _11115_/S vssd1 vssd1 vccd1 vccd1 _11161_/B sky130_fd_sc_hd__mux2_1
X_12095_ _15117_/Q _15085_/Q _15658_/Q _13392_/Q _12476_/S _12498_/A vssd1 vssd1 vccd1
+ vccd1 _12095_/X sky130_fd_sc_hd__mux4_1
XFILLER_96_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11046_ _11044_/Y _11045_/Y _11356_/B vssd1 vssd1 vccd1 vccd1 _11046_/X sky130_fd_sc_hd__mux2_1
XFILLER_7_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_212_clk clkbuf_5_17_0_clk/X vssd1 vssd1 vccd1 vccd1 _15226_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_49_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14805_ _15623_/CLK _14805_/D vssd1 vssd1 vccd1 vccd1 _14805_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_188_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12997_ _13086_/B2 _13039_/A2 _12996_/X _12944_/A vssd1 vssd1 vccd1 vccd1 _12997_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_188_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14736_ _15619_/CLK _14736_/D vssd1 vssd1 vccd1 vccd1 _14736_/Q sky130_fd_sc_hd__dfxtp_4
X_11948_ _12615_/A1 _11947_/X _12615_/B1 vssd1 vssd1 vccd1 vccd1 _11948_/X sky130_fd_sc_hd__a21o_1
XTAP_2970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_5_15_0_clk clkbuf_4_7_0_clk/X vssd1 vssd1 vccd1 vccd1 clkbuf_5_15_0_clk/X
+ sky130_fd_sc_hd__clkbuf_8
XTAP_2981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14667_ _15452_/CLK _14667_/D vssd1 vssd1 vccd1 vccd1 _14667_/Q sky130_fd_sc_hd__dfxtp_1
X_11879_ _15300_/Q _11879_/A1 _11883_/S vssd1 vssd1 vccd1 vccd1 _15300_/D sky130_fd_sc_hd__mux2_1
X_13618_ _15374_/CLK _13618_/D vssd1 vssd1 vccd1 vccd1 _13618_/Q sky130_fd_sc_hd__dfxtp_1
X_14598_ _15588_/CLK _14598_/D vssd1 vssd1 vccd1 vccd1 _14598_/Q sky130_fd_sc_hd__dfxtp_4
X_13549_ _13798_/CLK _13549_/D vssd1 vssd1 vccd1 vccd1 _13549_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07070_ _07069_/X _13602_/Q _12764_/S vssd1 vssd1 vccd1 vccd1 _07070_/X sky130_fd_sc_hd__mux2_1
XFILLER_173_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15219_ _15662_/CLK _15219_/D vssd1 vssd1 vccd1 vccd1 _15219_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07972_ _14751_/Q _07971_/A _07971_/Y _07987_/C1 vssd1 vssd1 vccd1 vccd1 _13558_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_102_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09711_ _13333_/A0 _14081_/Q _09723_/S vssd1 vssd1 vccd1 vccd1 _14081_/D sky130_fd_sc_hd__mux2_1
X_06923_ _06923_/A _06923_/B _06923_/C vssd1 vssd1 vccd1 vccd1 _06923_/X sky130_fd_sc_hd__or3_2
XFILLER_101_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_1095 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_203_clk clkbuf_5_16_0_clk/X vssd1 vssd1 vccd1 vccd1 _15295_/CLK sky130_fd_sc_hd__clkbuf_16
X_09642_ _14015_/Q _11689_/A0 _09660_/S vssd1 vssd1 vccd1 vccd1 _14015_/D sky130_fd_sc_hd__mux2_1
X_06854_ _14926_/Q _14925_/Q vssd1 vssd1 vccd1 vccd1 _06854_/X sky130_fd_sc_hd__xor2_1
X_09573_ _13949_/Q _13072_/B2 _09589_/S vssd1 vssd1 vccd1 vccd1 _13949_/D sky130_fd_sc_hd__mux2_1
X_06785_ _14586_/Q _08469_/A vssd1 vssd1 vccd1 vccd1 _08421_/A sky130_fd_sc_hd__nand2b_2
XFILLER_35_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08524_ _08537_/A _08532_/B vssd1 vssd1 vccd1 vccd1 _08524_/Y sky130_fd_sc_hd__nor2_4
XFILLER_64_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_322 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08455_ _14599_/Q _08773_/B vssd1 vssd1 vccd1 vccd1 _08455_/X sky130_fd_sc_hd__and2_1
XFILLER_168_327 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07406_ _14653_/Q _07490_/B _07482_/C vssd1 vssd1 vccd1 vccd1 _07406_/X sky130_fd_sc_hd__and3_1
XFILLER_50_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08386_ _08366_/A _08385_/Y _11318_/S vssd1 vssd1 vccd1 vccd1 _08386_/X sky130_fd_sc_hd__mux2_1
XFILLER_52_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07337_ _07337_/A _07337_/B vssd1 vssd1 vccd1 vccd1 _07337_/X sky130_fd_sc_hd__or2_1
XFILLER_167_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_177_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07268_ _07268_/A _07268_/B vssd1 vssd1 vccd1 vccd1 _07268_/Y sky130_fd_sc_hd__nand2_1
XFILLER_109_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09007_ _09511_/S1 _09005_/X _09006_/X vssd1 vssd1 vccd1 vccd1 _09008_/C sky130_fd_sc_hd__a21o_1
XFILLER_3_716 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07199_ _13936_/Q _15523_/Q _07334_/S vssd1 vssd1 vccd1 vccd1 _07228_/A sky130_fd_sc_hd__mux2_8
XFILLER_183_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout530 _09530_/S1 vssd1 vssd1 vccd1 vccd1 _09406_/S1 sky130_fd_sc_hd__buf_12
XFILLER_76_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout541 _08508_/B vssd1 vssd1 vccd1 vccd1 _13144_/A0 sky130_fd_sc_hd__buf_8
Xfanout552 _09438_/S0 vssd1 vssd1 vccd1 vccd1 _09444_/S sky130_fd_sc_hd__buf_12
X_09909_ _13072_/B2 _14270_/Q _09925_/S vssd1 vssd1 vccd1 vccd1 _14270_/D sky130_fd_sc_hd__mux2_1
Xfanout563 _09342_/S vssd1 vssd1 vccd1 vccd1 _09469_/S sky130_fd_sc_hd__buf_12
Xfanout574 _08405_/C vssd1 vssd1 vccd1 vccd1 _12616_/C1 sky130_fd_sc_hd__buf_12
XFILLER_59_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout585 _12061_/A vssd1 vssd1 vccd1 vccd1 _12498_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_74_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12920_ _15448_/Q _15634_/Q _12928_/S vssd1 vssd1 vccd1 vccd1 _15448_/D sky130_fd_sc_hd__mux2_1
Xfanout596 fanout600/X vssd1 vssd1 vccd1 vccd1 _12544_/A sky130_fd_sc_hd__buf_12
XFILLER_19_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12851_ _14745_/Q _15379_/Q _12866_/S vssd1 vssd1 vccd1 vccd1 _15379_/D sky130_fd_sc_hd__mux2_1
XTAP_2211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11802_ _15225_/Q _11868_/A1 _11816_/S vssd1 vssd1 vccd1 vccd1 _15225_/D sky130_fd_sc_hd__mux2_1
XTAP_2244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15570_ _15570_/CLK _15570_/D vssd1 vssd1 vccd1 vccd1 _15570_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12782_ _15359_/Q _12765_/B _12781_/X _12809_/C1 vssd1 vssd1 vccd1 vccd1 _15359_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_1521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14521_ _15303_/CLK _14521_/D vssd1 vssd1 vccd1 vccd1 _14521_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_42_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11733_ _15162_/Q _11874_/A1 _11742_/S vssd1 vssd1 vccd1 vccd1 _15162_/D sky130_fd_sc_hd__mux2_1
XTAP_1554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1034 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_826 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14452_ _15672_/CLK _14452_/D vssd1 vssd1 vccd1 vccd1 _14452_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11664_ _11872_/A1 _15096_/Q _11675_/S vssd1 vssd1 vccd1 vccd1 _15096_/D sky130_fd_sc_hd__mux2_1
XFILLER_109_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13403_ _15259_/CLK _13403_/D vssd1 vssd1 vccd1 vccd1 _13403_/Q sky130_fd_sc_hd__dfxtp_1
X_10615_ _14741_/Q _10614_/X _10615_/S vssd1 vssd1 vccd1 vccd1 _14741_/D sky130_fd_sc_hd__mux2_1
X_14383_ _15199_/CLK _14383_/D vssd1 vssd1 vccd1 vccd1 _14383_/Q sky130_fd_sc_hd__dfxtp_1
X_11595_ _11586_/A _11586_/B _11585_/A vssd1 vssd1 vccd1 vccd1 _11604_/B sky130_fd_sc_hd__a21oi_2
XFILLER_167_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13334_ _13334_/A0 _15664_/Q _13345_/S vssd1 vssd1 vccd1 vccd1 _15664_/D sky130_fd_sc_hd__mux2_1
X_10546_ _10543_/X _10544_/X _10478_/A vssd1 vssd1 vccd1 vccd1 _10546_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_182_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13265_ _15349_/Q _15596_/Q _13300_/S vssd1 vssd1 vccd1 vccd1 _15596_/D sky130_fd_sc_hd__mux2_1
XFILLER_108_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10477_ _11589_/B _13226_/B vssd1 vssd1 vccd1 vccd1 _10478_/B sky130_fd_sc_hd__or2_1
XFILLER_6_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15004_ _15006_/CLK _15004_/D vssd1 vssd1 vccd1 vccd1 _15004_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_142_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12216_ _12503_/A1 _12211_/X _12214_/X _12215_/X _12515_/C1 vssd1 vssd1 vccd1 vccd1
+ _12228_/B sky130_fd_sc_hd__a221o_1
XFILLER_155_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13196_ _06769_/Y _13195_/B _11475_/A _13219_/S vssd1 vssd1 vccd1 vccd1 _13196_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_29_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12147_ _12273_/A1 _12142_/X _12145_/X _12146_/X _08449_/A vssd1 vssd1 vccd1 vccd1
+ _12159_/B sky130_fd_sc_hd__a221o_2
XFILLER_116_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12078_ _12273_/A1 _12073_/X _12076_/X _12077_/X _08449_/A vssd1 vssd1 vccd1 vccd1
+ _12090_/B sky130_fd_sc_hd__a221o_1
XFILLER_77_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11029_ _11029_/A vssd1 vssd1 vccd1 vccd1 _11029_/Y sky130_fd_sc_hd__inv_2
XFILLER_38_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14719_ _15548_/CLK _14719_/D vssd1 vssd1 vccd1 vccd1 _14719_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08240_ _08240_/A _13806_/Q vssd1 vssd1 vccd1 vccd1 _08240_/X sky130_fd_sc_hd__and2_2
XFILLER_178_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_15 _11929_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_26 _14746_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_347 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_37 input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08171_ _08133_/S input17/X _08185_/A vssd1 vssd1 vccd1 vccd1 _08171_/X sky130_fd_sc_hd__and3b_1
XANTENNA_48 input28/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_59 _07168_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07122_ _14841_/Q _14833_/Q _07146_/S vssd1 vssd1 vccd1 vccd1 _07123_/B sky130_fd_sc_hd__mux2_1
XFILLER_146_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07053_ _07052_/X _14750_/Q _07077_/S vssd1 vssd1 vccd1 vccd1 _13596_/D sky130_fd_sc_hd__mux2_1
XFILLER_118_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput100 _07103_/X vssd1 vssd1 vccd1 vccd1 ext_write_strobe[1] sky130_fd_sc_hd__clkbuf_2
XFILLER_173_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07955_ _13553_/Q _07961_/C _13554_/Q vssd1 vssd1 vccd1 vccd1 _07955_/X sky130_fd_sc_hd__a21o_1
XFILLER_29_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06906_ _15380_/Q _06729_/Y _15379_/Q _06731_/Y _06905_/X vssd1 vssd1 vccd1 vccd1
+ _06906_/X sky130_fd_sc_hd__a221o_1
XFILLER_101_179 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_200 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07886_ _07886_/A vssd1 vssd1 vccd1 vccd1 _07886_/Y sky130_fd_sc_hd__inv_2
XFILLER_55_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09625_ _13999_/Q _13347_/A0 _09628_/S vssd1 vssd1 vccd1 vccd1 _13999_/D sky130_fd_sc_hd__mux2_1
XFILLER_56_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06837_ _08910_/S _06678_/Y _06834_/B _09382_/A _06836_/Y vssd1 vssd1 vccd1 vccd1
+ _06837_/X sky130_fd_sc_hd__o221a_1
XFILLER_56_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09556_ _15107_/Q _08497_/A _08508_/Y _13131_/A vssd1 vssd1 vccd1 vccd1 _09556_/X
+ sky130_fd_sc_hd__a31o_1
X_06768_ _15528_/Q vssd1 vssd1 vccd1 vccd1 _06768_/Y sky130_fd_sc_hd__inv_2
X_08507_ _08507_/A _09524_/A vssd1 vssd1 vccd1 vccd1 _08507_/Y sky130_fd_sc_hd__nor2_8
XFILLER_24_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06699_ _13472_/Q vssd1 vssd1 vccd1 vccd1 _06699_/Y sky130_fd_sc_hd__inv_2
X_09487_ _09554_/A _09487_/B _09487_/C vssd1 vssd1 vccd1 vccd1 _09487_/X sky130_fd_sc_hd__and3_1
XFILLER_178_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08438_ _13749_/Q _12878_/S _08426_/B _08437_/X vssd1 vssd1 vccd1 vccd1 _13749_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_169_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08369_ _08290_/X _11283_/B _11283_/A vssd1 vssd1 vccd1 vccd1 _08369_/X sky130_fd_sc_hd__mux2_2
XFILLER_149_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10400_ _08240_/A _13801_/Q _13769_/Q _08237_/A vssd1 vssd1 vccd1 vccd1 _10400_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_183_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11380_ _11380_/A _11389_/B vssd1 vssd1 vccd1 vccd1 _11383_/B sky130_fd_sc_hd__xnor2_2
XFILLER_164_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10331_ _14909_/Q _14716_/Q _10344_/S vssd1 vssd1 vccd1 vccd1 _14716_/D sky130_fd_sc_hd__mux2_1
X_13050_ _13050_/A _13050_/B _13050_/C vssd1 vssd1 vccd1 vccd1 _13051_/B sky130_fd_sc_hd__and3_1
X_10262_ _14647_/Q _14800_/Q _10735_/S vssd1 vssd1 vccd1 vccd1 _14647_/D sky130_fd_sc_hd__mux2_1
XFILLER_180_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12001_ _14459_/Q _14427_/Q _13848_/Q _14201_/Q _12407_/S _12406_/A vssd1 vssd1 vccd1
+ vccd1 _12001_/X sky130_fd_sc_hd__mux4_1
XFILLER_133_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10193_ _11879_/A1 _14577_/Q _10197_/S vssd1 vssd1 vccd1 vccd1 _14577_/D sky130_fd_sc_hd__mux2_1
XFILLER_160_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout382 _11349_/A vssd1 vssd1 vccd1 vccd1 _11259_/S sky130_fd_sc_hd__buf_12
X_13952_ _15315_/CLK _13952_/D vssd1 vssd1 vccd1 vccd1 _13952_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout393 _08230_/Y vssd1 vssd1 vccd1 vccd1 _11414_/A sky130_fd_sc_hd__buf_12
XFILLER_143_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12903_ _15431_/Q _15617_/Q _12904_/S vssd1 vssd1 vccd1 vccd1 _15431_/D sky130_fd_sc_hd__mux2_1
X_13883_ _15657_/CLK _13883_/D vssd1 vssd1 vccd1 vccd1 _13883_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_74_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_1014 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15622_ _15622_/CLK _15622_/D vssd1 vssd1 vccd1 vccd1 _15622_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12834_ _15074_/Q _12834_/B vssd1 vssd1 vccd1 vccd1 _12834_/X sky130_fd_sc_hd__or2_1
XFILLER_36_71 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15553_ _15553_/CLK _15553_/D vssd1 vssd1 vccd1 vccd1 _15553_/Q sky130_fd_sc_hd__dfxtp_1
X_12765_ _15357_/Q _12765_/B vssd1 vssd1 vccd1 vccd1 _12765_/X sky130_fd_sc_hd__or2_1
XTAP_2085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14504_ _15385_/CLK _14504_/D vssd1 vssd1 vccd1 vccd1 _14504_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11716_ _15145_/Q _11857_/A1 _11742_/S vssd1 vssd1 vccd1 vccd1 _15145_/D sky130_fd_sc_hd__mux2_1
XTAP_1384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15484_ _15499_/CLK _15484_/D vssd1 vssd1 vccd1 vccd1 _15484_/Q sky130_fd_sc_hd__dfxtp_1
X_12696_ _15055_/Q _12695_/X _12792_/B vssd1 vssd1 vccd1 vccd1 _12696_/X sky130_fd_sc_hd__mux2_1
XFILLER_175_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14435_ _15556_/CLK _14435_/D vssd1 vssd1 vccd1 vccd1 _14435_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11647_ _13322_/A0 _15079_/Q _11670_/S vssd1 vssd1 vccd1 vccd1 _15079_/D sky130_fd_sc_hd__mux2_1
Xinput13 ext_read_data[20] vssd1 vssd1 vccd1 vccd1 input13/X sky130_fd_sc_hd__clkbuf_4
XFILLER_30_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput24 ext_read_data[30] vssd1 vssd1 vccd1 vccd1 input24/X sky130_fd_sc_hd__clkbuf_16
XFILLER_128_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14366_ _15298_/CLK _14366_/D vssd1 vssd1 vccd1 vccd1 _14366_/Q sky130_fd_sc_hd__dfxtp_1
Xinput35 reset vssd1 vssd1 vccd1 vccd1 input35/X sky130_fd_sc_hd__buf_12
XFILLER_156_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11578_ _13226_/B _11572_/B _11577_/X vssd1 vssd1 vccd1 vccd1 _11578_/X sky130_fd_sc_hd__o21a_1
XFILLER_7_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_391 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_351 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13317_ _15648_/Q _10344_/S _10564_/A _15206_/Q vssd1 vssd1 vccd1 vccd1 _15648_/D
+ sky130_fd_sc_hd__a22o_1
X_10529_ _10529_/A _10529_/B vssd1 vssd1 vccd1 vccd1 _10558_/B sky130_fd_sc_hd__or2_2
XFILLER_6_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14297_ _15278_/CLK _14297_/D vssd1 vssd1 vccd1 vccd1 _14297_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_143_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13248_ _13242_/A _11349_/C _10530_/B vssd1 vssd1 vccd1 vccd1 _13248_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_112_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13179_ _15560_/Q _13252_/B _13177_/Y _13178_/Y vssd1 vssd1 vccd1 vccd1 _15560_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_35_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07740_ _07738_/Y _07746_/C _07750_/A vssd1 vssd1 vccd1 vccd1 _07740_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_111_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07671_ _13479_/Q _07672_/C _13480_/Q vssd1 vssd1 vccd1 vccd1 _07671_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_37_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09410_ _09421_/A1 _09406_/X _09409_/X _09405_/X vssd1 vssd1 vccd1 vccd1 _09411_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_179_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09341_ _14539_/Q _14152_/Q _14184_/Q _14120_/Q _09342_/S _09546_/S1 vssd1 vssd1
+ vccd1 vccd1 _09341_/X sky130_fd_sc_hd__mux4_1
XFILLER_33_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_978 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09272_ _14021_/Q _13989_/Q _09557_/S vssd1 vssd1 vccd1 vccd1 _09272_/X sky130_fd_sc_hd__mux2_1
XFILLER_178_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_488 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08223_ _14929_/D _14928_/D _14927_/D vssd1 vssd1 vccd1 vccd1 _08223_/X sky130_fd_sc_hd__or3b_4
XFILLER_20_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08154_ _08185_/A _08154_/B vssd1 vssd1 vccd1 vccd1 _08154_/X sky130_fd_sc_hd__and2_1
XFILLER_146_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07105_ _14900_/Q _07163_/A _07104_/X vssd1 vssd1 vccd1 vccd1 _07105_/X sky130_fd_sc_hd__a21o_4
XFILLER_147_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08085_ _15305_/Q _13647_/Q _08085_/S vssd1 vssd1 vccd1 vccd1 _08086_/B sky130_fd_sc_hd__mux2_1
XFILLER_119_599 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07036_ _14624_/Q _14656_/Q _07078_/S vssd1 vssd1 vccd1 vccd1 _07036_/X sky130_fd_sc_hd__mux2_1
XFILLER_161_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_399 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_742 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08987_ _15653_/Q _13387_/Q _09132_/S vssd1 vssd1 vccd1 vccd1 _08987_/X sky130_fd_sc_hd__mux2_1
XFILLER_87_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_4_5_0_clk clkbuf_4_5_0_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_5_0_clk/X sky130_fd_sc_hd__clkbuf_8
XFILLER_102_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07938_ _14742_/Q _08012_/A2 _07937_/Y _07938_/C1 vssd1 vssd1 vccd1 vccd1 _13549_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_69_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07869_ _13532_/Q _13531_/Q _13530_/Q _07869_/D vssd1 vssd1 vccd1 vccd1 _07884_/C
+ sky130_fd_sc_hd__and4_4
XFILLER_90_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09608_ _13982_/Q _13074_/B2 _09627_/S vssd1 vssd1 vccd1 vccd1 _13982_/D sky130_fd_sc_hd__mux2_1
XFILLER_16_439 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10880_ _14912_/Q _15543_/Q _13134_/A vssd1 vssd1 vccd1 vccd1 _14912_/D sky130_fd_sc_hd__mux2_1
XFILLER_113_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_208 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09539_ _12596_/A _09539_/B _09539_/C vssd1 vssd1 vccd1 vccd1 _09539_/X sky130_fd_sc_hd__and3_1
XFILLER_71_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1072 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_910 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12550_ _12573_/A _12550_/B _12550_/C vssd1 vssd1 vccd1 vccd1 _12550_/X sky130_fd_sc_hd__and3_1
XFILLER_12_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11501_ _11501_/A _11501_/B vssd1 vssd1 vccd1 vccd1 _11546_/A sky130_fd_sc_hd__and2_2
XFILLER_19_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_1048 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12481_ _12481_/A _12481_/B _12481_/C vssd1 vssd1 vccd1 vccd1 _12481_/X sky130_fd_sc_hd__and3_1
XFILLER_156_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14220_ _15518_/CLK _14220_/D vssd1 vssd1 vccd1 vccd1 _14220_/Q sky130_fd_sc_hd__dfxtp_1
X_11432_ _11432_/A _11441_/A vssd1 vssd1 vccd1 vccd1 _11460_/B sky130_fd_sc_hd__nor2_1
XFILLER_137_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14151_ _15096_/CLK _14151_/D vssd1 vssd1 vccd1 vccd1 _14151_/Q sky130_fd_sc_hd__dfxtp_1
X_11363_ _13162_/B _11363_/B _11363_/C vssd1 vssd1 vccd1 vccd1 _11363_/X sky130_fd_sc_hd__and3b_1
XFILLER_180_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13102_ _13020_/X _13104_/A2 _13104_/B1 _13344_/A0 vssd1 vssd1 vccd1 vccd1 _13102_/X
+ sky130_fd_sc_hd__a22o_1
X_10314_ _14699_/Q _14884_/Q _10695_/S vssd1 vssd1 vccd1 vccd1 _14699_/D sky130_fd_sc_hd__mux2_1
X_14082_ _15088_/CLK _14082_/D vssd1 vssd1 vccd1 vccd1 _14082_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11294_ _11294_/A _11294_/B vssd1 vssd1 vccd1 vccd1 _11294_/Y sky130_fd_sc_hd__nand2_1
XFILLER_152_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13033_ _13110_/B2 _13039_/A2 _13032_/X _12936_/X vssd1 vssd1 vccd1 vccd1 _13033_/X
+ sky130_fd_sc_hd__a22o_1
X_10245_ _14630_/Q _14783_/Q _10665_/S vssd1 vssd1 vccd1 vccd1 _14630_/D sky130_fd_sc_hd__mux2_1
XFILLER_152_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_1087 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10176_ _13329_/A0 _14560_/Q _10192_/S vssd1 vssd1 vccd1 vccd1 _14560_/D sky130_fd_sc_hd__mux2_1
XFILLER_79_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_1019 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14984_ _15582_/CLK _14984_/D vssd1 vssd1 vccd1 vccd1 _14984_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_93_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout190 _09997_/X vssd1 vssd1 vccd1 vccd1 _10029_/S sky130_fd_sc_hd__buf_12
X_13935_ _15326_/CLK _13935_/D vssd1 vssd1 vccd1 vccd1 _13935_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_35_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13866_ _15336_/CLK _13866_/D vssd1 vssd1 vccd1 vccd1 _13866_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15605_ _15638_/CLK _15605_/D vssd1 vssd1 vccd1 vccd1 _15605_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_179_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12817_ _15364_/Q _12759_/B _12816_/X _12832_/C1 vssd1 vssd1 vccd1 vccd1 _15364_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_37_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13797_ _15422_/CLK _13797_/D vssd1 vssd1 vccd1 vccd1 _13797_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15536_ _15536_/CLK _15536_/D vssd1 vssd1 vccd1 vccd1 _15536_/Q sky130_fd_sc_hd__dfxtp_1
X_12748_ _15062_/Q _12747_/Y _12792_/B vssd1 vssd1 vccd1 vccd1 _12748_/X sky130_fd_sc_hd__mux2_1
XTAP_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15467_ _15499_/CLK _15467_/D vssd1 vssd1 vccd1 vccd1 _15467_/Q sky130_fd_sc_hd__dfxtp_1
X_12679_ _15346_/Q _15345_/Q _12679_/C vssd1 vssd1 vccd1 vccd1 _12688_/B sky130_fd_sc_hd__and3_2
XFILLER_8_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14418_ _15677_/CLK _14418_/D vssd1 vssd1 vccd1 vccd1 _14418_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_163_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15398_ _15398_/CLK _15398_/D vssd1 vssd1 vccd1 vccd1 _15398_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_184_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14349_ _15286_/CLK _14349_/D vssd1 vssd1 vccd1 vccd1 _14349_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_156_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08910_ _13844_/Q _14197_/Q _08910_/S vssd1 vssd1 vccd1 vccd1 _08910_/X sky130_fd_sc_hd__mux2_1
XFILLER_98_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09890_ _11876_/A1 _14252_/Q _09892_/S vssd1 vssd1 vccd1 vccd1 _14252_/D sky130_fd_sc_hd__mux2_1
XFILLER_98_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08841_ _13864_/Q _11873_/A1 _08851_/S vssd1 vssd1 vccd1 vccd1 _13864_/D sky130_fd_sc_hd__mux2_1
XTAP_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08772_ _08772_/A _08772_/B _08779_/A _08771_/X vssd1 vssd1 vccd1 vccd1 _08772_/X
+ sky130_fd_sc_hd__or4b_2
XFILLER_111_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07723_ _13493_/Q _07724_/C _13494_/Q vssd1 vssd1 vccd1 vccd1 _07723_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_72_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07654_ _13476_/Q _13475_/Q _13474_/Q _13473_/Q vssd1 vssd1 vccd1 vccd1 _07655_/C
+ sky130_fd_sc_hd__and4_1
XFILLER_25_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_1075 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07585_ _07583_/Y _07587_/B _07607_/A vssd1 vssd1 vccd1 vccd1 _07585_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_81_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09324_ _13927_/Q _09323_/X _12573_/A vssd1 vssd1 vccd1 vccd1 _13927_/D sky130_fd_sc_hd__mux2_1
XFILLER_80_397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09255_ _09511_/S1 _08519_/B _09254_/X _08501_/A vssd1 vssd1 vccd1 vccd1 _09255_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_166_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08206_ _13697_/Q _13335_/A0 _08216_/S vssd1 vssd1 vccd1 vccd1 _13697_/D sky130_fd_sc_hd__mux2_1
X_09186_ _09419_/A2 _09184_/X _09185_/X _09421_/A1 _09183_/X vssd1 vssd1 vccd1 vccd1
+ _09186_/X sky130_fd_sc_hd__a221o_4
XFILLER_147_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08137_ input4/X input13/X _08150_/S vssd1 vssd1 vccd1 vccd1 _08137_/X sky130_fd_sc_hd__mux2_1
XFILLER_161_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08068_ _14761_/Q _13639_/Q _08072_/S vssd1 vssd1 vccd1 vccd1 _13639_/D sky130_fd_sc_hd__mux2_1
XFILLER_108_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07019_ _07018_/X _13585_/Q _12640_/S vssd1 vssd1 vccd1 vccd1 _07019_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10030_ _12832_/C1 _13580_/Q _08030_/Y _06997_/B _14388_/Q vssd1 vssd1 vccd1 vccd1
+ _14388_/D sky130_fd_sc_hd__a32o_1
XFILLER_49_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11981_ _11977_/X _11978_/X _12260_/A vssd1 vssd1 vccd1 vccd1 _11981_/X sky130_fd_sc_hd__mux2_1
XFILLER_1_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13720_ _14966_/CLK _13720_/D vssd1 vssd1 vccd1 vccd1 _13720_/Q sky130_fd_sc_hd__dfxtp_2
X_10932_ _14949_/Q _10931_/Y _10944_/B vssd1 vssd1 vccd1 vccd1 _14949_/D sky130_fd_sc_hd__mux2_1
XFILLER_56_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13651_ _15616_/CLK _13651_/D vssd1 vssd1 vccd1 vccd1 _13651_/Q sky130_fd_sc_hd__dfxtp_1
X_10863_ _14895_/Q hold1/X _10871_/S vssd1 vssd1 vccd1 vccd1 _14895_/D sky130_fd_sc_hd__mux2_1
XFILLER_44_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12602_ _12598_/X _12599_/X _12617_/S vssd1 vssd1 vccd1 vccd1 _12602_/X sky130_fd_sc_hd__mux2_1
XPHY_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13582_ _15618_/CLK _13582_/D vssd1 vssd1 vccd1 vccd1 _13582_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10794_ _14826_/Q _15458_/Q _12933_/S vssd1 vssd1 vccd1 vccd1 _14826_/D sky130_fd_sc_hd__mux2_1
XPHY_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15321_ _15664_/CLK _15321_/D vssd1 vssd1 vccd1 vccd1 _15321_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12533_ _12529_/X _12530_/X _12548_/S vssd1 vssd1 vccd1 vccd1 _12533_/X sky130_fd_sc_hd__mux2_1
XFILLER_157_425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15252_ _15284_/CLK _15252_/D vssd1 vssd1 vccd1 vccd1 _15252_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12464_ _12460_/X _12461_/X _12490_/A vssd1 vssd1 vccd1 vccd1 _12464_/X sky130_fd_sc_hd__mux2_1
XFILLER_149_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14203_ _15284_/CLK _14203_/D vssd1 vssd1 vccd1 vccd1 _14203_/Q sky130_fd_sc_hd__dfxtp_1
X_11415_ _11437_/A _11437_/B _13229_/A vssd1 vssd1 vccd1 vccd1 _11416_/B sky130_fd_sc_hd__a21oi_1
X_15183_ _15220_/CLK _15183_/D vssd1 vssd1 vccd1 vccd1 _15183_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12395_ _12391_/X _12392_/X _12594_/S vssd1 vssd1 vccd1 vccd1 _12395_/X sky130_fd_sc_hd__mux2_1
XFILLER_67_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14134_ _15202_/CLK _14134_/D vssd1 vssd1 vccd1 vccd1 _14134_/Q sky130_fd_sc_hd__dfxtp_1
X_11346_ _15041_/Q _11346_/A2 _11345_/X vssd1 vssd1 vccd1 vccd1 _15041_/D sky130_fd_sc_hd__a21o_1
XFILLER_4_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_152_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14065_ _14420_/CLK _14065_/D vssd1 vssd1 vccd1 vccd1 _14065_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_106_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11277_ _11283_/A _11344_/A _08282_/X _11346_/A2 vssd1 vssd1 vccd1 vccd1 _11277_/X
+ sky130_fd_sc_hd__a31o_1
X_13016_ _15485_/Q _13119_/S _13116_/C _13015_/X vssd1 vssd1 vccd1 vccd1 _15485_/D
+ sky130_fd_sc_hd__a22o_1
X_10228_ input24/X _14613_/Q _13291_/S vssd1 vssd1 vccd1 vccd1 _14613_/D sky130_fd_sc_hd__mux2_1
XFILLER_67_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2 hold2/A vssd1 vssd1 vccd1 vccd1 hold2/X sky130_fd_sc_hd__bufbuf_16
XFILLER_66_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10159_ _14544_/Q _13345_/A0 _10159_/S vssd1 vssd1 vccd1 vccd1 _14544_/D sky130_fd_sc_hd__mux2_1
XFILLER_181_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14967_ _15000_/CLK _14967_/D vssd1 vssd1 vccd1 vccd1 _14967_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13918_ _15507_/CLK _13918_/D vssd1 vssd1 vccd1 vccd1 _13918_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14898_ _15616_/CLK _14898_/D vssd1 vssd1 vccd1 vccd1 _14898_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_74_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13849_ _14462_/CLK _13849_/D vssd1 vssd1 vccd1 vccd1 _13849_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_386 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07370_ _14714_/Q _14715_/Q _13318_/C _11710_/A vssd1 vssd1 vccd1 vccd1 _07370_/X
+ sky130_fd_sc_hd__or4_4
XFILLER_188_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_572 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15519_ _15519_/CLK _15519_/D vssd1 vssd1 vccd1 vccd1 _15519_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_175_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09040_ _09445_/C1 _09039_/X _09038_/X _09130_/A vssd1 vssd1 vccd1 vccd1 _09040_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_129_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09942_ _13072_/B2 _14302_/Q _09958_/S vssd1 vssd1 vccd1 vccd1 _14302_/D sky130_fd_sc_hd__mux2_1
XFILLER_132_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09873_ _12967_/A1 _14235_/Q _09892_/S vssd1 vssd1 vccd1 vccd1 _14235_/D sky130_fd_sc_hd__mux2_1
XTAP_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08824_ _13847_/Q _13323_/A0 _08846_/S vssd1 vssd1 vccd1 vccd1 _13847_/D sky130_fd_sc_hd__mux2_1
XTAP_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08755_ _08754_/A _08765_/A _08753_/X _08754_/Y vssd1 vssd1 vccd1 vccd1 _08755_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_2607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07706_ _07713_/A _07706_/B vssd1 vssd1 vccd1 vccd1 _07706_/Y sky130_fd_sc_hd__nand2_1
XTAP_2618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08686_ _15377_/Q _08690_/A2 _08690_/B1 _13422_/Q vssd1 vssd1 vccd1 vccd1 _08686_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_81_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07637_ _14760_/Q _07651_/A _07636_/Y _08012_/C1 vssd1 vssd1 vccd1 vccd1 _13471_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_54_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07568_ _07629_/A _07568_/B vssd1 vssd1 vccd1 vccd1 _07568_/Y sky130_fd_sc_hd__nand2_1
XFILLER_179_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09307_ _08507_/A _09304_/X _09306_/X _09554_/A vssd1 vssd1 vccd1 vccd1 _09307_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_142_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07499_ _13680_/Q _07499_/A2 _07499_/B1 _14708_/Q _07498_/X vssd1 vssd1 vccd1 vccd1
+ _07499_/X sky130_fd_sc_hd__a221o_1
XFILLER_186_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09238_ _13923_/Q _09237_/X _12596_/A vssd1 vssd1 vccd1 vccd1 _13923_/D sky130_fd_sc_hd__mux2_1
XFILLER_148_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09169_ _14016_/Q _13984_/Q _09441_/S vssd1 vssd1 vccd1 vccd1 _09169_/X sky130_fd_sc_hd__mux2_1
XFILLER_5_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11200_ _14992_/Q _11202_/A _11170_/X _11199_/Y vssd1 vssd1 vccd1 vccd1 _14992_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_163_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12180_ _12163_/X _12164_/X _12502_/S vssd1 vssd1 vccd1 vccd1 _12180_/X sky130_fd_sc_hd__mux2_1
XFILLER_134_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11131_ _11199_/A _11187_/B vssd1 vssd1 vccd1 vccd1 _11131_/Y sky130_fd_sc_hd__nand2_1
XFILLER_150_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11062_ _11059_/X _11061_/A _11252_/A vssd1 vssd1 vccd1 vccd1 _11062_/X sky130_fd_sc_hd__mux2_1
XFILLER_1_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_74 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10013_ _13334_/A0 _14371_/Q _10028_/S vssd1 vssd1 vccd1 vccd1 _14371_/D sky130_fd_sc_hd__mux2_1
XFILLER_62_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_1079 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14821_ _15641_/CLK _14821_/D vssd1 vssd1 vccd1 vccd1 _14821_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14752_ _15452_/CLK _14752_/D vssd1 vssd1 vccd1 vccd1 _14752_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_151_62 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11964_ _13942_/Q _13684_/Q _12079_/S vssd1 vssd1 vccd1 vccd1 _11965_/B sky130_fd_sc_hd__mux2_1
XTAP_3875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13703_ _15651_/CLK _13703_/D vssd1 vssd1 vccd1 vccd1 _13703_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10915_ _14940_/Q _10944_/B _10914_/Y _11440_/A vssd1 vssd1 vccd1 vccd1 _14940_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_60_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14683_ _14892_/CLK _14683_/D vssd1 vssd1 vccd1 vccd1 _14683_/Q sky130_fd_sc_hd__dfxtp_1
X_11895_ _13939_/Q _13681_/Q _12269_/S vssd1 vssd1 vccd1 vccd1 _11896_/B sky130_fd_sc_hd__mux2_1
X_13634_ _14510_/CLK _13634_/D vssd1 vssd1 vccd1 vccd1 _13634_/Q sky130_fd_sc_hd__dfxtp_1
X_10846_ _14878_/Q _13790_/Q _12927_/S vssd1 vssd1 vccd1 vccd1 _14878_/D sky130_fd_sc_hd__mux2_1
XFILLER_158_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_740 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13565_ _13565_/CLK _13565_/D vssd1 vssd1 vccd1 vccd1 _13565_/Q sky130_fd_sc_hd__dfxtp_1
X_10777_ _14809_/Q _15441_/Q _12918_/S vssd1 vssd1 vccd1 vccd1 _14809_/D sky130_fd_sc_hd__mux2_1
XFILLER_157_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15304_ _15304_/CLK _15304_/D vssd1 vssd1 vccd1 vccd1 _15304_/Q sky130_fd_sc_hd__dfxtp_1
X_12516_ _13966_/Q _13708_/Q _12522_/S vssd1 vssd1 vccd1 vccd1 _12517_/B sky130_fd_sc_hd__mux2_1
X_13496_ _13632_/CLK _13496_/D vssd1 vssd1 vccd1 vccd1 _13496_/Q sky130_fd_sc_hd__dfxtp_1
X_15235_ _15235_/CLK _15235_/D vssd1 vssd1 vccd1 vccd1 _15235_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_157_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12447_ _13963_/Q _13705_/Q _12453_/S vssd1 vssd1 vccd1 vccd1 _12448_/B sky130_fd_sc_hd__mux2_1
X_15166_ _15235_/CLK _15166_/D vssd1 vssd1 vccd1 vccd1 _15166_/Q sky130_fd_sc_hd__dfxtp_1
X_12378_ _13960_/Q _13702_/Q _12518_/S vssd1 vssd1 vccd1 vccd1 _12379_/B sky130_fd_sc_hd__mux2_1
XFILLER_99_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14117_ _14439_/CLK _14117_/D vssd1 vssd1 vccd1 vccd1 _14117_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11329_ _11329_/A _11329_/B vssd1 vssd1 vccd1 vccd1 _11329_/Y sky130_fd_sc_hd__nor2_1
XFILLER_140_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15097_ _15544_/CLK _15097_/D vssd1 vssd1 vccd1 vccd1 _15097_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14048_ _15331_/CLK _14048_/D vssd1 vssd1 vccd1 vccd1 _14048_/Q sky130_fd_sc_hd__dfxtp_1
X_06870_ _06700_/Y _13503_/Q _14511_/Q _06703_/Y vssd1 vssd1 vccd1 vccd1 _06871_/B
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_83_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08540_ _08724_/C _08540_/B vssd1 vssd1 vccd1 vccd1 _08540_/X sky130_fd_sc_hd__and2_4
XFILLER_54_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08471_ _13764_/Q _10764_/S _08470_/X _14613_/Q vssd1 vssd1 vccd1 vccd1 _13764_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_39_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07422_ _14657_/Q _07474_/B _07482_/C vssd1 vssd1 vccd1 vccd1 _07422_/X sky130_fd_sc_hd__and3_1
XFILLER_165_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07353_ _07347_/X _07363_/B _07352_/Y _07311_/X _07278_/X vssd1 vssd1 vccd1 vccd1
+ _07353_/X sky130_fd_sc_hd__o32a_1
XFILLER_176_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_929 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07284_ _07284_/A vssd1 vssd1 vccd1 vccd1 _07287_/A sky130_fd_sc_hd__inv_2
XFILLER_148_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09023_ _14460_/Q _09536_/A2 _09022_/X _06676_/A vssd1 vssd1 vccd1 vccd1 _09023_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_40_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09925_ _13104_/B2 _14286_/Q _09925_/S vssd1 vssd1 vccd1 vccd1 _14286_/D sky130_fd_sc_hd__mux2_1
XFILLER_160_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09856_ _14220_/Q _13343_/A0 _09858_/S vssd1 vssd1 vccd1 vccd1 _14220_/D sky130_fd_sc_hd__mux2_1
XFILLER_59_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08807_ _11874_/A1 _13833_/Q _08816_/S vssd1 vssd1 vccd1 vccd1 _13833_/D sky130_fd_sc_hd__mux2_1
XFILLER_65_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09787_ _14154_/Q _13342_/A0 _09795_/S vssd1 vssd1 vccd1 vccd1 _14154_/D sky130_fd_sc_hd__mux2_1
XTAP_3127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06999_ _14722_/Q _14721_/Q _14723_/Q vssd1 vssd1 vccd1 vccd1 _10098_/A sky130_fd_sc_hd__or3b_4
XTAP_3138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08738_ _13614_/Q _08750_/B1 _08737_/X _13154_/S vssd1 vssd1 vccd1 vccd1 _08738_/X
+ sky130_fd_sc_hd__a211o_1
XANTENNA_105 _14750_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_116 _07184_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_127 _08453_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08669_ _13456_/Q _08684_/A2 _08685_/A2 _13552_/Q vssd1 vssd1 vccd1 vccd1 _08669_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_42_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10700_ _14758_/Q _10699_/X _10710_/S vssd1 vssd1 vccd1 vccd1 _14758_/D sky130_fd_sc_hd__mux2_1
XFILLER_14_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_492 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11680_ _11680_/A0 _15111_/Q _11703_/S vssd1 vssd1 vccd1 vccd1 _15111_/D sky130_fd_sc_hd__mux2_1
XTAP_1769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_98 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10631_ _15005_/Q _10717_/A2 _10722_/B1 _14941_/Q _10717_/C1 vssd1 vssd1 vccd1 vccd1
+ _10631_/X sky130_fd_sc_hd__a221o_1
XFILLER_179_380 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_63 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13350_ _13350_/A0 _15680_/Q _13350_/S vssd1 vssd1 vccd1 vccd1 _15680_/D sky130_fd_sc_hd__mux2_1
XFILLER_139_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10562_ _14924_/Q _06857_/C _07115_/B _10730_/S vssd1 vssd1 vccd1 vccd1 _10563_/B
+ sky130_fd_sc_hd__o31a_2
XFILLER_167_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12301_ _14536_/Q _14149_/Q _14181_/Q _14117_/Q _12612_/S _12383_/A vssd1 vssd1 vccd1
+ vccd1 _12301_/X sky130_fd_sc_hd__mux4_1
XFILLER_127_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13281_ _15365_/Q _15612_/Q _13282_/S vssd1 vssd1 vccd1 vccd1 _15612_/D sky130_fd_sc_hd__mux2_1
X_10493_ _07256_/X _08225_/Y _10492_/X vssd1 vssd1 vccd1 vccd1 _11536_/B sky130_fd_sc_hd__a21oi_4
X_15020_ _15020_/CLK _15020_/D vssd1 vssd1 vccd1 vccd1 _15020_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12232_ _14533_/Q _14146_/Q _14178_/Q _14114_/Q _12499_/S _12489_/S1 vssd1 vssd1
+ vccd1 vccd1 _12232_/X sky130_fd_sc_hd__mux4_1
XFILLER_182_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12163_ _14530_/Q _14143_/Q _14175_/Q _14111_/Q _12246_/S _12452_/A vssd1 vssd1 vccd1
+ vccd1 _12163_/X sky130_fd_sc_hd__mux4_1
XFILLER_162_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11114_ _11112_/X _11113_/X _11371_/A vssd1 vssd1 vccd1 vccd1 _11114_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12094_ _14527_/Q _14140_/Q _14172_/Q _14108_/Q _12476_/S _12498_/A vssd1 vssd1 vccd1
+ vccd1 _12094_/X sky130_fd_sc_hd__mux4_1
XFILLER_110_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11045_ _11045_/A _11045_/B vssd1 vssd1 vccd1 vccd1 _11045_/Y sky130_fd_sc_hd__nor2_1
XFILLER_39_71 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14804_ _15612_/CLK _14804_/D vssd1 vssd1 vccd1 vccd1 _14804_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12996_ _10664_/X _14879_/Q _13038_/S vssd1 vssd1 vccd1 vccd1 _12996_/X sky130_fd_sc_hd__mux2_8
XTAP_3661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11947_ _14069_/Q _14037_/Q _12407_/S vssd1 vssd1 vccd1 vccd1 _11947_/X sky130_fd_sc_hd__mux2_1
XFILLER_45_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14735_ _15616_/CLK _14735_/D vssd1 vssd1 vccd1 vccd1 _14735_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_3694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14666_ _15375_/CLK _14666_/D vssd1 vssd1 vccd1 vccd1 _14666_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11878_ _15299_/Q _13345_/A0 _11878_/S vssd1 vssd1 vccd1 vccd1 _15299_/D sky130_fd_sc_hd__mux2_1
X_13617_ _15374_/CLK _13617_/D vssd1 vssd1 vccd1 vccd1 _13617_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10829_ _14861_/Q _07197_/A _12906_/S vssd1 vssd1 vccd1 vccd1 _14861_/D sky130_fd_sc_hd__mux2_1
X_14597_ _14892_/CLK _14597_/D vssd1 vssd1 vccd1 vccd1 _14597_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_186_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13548_ _13798_/CLK _13548_/D vssd1 vssd1 vccd1 vccd1 _13548_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_158_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13479_ _14517_/CLK _13479_/D vssd1 vssd1 vccd1 vccd1 _13479_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_65_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15218_ _15218_/CLK _15218_/D vssd1 vssd1 vccd1 vccd1 _15218_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_962 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15149_ _15218_/CLK _15149_/D vssd1 vssd1 vccd1 vccd1 _15149_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_290 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07971_ _07971_/A _07971_/B vssd1 vssd1 vccd1 vccd1 _07971_/Y sky130_fd_sc_hd__nand2_1
XFILLER_113_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09710_ _13078_/B2 _14080_/Q _09723_/S vssd1 vssd1 vccd1 vccd1 _14080_/D sky130_fd_sc_hd__mux2_1
X_06922_ _06922_/A _06922_/B _06922_/C vssd1 vssd1 vccd1 vccd1 _06923_/C sky130_fd_sc_hd__or3_1
XFILLER_45_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09641_ _14014_/Q _13074_/B2 _09660_/S vssd1 vssd1 vccd1 vccd1 _14014_/D sky130_fd_sc_hd__mux2_1
X_06853_ _13309_/A vssd1 vssd1 vccd1 vccd1 _13316_/S sky130_fd_sc_hd__inv_8
XFILLER_68_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09572_ _13948_/Q _13328_/A0 _09589_/S vssd1 vssd1 vccd1 vccd1 _13948_/D sky130_fd_sc_hd__mux2_1
XFILLER_71_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06784_ _14587_/Q _06987_/D _14589_/Q _14588_/Q vssd1 vssd1 vccd1 vccd1 _08469_/A
+ sky130_fd_sc_hd__and4b_4
XFILLER_35_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08523_ _08529_/B _08532_/B vssd1 vssd1 vccd1 vccd1 _08523_/Y sky130_fd_sc_hd__nor2_4
XFILLER_24_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08454_ _13757_/Q _12878_/S _08426_/X _08453_/X vssd1 vssd1 vccd1 vccd1 _13757_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_23_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07405_ _13326_/A0 _13390_/Q _07481_/S vssd1 vssd1 vccd1 vccd1 _13390_/D sky130_fd_sc_hd__mux2_1
XFILLER_168_339 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08385_ _11025_/A _13202_/B _11036_/B vssd1 vssd1 vccd1 vccd1 _08385_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_149_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07336_ _07336_/A vssd1 vssd1 vccd1 vccd1 _07337_/B sky130_fd_sc_hd__inv_2
XFILLER_167_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07267_ _07237_/Y _07238_/X _07242_/X _07244_/Y vssd1 vssd1 vccd1 vccd1 _07268_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_09006_ _14072_/Q _09522_/A2 _09519_/B1 _14040_/Q _09532_/A vssd1 vssd1 vccd1 vccd1
+ _09006_/X sky130_fd_sc_hd__a221o_1
XFILLER_136_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07198_ _06768_/Y _07197_/X _15529_/Q vssd1 vssd1 vccd1 vccd1 _07365_/A sky130_fd_sc_hd__a21bo_1
XFILLER_183_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout520 _09435_/A vssd1 vssd1 vccd1 vccd1 _09391_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_104_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout531 _08487_/A vssd1 vssd1 vccd1 vccd1 _09530_/S1 sky130_fd_sc_hd__clkbuf_16
XFILLER_116_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout542 _08487_/A vssd1 vssd1 vccd1 vccd1 _08508_/B sky130_fd_sc_hd__buf_12
X_09908_ _11861_/A1 _14269_/Q _09925_/S vssd1 vssd1 vccd1 vccd1 _14269_/D sky130_fd_sc_hd__mux2_1
Xfanout553 _09438_/S0 vssd1 vssd1 vccd1 vccd1 _09441_/S sky130_fd_sc_hd__buf_6
Xfanout564 _08910_/S vssd1 vssd1 vccd1 vccd1 _09342_/S sky130_fd_sc_hd__buf_8
XFILLER_58_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout575 _14601_/Q vssd1 vssd1 vccd1 vccd1 _08405_/C sky130_fd_sc_hd__buf_12
Xfanout586 _12061_/A vssd1 vssd1 vccd1 vccd1 _12268_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_58_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout597 fanout600/X vssd1 vssd1 vccd1 vccd1 _12540_/A sky130_fd_sc_hd__buf_4
X_09839_ _14203_/Q _12967_/A1 _09858_/S vssd1 vssd1 vccd1 vccd1 _14203_/D sky130_fd_sc_hd__mux2_1
XFILLER_47_938 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12850_ _14744_/Q _15378_/Q _12866_/S vssd1 vssd1 vccd1 vccd1 _15378_/D sky130_fd_sc_hd__mux2_1
XFILLER_74_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11801_ _15224_/Q _13082_/B2 _11816_/S vssd1 vssd1 vccd1 vccd1 _15224_/D sky130_fd_sc_hd__mux2_1
XFILLER_73_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12781_ _06861_/Y _12778_/X _12779_/X _12780_/X vssd1 vssd1 vccd1 vccd1 _12781_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_27_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14520_ _15211_/CLK _14520_/D vssd1 vssd1 vccd1 vccd1 _14520_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11732_ _15161_/Q _13340_/A0 _11742_/S vssd1 vssd1 vccd1 vccd1 _15161_/D sky130_fd_sc_hd__mux2_1
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1046 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14451_ _15650_/CLK _14451_/D vssd1 vssd1 vccd1 vccd1 _14451_/Q sky130_fd_sc_hd__dfxtp_1
X_11663_ _13338_/A0 _15095_/Q _11675_/S vssd1 vssd1 vccd1 vccd1 _15095_/D sky130_fd_sc_hd__mux2_1
XFILLER_30_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13402_ _15668_/CLK _13402_/D vssd1 vssd1 vccd1 vccd1 _13402_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_174_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10614_ _15050_/Q _10734_/A2 _10611_/X _10613_/X vssd1 vssd1 vccd1 vccd1 _10614_/X
+ sky130_fd_sc_hd__o22a_1
X_14382_ _15267_/CLK _14382_/D vssd1 vssd1 vccd1 vccd1 _14382_/Q sky130_fd_sc_hd__dfxtp_1
X_11594_ _11606_/A _11604_/A vssd1 vssd1 vccd1 vccd1 _11596_/A sky130_fd_sc_hd__nor2_1
XFILLER_168_895 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13333_ _13333_/A0 _15663_/Q _13345_/S vssd1 vssd1 vccd1 vccd1 _15663_/D sky130_fd_sc_hd__mux2_1
X_10545_ _10365_/B _10417_/X _10418_/Y _10558_/B vssd1 vssd1 vccd1 vccd1 _10545_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_6_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_130_clk clkbuf_5_30_0_clk/X vssd1 vssd1 vccd1 vccd1 _15393_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_6_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13264_ _15348_/Q _15595_/Q _13300_/S vssd1 vssd1 vccd1 vccd1 _15595_/D sky130_fd_sc_hd__mux2_1
X_10476_ _11589_/B _13226_/B vssd1 vssd1 vccd1 vccd1 _10478_/A sky130_fd_sc_hd__nand2_1
XFILLER_143_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15003_ _15006_/CLK _15003_/D vssd1 vssd1 vccd1 vccd1 _15003_/Q sky130_fd_sc_hd__dfxtp_1
X_12215_ _08453_/A _12212_/X _08451_/A vssd1 vssd1 vccd1 vccd1 _12215_/X sky130_fd_sc_hd__o21a_1
XFILLER_108_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13195_ _13217_/A _13195_/B vssd1 vssd1 vccd1 vccd1 _13195_/Y sky130_fd_sc_hd__nand2_1
XFILLER_155_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12146_ _12500_/B1 _12143_/X _12501_/C1 vssd1 vssd1 vccd1 vccd1 _12146_/X sky130_fd_sc_hd__o21a_1
XFILLER_150_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12077_ _12468_/A1 _12074_/X _12455_/C1 vssd1 vssd1 vccd1 vccd1 _12077_/X sky130_fd_sc_hd__o21a_1
XFILLER_1_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11028_ _11024_/X _11027_/X _11259_/S vssd1 vssd1 vccd1 vccd1 _11029_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_197_clk clkbuf_5_17_0_clk/X vssd1 vssd1 vccd1 vccd1 _15651_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_2_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12979_ _13074_/B2 _13024_/A2 _12978_/X _13024_/B2 vssd1 vssd1 vccd1 vccd1 _12979_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_3491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14718_ _15542_/CLK _14718_/D vssd1 vssd1 vccd1 vccd1 _14718_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_33_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_177_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14649_ _14649_/CLK _14649_/D vssd1 vssd1 vccd1 vccd1 _14649_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_16 _15054_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_27 _14746_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08170_ _13672_/Q _10285_/S _08155_/X _08169_/X vssd1 vssd1 vccd1 vccd1 _13672_/D
+ sky130_fd_sc_hd__o22a_1
XANTENNA_38 input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_49 _07177_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07121_ _07131_/A _07121_/B vssd1 vssd1 vccd1 vccd1 _07121_/X sky130_fd_sc_hd__and2_2
Xclkbuf_leaf_121_clk clkbuf_5_30_0_clk/X vssd1 vssd1 vccd1 vccd1 _15383_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_119_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07052_ _07051_/X _13596_/Q _12728_/S vssd1 vssd1 vccd1 vccd1 _07052_/X sky130_fd_sc_hd__mux2_1
XFILLER_146_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput101 _07105_/X vssd1 vssd1 vccd1 vccd1 ext_write_strobe[2] sky130_fd_sc_hd__clkbuf_2
XFILLER_161_526 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_442 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07954_ _07961_/C _07961_/D vssd1 vssd1 vccd1 vccd1 _07958_/B sky130_fd_sc_hd__nand2_1
X_06905_ _15379_/Q _06731_/Y _15378_/Q _06733_/Y _06904_/X vssd1 vssd1 vccd1 vccd1
+ _06905_/X sky130_fd_sc_hd__o221a_1
XFILLER_101_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07885_ _13535_/Q _07884_/C _07884_/D _13536_/Q vssd1 vssd1 vccd1 vccd1 _07886_/A
+ sky130_fd_sc_hd__a31o_1
Xclkbuf_leaf_188_clk clkbuf_5_21_0_clk/X vssd1 vssd1 vccd1 vccd1 _15192_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_55_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09624_ _13998_/Q _13346_/A0 _09628_/S vssd1 vssd1 vccd1 vccd1 _13998_/D sky130_fd_sc_hd__mux2_1
XFILLER_56_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06836_ _09466_/A _14907_/Q vssd1 vssd1 vccd1 vccd1 _06836_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_55_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09555_ _14549_/Q _14162_/Q _14194_/Q _14130_/Q _09557_/S _13144_/A0 vssd1 vssd1
+ vccd1 vccd1 _09555_/X sky130_fd_sc_hd__mux4_1
X_06767_ _14928_/Q vssd1 vssd1 vccd1 vccd1 _10581_/B sky130_fd_sc_hd__inv_2
XFILLER_70_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08506_ _08517_/A _13127_/C vssd1 vssd1 vccd1 vccd1 _08724_/C sky130_fd_sc_hd__nor2_4
X_09486_ _09550_/A1 _09484_/X _09485_/X vssd1 vssd1 vccd1 vccd1 _09487_/C sky130_fd_sc_hd__a21o_1
X_06698_ _13504_/Q vssd1 vssd1 vccd1 vccd1 _06698_/Y sky130_fd_sc_hd__inv_2
XFILLER_23_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08437_ _14608_/Q _08390_/C _08425_/X _10764_/S vssd1 vssd1 vccd1 vccd1 _08437_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_23_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08368_ _08329_/X _08367_/X _11297_/S vssd1 vssd1 vccd1 vccd1 _11283_/B sky130_fd_sc_hd__mux2_1
XFILLER_108_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07319_ _13912_/Q _15499_/Q _07334_/S vssd1 vssd1 vccd1 vccd1 _07319_/X sky130_fd_sc_hd__mux2_8
XFILLER_109_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08299_ _11329_/A _08299_/B _08299_/C vssd1 vssd1 vccd1 vccd1 _08299_/X sky130_fd_sc_hd__and3_1
XFILLER_20_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_165_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10330_ _14908_/Q _14715_/Q _10566_/B vssd1 vssd1 vccd1 vccd1 _14715_/D sky130_fd_sc_hd__mux2_1
XFILLER_125_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10261_ _14646_/Q _14799_/Q _10730_/S vssd1 vssd1 vccd1 vccd1 _14646_/D sky130_fd_sc_hd__mux2_1
XFILLER_133_740 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12000_ _14233_/Q _14265_/Q _14297_/Q _14329_/Q _12407_/S _12406_/A vssd1 vssd1 vccd1
+ vccd1 _12000_/X sky130_fd_sc_hd__mux4_1
Xclkbuf_5_14_0_clk clkbuf_4_7_0_clk/X vssd1 vssd1 vccd1 vccd1 clkbuf_5_14_0_clk/X
+ sky130_fd_sc_hd__clkbuf_8
X_10192_ _13345_/A0 _14576_/Q _10192_/S vssd1 vssd1 vccd1 vccd1 _14576_/D sky130_fd_sc_hd__mux2_1
XFILLER_120_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout350 _12834_/B vssd1 vssd1 vccd1 vccd1 _12792_/B sky130_fd_sc_hd__buf_12
Xfanout361 _08519_/X vssd1 vssd1 vccd1 vccd1 _08520_/B sky130_fd_sc_hd__buf_12
XFILLER_143_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout372 _11013_/A vssd1 vssd1 vccd1 vccd1 _11037_/A sky130_fd_sc_hd__buf_6
Xclkbuf_leaf_179_clk clkbuf_5_22_0_clk/X vssd1 vssd1 vccd1 vccd1 _15667_/CLK sky130_fd_sc_hd__clkbuf_16
X_13951_ _15233_/CLK _13951_/D vssd1 vssd1 vccd1 vccd1 _13951_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout383 _08238_/Y vssd1 vssd1 vccd1 vccd1 _11349_/A sky130_fd_sc_hd__buf_6
XFILLER_101_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout394 _11371_/A vssd1 vssd1 vccd1 vccd1 _11347_/A sky130_fd_sc_hd__buf_8
XFILLER_19_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_143_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12902_ _15430_/Q _15616_/Q _12906_/S vssd1 vssd1 vccd1 vccd1 _15430_/D sky130_fd_sc_hd__mux2_1
Xclkbuf_5_29_0_clk clkbuf_5_29_0_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_5_29_0_clk/X
+ sky130_fd_sc_hd__clkbuf_8
X_13882_ _15656_/CLK _13882_/D vssd1 vssd1 vccd1 vccd1 _13882_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_919 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_1026 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15621_ _15646_/CLK _15621_/D vssd1 vssd1 vccd1 vccd1 _15621_/Q sky130_fd_sc_hd__dfxtp_1
X_12833_ _15367_/Q _12833_/B vssd1 vssd1 vccd1 vccd1 _12833_/Y sky130_fd_sc_hd__xnor2_1
XTAP_2031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12764_ _13434_/Q _12763_/X _12764_/S vssd1 vssd1 vccd1 vccd1 _12764_/X sky130_fd_sc_hd__mux2_1
XFILLER_14_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15552_ _15552_/CLK _15552_/D vssd1 vssd1 vccd1 vccd1 _15552_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14503_ _15386_/CLK _14503_/D vssd1 vssd1 vccd1 vccd1 _14503_/Q sky130_fd_sc_hd__dfxtp_1
X_11715_ _15144_/Q _13323_/A0 _11741_/S vssd1 vssd1 vccd1 vccd1 _15144_/D sky130_fd_sc_hd__mux2_1
XFILLER_159_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15483_ _15489_/CLK _15483_/D vssd1 vssd1 vccd1 vccd1 _15483_/Q sky130_fd_sc_hd__dfxtp_1
X_12695_ _15348_/Q _12701_/C vssd1 vssd1 vccd1 vccd1 _12695_/X sky130_fd_sc_hd__xor2_2
XFILLER_159_136 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_495 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14434_ _15285_/CLK _14434_/D vssd1 vssd1 vccd1 vccd1 _14434_/Q sky130_fd_sc_hd__dfxtp_1
X_11646_ _13321_/A0 _15078_/Q _11675_/S vssd1 vssd1 vccd1 vccd1 _15078_/D sky130_fd_sc_hd__mux2_1
XFILLER_156_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput14 ext_read_data[21] vssd1 vssd1 vccd1 vccd1 input14/X sky130_fd_sc_hd__buf_4
Xinput25 ext_read_data[31] vssd1 vssd1 vccd1 vccd1 input25/X sky130_fd_sc_hd__buf_6
XFILLER_174_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14365_ _15218_/CLK _14365_/D vssd1 vssd1 vccd1 vccd1 _14365_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_183_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11577_ _13226_/B _11572_/B _11564_/A vssd1 vssd1 vccd1 vccd1 _11577_/X sky130_fd_sc_hd__a21bo_1
Xclkbuf_leaf_103_clk clkbuf_5_26_0_clk/X vssd1 vssd1 vccd1 vccd1 _15624_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_116_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13316_ _15647_/Q _12833_/Y _13316_/S vssd1 vssd1 vccd1 vccd1 _15647_/D sky130_fd_sc_hd__mux2_1
XFILLER_183_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10528_ _10528_/A _10528_/B _10528_/C _10528_/D vssd1 vssd1 vccd1 vccd1 _10529_/B
+ sky130_fd_sc_hd__or4_1
XFILLER_155_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14296_ _15284_/CLK _14296_/D vssd1 vssd1 vccd1 vccd1 _14296_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_526 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13247_ _15582_/Q _13214_/B _13245_/X _13246_/Y vssd1 vssd1 vccd1 vccd1 _15582_/D
+ sky130_fd_sc_hd__a22o_1
X_10459_ _07215_/A _10481_/B _10458_/X vssd1 vssd1 vccd1 vccd1 wire360/A sky130_fd_sc_hd__a21oi_2
X_13178_ _13242_/A _13178_/B vssd1 vssd1 vccd1 vccd1 _13178_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_69_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12129_ _14013_/Q _13981_/Q _12476_/S vssd1 vssd1 vccd1 vccd1 _12130_/B sky130_fd_sc_hd__mux2_1
XFILLER_112_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_990 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07670_ _14736_/Q _07777_/A _07669_/Y _08016_/C1 vssd1 vssd1 vccd1 vccd1 _13479_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_92_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09340_ _09382_/A _09340_/B _09340_/C vssd1 vssd1 vccd1 vccd1 _09340_/X sky130_fd_sc_hd__and3_1
XFILLER_34_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09271_ _09550_/A1 _09269_/X _09270_/X vssd1 vssd1 vccd1 vccd1 _09275_/B sky130_fd_sc_hd__a21o_1
XFILLER_21_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08222_ _14929_/D _14928_/D _14927_/D vssd1 vssd1 vccd1 vccd1 wire438/A sky130_fd_sc_hd__nor3b_4
XFILLER_138_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08153_ _13664_/Q _10710_/S _08152_/X vssd1 vssd1 vccd1 vccd1 _13664_/D sky130_fd_sc_hd__o21a_1
XFILLER_147_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07104_ _07146_/S _07163_/A _07104_/C vssd1 vssd1 vccd1 vccd1 _07104_/X sky130_fd_sc_hd__and3b_4
XFILLER_180_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08084_ _14736_/Q _08083_/A _08083_/Y _08084_/C1 vssd1 vssd1 vccd1 vccd1 _13646_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_134_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07035_ _07034_/X _14744_/Q _07077_/S vssd1 vssd1 vccd1 vccd1 _13590_/D sky130_fd_sc_hd__mux2_1
XFILLER_164_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08986_ _14522_/Q _14135_/Q _14167_/Q _14103_/Q _09132_/S _08988_/A1 vssd1 vssd1
+ vccd1 vccd1 _08986_/X sky130_fd_sc_hd__mux4_1
XFILLER_88_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07937_ _07946_/D _07936_/Y _08012_/A2 vssd1 vssd1 vccd1 vccd1 _07937_/Y sky130_fd_sc_hd__o21ai_1
X_07868_ _14756_/Q _07874_/A _07867_/Y vssd1 vssd1 vccd1 vccd1 _13531_/D sky130_fd_sc_hd__o21a_1
XFILLER_56_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09607_ _13981_/Q _13072_/B2 _09627_/S vssd1 vssd1 vccd1 vccd1 _13981_/D sky130_fd_sc_hd__mux2_1
X_06819_ _13574_/Q _13579_/Q _13578_/Q vssd1 vssd1 vccd1 vccd1 _06819_/X sky130_fd_sc_hd__and3_1
X_07799_ _07816_/A _07799_/B vssd1 vssd1 vccd1 vccd1 _07799_/Y sky130_fd_sc_hd__nand2_1
X_09538_ _08520_/B _09535_/X _09537_/X _09533_/X vssd1 vssd1 vccd1 vccd1 _09539_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_24_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09469_ _13870_/Q _14223_/Q _09469_/S vssd1 vssd1 vccd1 vccd1 _09469_/X sky130_fd_sc_hd__mux2_1
XFILLER_12_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11500_ _11500_/A _11500_/B vssd1 vssd1 vccd1 vccd1 _11501_/B sky130_fd_sc_hd__or2_1
XFILLER_40_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12480_ _12503_/A1 _12479_/X _12478_/X _12503_/C1 vssd1 vssd1 vccd1 vccd1 _12481_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_156_106 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_628 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11431_ _11431_/A _11431_/B vssd1 vssd1 vccd1 vccd1 _11441_/A sky130_fd_sc_hd__and2_1
XFILLER_22_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14150_ _15127_/CLK _14150_/D vssd1 vssd1 vccd1 vccd1 _14150_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_165_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11362_ _13251_/A _11362_/B _11362_/C vssd1 vssd1 vccd1 vccd1 _11363_/C sky130_fd_sc_hd__or3_1
XFILLER_137_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13101_ _15518_/Q _13119_/S _13105_/B1 _13100_/X vssd1 vssd1 vccd1 vccd1 _15518_/D
+ sky130_fd_sc_hd__a22o_1
X_10313_ _14698_/Q _14883_/Q _10715_/S vssd1 vssd1 vccd1 vccd1 _14698_/D sky130_fd_sc_hd__mux2_1
XFILLER_138_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14081_ _15133_/CLK _14081_/D vssd1 vssd1 vccd1 vccd1 _14081_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_125_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11293_ _15033_/Q _08232_/A _11292_/X vssd1 vssd1 vccd1 vccd1 _15033_/D sky130_fd_sc_hd__a21o_1
XFILLER_4_856 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13032_ _10724_/X _14891_/Q _13038_/S vssd1 vssd1 vccd1 vccd1 _13032_/X sky130_fd_sc_hd__mux2_4
X_10244_ _14629_/Q _14782_/Q _10244_/S vssd1 vssd1 vccd1 vccd1 _14629_/D sky130_fd_sc_hd__mux2_1
XFILLER_180_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10175_ _11861_/A1 _14559_/Q _10192_/S vssd1 vssd1 vccd1 vccd1 _14559_/D sky130_fd_sc_hd__mux2_1
XFILLER_65_1099 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14983_ _15582_/CLK _14983_/D vssd1 vssd1 vccd1 vccd1 _14983_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout180 _11643_/X vssd1 vssd1 vccd1 vccd1 _11675_/S sky130_fd_sc_hd__buf_12
Xfanout191 _09964_/Y vssd1 vssd1 vccd1 vccd1 _09991_/S sky130_fd_sc_hd__buf_12
XFILLER_75_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13934_ _15670_/CLK _13934_/D vssd1 vssd1 vccd1 vccd1 _13934_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_75_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13865_ _15081_/CLK _13865_/D vssd1 vssd1 vccd1 vccd1 _13865_/Q sky130_fd_sc_hd__dfxtp_1
X_15604_ _15638_/CLK _15604_/D vssd1 vssd1 vccd1 vccd1 _15604_/Q sky130_fd_sc_hd__dfxtp_1
X_12816_ _06861_/Y _12813_/X _12814_/X _12815_/X vssd1 vssd1 vccd1 vccd1 _12816_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_188_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13796_ _15422_/CLK _13796_/D vssd1 vssd1 vccd1 vccd1 _13796_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15535_ _15616_/CLK _15535_/D vssd1 vssd1 vccd1 vccd1 _15535_/Q sky130_fd_sc_hd__dfxtp_1
X_12747_ _12754_/B _12747_/B vssd1 vssd1 vccd1 vccd1 _12747_/Y sky130_fd_sc_hd__nor2_1
XFILLER_31_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_798 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12678_ _15345_/Q _12765_/B _12677_/X _12809_/C1 vssd1 vssd1 vccd1 vccd1 _15345_/D
+ sky130_fd_sc_hd__o211a_1
X_15466_ _15507_/CLK _15466_/D vssd1 vssd1 vccd1 vccd1 _15466_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14417_ _15161_/CLK _14417_/D vssd1 vssd1 vccd1 vccd1 _14417_/Q sky130_fd_sc_hd__dfxtp_1
X_11629_ _11629_/A _11629_/B vssd1 vssd1 vccd1 vccd1 _11629_/Y sky130_fd_sc_hd__xnor2_1
X_15397_ _15397_/CLK _15397_/D vssd1 vssd1 vccd1 vccd1 _15397_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_144_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14348_ _15518_/CLK _14348_/D vssd1 vssd1 vccd1 vccd1 _14348_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14279_ _15292_/CLK _14279_/D vssd1 vssd1 vccd1 vccd1 _14279_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_170_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08840_ _13863_/Q _11872_/A1 _08851_/S vssd1 vssd1 vccd1 vccd1 _13863_/D sky130_fd_sc_hd__mux2_1
XTAP_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08771_ _08530_/B _08769_/X _08777_/B _14611_/Q _06685_/Y vssd1 vssd1 vccd1 vccd1
+ _08771_/X sky130_fd_sc_hd__o2111a_1
XFILLER_100_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07722_ _14750_/Q _07750_/A _07721_/Y _07987_/C1 vssd1 vssd1 vccd1 vccd1 _13493_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_84_159 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07653_ _13475_/Q _07650_/B _13476_/Q vssd1 vssd1 vccd1 vccd1 _07653_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_53_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_343 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07584_ _13457_/Q _13456_/Q _07588_/D vssd1 vssd1 vccd1 vccd1 _07587_/B sky130_fd_sc_hd__and3_1
XFILLER_168_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09323_ _09307_/X _09310_/X _09317_/X _09322_/X vssd1 vssd1 vccd1 vccd1 _09323_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_22_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_178_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09254_ _15666_/Q _13400_/Q _09512_/S vssd1 vssd1 vccd1 vccd1 _09254_/X sky130_fd_sc_hd__mux2_1
X_08205_ _13696_/Q _13082_/B2 _08216_/S vssd1 vssd1 vccd1 vccd1 _13696_/D sky130_fd_sc_hd__mux2_1
XFILLER_18_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09185_ _14242_/Q _14274_/Q _14306_/Q _14338_/Q _09438_/S0 _09448_/S1 vssd1 vssd1
+ vccd1 vccd1 _09185_/X sky130_fd_sc_hd__mux4_2
XFILLER_119_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08136_ _13660_/Q _10730_/S _08119_/X _08135_/X vssd1 vssd1 vccd1 vccd1 _13660_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_175_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08067_ _14760_/Q _13638_/Q _08072_/S vssd1 vssd1 vccd1 vccd1 _13638_/D sky130_fd_sc_hd__mux2_1
XFILLER_107_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07018_ _14618_/Q _14650_/Q _07096_/S vssd1 vssd1 vccd1 vccd1 _07018_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08969_ _09130_/A _08962_/X _08965_/X _09450_/B1 vssd1 vssd1 vccd1 vccd1 _08969_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_57_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11980_ _15112_/Q _15080_/Q _15653_/Q _13387_/Q _11993_/S _11992_/A vssd1 vssd1 vccd1
+ vccd1 _11980_/X sky130_fd_sc_hd__mux4_1
XFILLER_72_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10931_ _13214_/A _13215_/B vssd1 vssd1 vccd1 vccd1 _10931_/Y sky130_fd_sc_hd__nand2_1
XFILLER_29_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_215 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10862_ _14894_/Q _15530_/Q _10871_/S vssd1 vssd1 vccd1 vccd1 _14894_/D sky130_fd_sc_hd__mux2_1
X_13650_ _15620_/CLK _13650_/D vssd1 vssd1 vccd1 vccd1 _13650_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12601_ _15139_/Q _15107_/Q _15680_/Q _13414_/Q _12612_/S _12613_/A vssd1 vssd1 vccd1
+ vccd1 _12601_/X sky130_fd_sc_hd__mux4_1
X_13581_ _15534_/CLK _13581_/D vssd1 vssd1 vccd1 vccd1 _13581_/Q sky130_fd_sc_hd__dfxtp_2
XPHY_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10793_ _14825_/Q _15457_/Q _12929_/S vssd1 vssd1 vccd1 vccd1 _14825_/D sky130_fd_sc_hd__mux2_1
XFILLER_12_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12532_ _15136_/Q _15104_/Q _15677_/Q _13411_/Q _12612_/S _12383_/A vssd1 vssd1 vccd1
+ vccd1 _12532_/X sky130_fd_sc_hd__mux4_1
X_15320_ _15332_/CLK _15320_/D vssd1 vssd1 vccd1 vccd1 _15320_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12463_ _15133_/Q _15101_/Q _15674_/Q _13408_/Q _12472_/S _12465_/S1 vssd1 vssd1
+ vccd1 vccd1 _12463_/X sky130_fd_sc_hd__mux4_1
X_15251_ _15298_/CLK _15251_/D vssd1 vssd1 vccd1 vccd1 _15251_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_184_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14202_ _14462_/CLK _14202_/D vssd1 vssd1 vccd1 vccd1 _14202_/Q sky130_fd_sc_hd__dfxtp_1
X_11414_ _11414_/A _13177_/A _11414_/C _11414_/D vssd1 vssd1 vccd1 vccd1 _11437_/B
+ sky130_fd_sc_hd__and4_4
XFILLER_126_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15182_ _15298_/CLK _15182_/D vssd1 vssd1 vccd1 vccd1 _15182_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_184_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12394_ _15130_/Q _15098_/Q _15671_/Q _13405_/Q _12591_/S _12590_/A vssd1 vssd1 vccd1
+ vccd1 _12394_/X sky130_fd_sc_hd__mux4_1
XFILLER_137_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14133_ _15211_/CLK _14133_/D vssd1 vssd1 vccd1 vccd1 _14133_/Q sky130_fd_sc_hd__dfxtp_1
X_11345_ _08233_/B _08379_/X _11344_/X wire438/X vssd1 vssd1 vccd1 vccd1 _11345_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_125_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14064_ _15226_/CLK _14064_/D vssd1 vssd1 vccd1 vccd1 _14064_/Q sky130_fd_sc_hd__dfxtp_1
X_11276_ _11329_/A _08358_/X _11275_/Y _08233_/B vssd1 vssd1 vccd1 vccd1 _11276_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_79_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13015_ _13098_/B2 _13039_/A2 _13014_/X _12944_/A vssd1 vssd1 vccd1 vccd1 _13015_/X
+ sky130_fd_sc_hd__a22o_1
X_10227_ input22/X _14612_/Q _13284_/S vssd1 vssd1 vccd1 vccd1 _14612_/D sky130_fd_sc_hd__mux2_1
XFILLER_79_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_318 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10158_ _14543_/Q _11877_/A1 _10159_/S vssd1 vssd1 vccd1 vccd1 _14543_/D sky130_fd_sc_hd__mux2_1
XFILLER_121_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold3 hold3/A vssd1 vssd1 vccd1 vccd1 hold3/X sky130_fd_sc_hd__bufbuf_16
XFILLER_181_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10089_ _14445_/Q _13098_/B2 _10097_/S vssd1 vssd1 vccd1 vccd1 _14445_/D sky130_fd_sc_hd__mux2_1
X_14966_ _14966_/CLK _14966_/D vssd1 vssd1 vccd1 vccd1 _14966_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13917_ _15507_/CLK _13917_/D vssd1 vssd1 vccd1 vccd1 _13917_/Q sky130_fd_sc_hd__dfxtp_1
X_14897_ _15616_/CLK _14897_/D vssd1 vssd1 vccd1 vccd1 _14897_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_546 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13848_ _15211_/CLK _13848_/D vssd1 vssd1 vccd1 vccd1 _13848_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_74_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13779_ _15397_/CLK _13779_/D vssd1 vssd1 vccd1 vccd1 _13779_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_95_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15518_ _15518_/CLK _15518_/D vssd1 vssd1 vccd1 vccd1 _15518_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_595 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15449_ _15635_/CLK _15449_/D vssd1 vssd1 vccd1 vccd1 _15449_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_4_4_0_clk clkbuf_4_5_0_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_5_9_0_clk/A sky130_fd_sc_hd__clkbuf_8
XFILLER_163_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_175_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09941_ _11861_/A1 _14301_/Q _09958_/S vssd1 vssd1 vccd1 vccd1 _14301_/D sky130_fd_sc_hd__mux2_1
XFILLER_48_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09872_ _11858_/A1 _14234_/Q _09892_/S vssd1 vssd1 vccd1 vccd1 _14234_/D sky130_fd_sc_hd__mux2_1
XFILLER_174_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08823_ _13846_/Q _13322_/A0 _08846_/S vssd1 vssd1 vccd1 vccd1 _13846_/D sky130_fd_sc_hd__mux2_1
XTAP_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08754_ _08754_/A _09829_/B vssd1 vssd1 vccd1 vccd1 _08754_/Y sky130_fd_sc_hd__nand2_1
XFILLER_38_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07705_ _13489_/Q _07732_/A vssd1 vssd1 vccd1 vccd1 _07706_/B sky130_fd_sc_hd__xnor2_1
XFILLER_38_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08685_ _13550_/Q _08685_/A2 _08691_/B1 _13486_/Q vssd1 vssd1 vccd1 vccd1 _08685_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_2619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_92_clk clkbuf_5_24_0_clk/X vssd1 vssd1 vccd1 vccd1 _15616_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_1907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07636_ _07651_/A _07636_/B vssd1 vssd1 vccd1 vccd1 _07636_/Y sky130_fd_sc_hd__nand2_1
XFILLER_54_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07567_ _07571_/B _07567_/B vssd1 vssd1 vccd1 vccd1 _07568_/B sky130_fd_sc_hd__xnor2_1
X_09306_ _09543_/A _09306_/B vssd1 vssd1 vccd1 vccd1 _09306_/X sky130_fd_sc_hd__or2_1
XFILLER_55_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07498_ _14676_/Q _07498_/B _07498_/C vssd1 vssd1 vccd1 vccd1 _07498_/X sky130_fd_sc_hd__and3_1
XFILLER_10_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09237_ _06676_/A _09226_/X _09235_/X _09236_/X vssd1 vssd1 vccd1 vccd1 _09237_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_186_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_407 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09168_ _09446_/A1 _09166_/X _09167_/X vssd1 vssd1 vccd1 vccd1 _09172_/B sky130_fd_sc_hd__a21o_1
XFILLER_163_930 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08119_ _06661_/Y _06771_/C _14901_/Q _08117_/X _10344_/S vssd1 vssd1 vccd1 vccd1
+ _08119_/X sky130_fd_sc_hd__a41o_4
XFILLER_119_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09099_ _09435_/A _09099_/B vssd1 vssd1 vccd1 vccd1 _09099_/X sky130_fd_sc_hd__or2_1
XFILLER_79_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11130_ _11129_/A _10965_/X _11129_/Y vssd1 vssd1 vccd1 vccd1 _11187_/B sky130_fd_sc_hd__a21oi_1
XFILLER_122_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_827 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11061_ _11061_/A vssd1 vssd1 vccd1 vccd1 _11061_/Y sky130_fd_sc_hd__inv_2
XFILLER_135_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10012_ _13080_/B2 _14370_/Q _10028_/S vssd1 vssd1 vccd1 vccd1 _14370_/D sky130_fd_sc_hd__mux2_1
XFILLER_89_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14820_ _15452_/CLK _14820_/D vssd1 vssd1 vccd1 vccd1 _14820_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14751_ _15643_/CLK _14751_/D vssd1 vssd1 vccd1 vccd1 _14751_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_3854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_74 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11963_ _12273_/A1 _11958_/X _11961_/X _11962_/X _08449_/A vssd1 vssd1 vccd1 vccd1
+ _11975_/B sky130_fd_sc_hd__a221o_1
XFILLER_91_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_83_clk clkbuf_5_14_0_clk/X vssd1 vssd1 vccd1 vccd1 _15591_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_3887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13702_ _15304_/CLK _13702_/D vssd1 vssd1 vccd1 vccd1 _13702_/Q sky130_fd_sc_hd__dfxtp_1
X_10914_ _11476_/B _10944_/B vssd1 vssd1 vccd1 vccd1 _10914_/Y sky130_fd_sc_hd__nand2_1
XTAP_3898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11894_ _12273_/A1 _11889_/X _11892_/X _11893_/X _08449_/A vssd1 vssd1 vccd1 vccd1
+ _11906_/B sky130_fd_sc_hd__a221o_1
X_14682_ _15620_/CLK _14682_/D vssd1 vssd1 vccd1 vccd1 _14682_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10845_ _14877_/Q _13791_/Q _12927_/S vssd1 vssd1 vccd1 vccd1 _14877_/D sky130_fd_sc_hd__mux2_1
X_13633_ _14506_/CLK _13633_/D vssd1 vssd1 vccd1 vccd1 _13633_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10776_ _14808_/Q _15440_/Q _12918_/S vssd1 vssd1 vccd1 vccd1 _14808_/D sky130_fd_sc_hd__mux2_1
X_13564_ _13565_/CLK _13564_/D vssd1 vssd1 vccd1 vccd1 _13564_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15303_ _15303_/CLK _15303_/D vssd1 vssd1 vccd1 vccd1 _15303_/Q sky130_fd_sc_hd__dfxtp_1
X_12515_ _12618_/A1 _12510_/X _12513_/X _12514_/X _12515_/C1 vssd1 vssd1 vccd1 vccd1
+ _12527_/B sky130_fd_sc_hd__a221o_1
X_13495_ _13632_/CLK _13495_/D vssd1 vssd1 vccd1 vccd1 _13495_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_12_284 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12446_ _12503_/A1 _12441_/X _12444_/X _12445_/X _08449_/A vssd1 vssd1 vccd1 vccd1
+ _12458_/B sky130_fd_sc_hd__a221o_1
X_15234_ _15298_/CLK _15234_/D vssd1 vssd1 vccd1 vccd1 _15234_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_138_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15165_ _15298_/CLK _15165_/D vssd1 vssd1 vccd1 vccd1 _15165_/Q sky130_fd_sc_hd__dfxtp_1
X_12377_ _12618_/A1 _12372_/X _12375_/X _12376_/X _12515_/C1 vssd1 vssd1 vccd1 vccd1
+ _12389_/B sky130_fd_sc_hd__a221o_1
XFILLER_154_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11328_ _15038_/Q _11302_/A _08349_/X _11303_/A _11327_/X vssd1 vssd1 vccd1 vccd1
+ _15038_/D sky130_fd_sc_hd__o221a_1
XFILLER_5_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14116_ _14225_/CLK _14116_/D vssd1 vssd1 vccd1 vccd1 _14116_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15096_ _15096_/CLK _15096_/D vssd1 vssd1 vccd1 vccd1 _15096_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11259_ _11242_/Y _11258_/Y _11259_/S vssd1 vssd1 vccd1 vccd1 _11259_/X sky130_fd_sc_hd__mux2_1
X_14047_ _15656_/CLK _14047_/D vssd1 vssd1 vccd1 vccd1 _14047_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_991 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14949_ _15014_/CLK _14949_/D vssd1 vssd1 vccd1 vccd1 _14949_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_74_clk clkbuf_5_15_0_clk/X vssd1 vssd1 vccd1 vccd1 _15628_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_91_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08470_ _08465_/B _08487_/B _12906_/S vssd1 vssd1 vccd1 vccd1 _08470_/X sky130_fd_sc_hd__o21a_4
XFILLER_51_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07421_ _13330_/A0 _13394_/Q _07481_/S vssd1 vssd1 vccd1 vccd1 _13394_/D sky130_fd_sc_hd__mux2_1
XFILLER_51_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07352_ _07352_/A _07352_/B vssd1 vssd1 vccd1 vccd1 _07352_/Y sky130_fd_sc_hd__nor2_1
XFILLER_148_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07283_ _13920_/Q _15507_/Q _07339_/S vssd1 vssd1 vccd1 vccd1 _07284_/A sky130_fd_sc_hd__mux2_8
X_09022_ _14428_/Q _13130_/B1 _08520_/B _09021_/X vssd1 vssd1 vccd1 vccd1 _09022_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_136_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09924_ _13344_/A0 _14285_/Q _09925_/S vssd1 vssd1 vccd1 vccd1 _14285_/D sky130_fd_sc_hd__mux2_1
XFILLER_59_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09855_ _14219_/Q _13098_/B2 _09863_/S vssd1 vssd1 vccd1 vccd1 _14219_/D sky130_fd_sc_hd__mux2_1
XTAP_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08806_ _11873_/A1 _13832_/Q _08816_/S vssd1 vssd1 vccd1 vccd1 _13832_/D sky130_fd_sc_hd__mux2_1
XFILLER_85_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09786_ _14153_/Q _13341_/A0 _09795_/S vssd1 vssd1 vccd1 vccd1 _14153_/D sky130_fd_sc_hd__mux2_1
X_06998_ _14727_/Q _14728_/Q _14726_/Q _14725_/Q vssd1 vssd1 vccd1 vccd1 _07504_/B
+ sky130_fd_sc_hd__or4bb_4
XTAP_3117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08737_ _13646_/Q _08523_/Y _08747_/B1 _13479_/Q vssd1 vssd1 vccd1 vccd1 _08737_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_73_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_65_clk clkbuf_5_11_0_clk/X vssd1 vssd1 vccd1 vccd1 _15577_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_2427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_106 _14741_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_332 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_117 _07192_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_128 _08453_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08668_ _08532_/B _08668_/B _08668_/C _08668_/D vssd1 vssd1 vccd1 vccd1 _08668_/X
+ sky130_fd_sc_hd__and4b_4
XTAP_2449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07619_ _14755_/Q _07629_/A _07618_/X _07949_/C1 vssd1 vssd1 vccd1 vccd1 _13466_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_1748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08599_ _13784_/Q _08626_/S _08598_/X vssd1 vssd1 vccd1 vccd1 _13784_/D sky130_fd_sc_hd__o21a_1
XTAP_1759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10630_ _14744_/Q _10629_/X _10630_/S vssd1 vssd1 vccd1 vccd1 _14744_/D sky130_fd_sc_hd__mux2_1
XFILLER_14_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10561_ _14924_/Q _10561_/B _10561_/C vssd1 vssd1 vccd1 vccd1 _11777_/B sky130_fd_sc_hd__nor3_4
XFILLER_10_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12300_ _14472_/Q _14440_/Q _13861_/Q _14214_/Q _12612_/S _12383_/A vssd1 vssd1 vccd1
+ vccd1 _12300_/X sky130_fd_sc_hd__mux4_1
XFILLER_155_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13280_ _15364_/Q _15611_/Q _13309_/A vssd1 vssd1 vccd1 vccd1 _15611_/D sky130_fd_sc_hd__mux2_1
X_10492_ _10520_/A1 _13790_/Q _13758_/Q _10520_/B2 vssd1 vssd1 vccd1 vccd1 _10492_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_10_788 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12231_ _14469_/Q _14437_/Q _13858_/Q _14211_/Q _12499_/S _12486_/S1 vssd1 vssd1
+ vccd1 vccd1 _12231_/X sky130_fd_sc_hd__mux4_1
XFILLER_163_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12162_ _14466_/Q _14434_/Q _13855_/Q _14208_/Q _12246_/S _12452_/A vssd1 vssd1 vccd1
+ vccd1 _12162_/X sky130_fd_sc_hd__mux4_1
XFILLER_108_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_943 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11113_ _11115_/S _11056_/X _11094_/Y vssd1 vssd1 vccd1 vccd1 _11113_/X sky130_fd_sc_hd__a21o_1
XFILLER_123_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12093_ _14463_/Q _14431_/Q _13852_/Q _14205_/Q _12472_/S _12465_/S1 vssd1 vssd1
+ vccd1 vccd1 _12093_/X sky130_fd_sc_hd__mux4_1
X_11044_ _11044_/A _11044_/B vssd1 vssd1 vccd1 vccd1 _11044_/Y sky130_fd_sc_hd__nor2_1
XFILLER_89_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14803_ _15646_/CLK _14803_/D vssd1 vssd1 vccd1 vccd1 _14803_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_76_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_56_clk clkbuf_5_11_0_clk/X vssd1 vssd1 vccd1 vccd1 _15017_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_29_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12995_ _15478_/Q _13119_/S _13025_/B1 _12994_/X vssd1 vssd1 vccd1 vccd1 _15478_/D
+ sky130_fd_sc_hd__a22o_1
XTAP_3662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14734_ _15462_/CLK _14734_/D vssd1 vssd1 vccd1 vccd1 _14734_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_3684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11946_ _12406_/A _11946_/B vssd1 vssd1 vccd1 vccd1 _11946_/X sky130_fd_sc_hd__and2_1
XTAP_3695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14665_ _15636_/CLK _14665_/D vssd1 vssd1 vccd1 vccd1 _14665_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11877_ _15298_/Q _11877_/A1 _11878_/S vssd1 vssd1 vccd1 vccd1 _15298_/D sky130_fd_sc_hd__mux2_1
XTAP_2994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13616_ _15372_/CLK _13616_/D vssd1 vssd1 vccd1 vccd1 _13616_/Q sky130_fd_sc_hd__dfxtp_1
X_10828_ _14860_/Q _07225_/A _10868_/S vssd1 vssd1 vccd1 vccd1 _14860_/D sky130_fd_sc_hd__mux2_1
X_14596_ _15536_/CLK _14596_/D vssd1 vssd1 vccd1 vccd1 _14596_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_38_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13547_ _15374_/CLK _13547_/D vssd1 vssd1 vccd1 vccd1 _13547_/Q sky130_fd_sc_hd__dfxtp_1
X_10759_ _15423_/Q _14791_/Q _10759_/S vssd1 vssd1 vccd1 vccd1 _14791_/D sky130_fd_sc_hd__mux2_1
XFILLER_173_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13478_ _15542_/CLK _13478_/D vssd1 vssd1 vccd1 vccd1 _13478_/Q sky130_fd_sc_hd__dfxtp_4
X_15217_ _15281_/CLK _15217_/D vssd1 vssd1 vccd1 vccd1 _15217_/Q sky130_fd_sc_hd__dfxtp_1
X_12429_ _12563_/A _12429_/B vssd1 vssd1 vccd1 vccd1 _12429_/X sky130_fd_sc_hd__and2_1
XFILLER_127_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_911 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15148_ _15281_/CLK _15148_/D vssd1 vssd1 vccd1 vccd1 _15148_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_181_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07970_ _13558_/Q _07970_/B vssd1 vssd1 vccd1 vccd1 _07971_/B sky130_fd_sc_hd__xor2_1
X_15079_ _15652_/CLK _15079_/D vssd1 vssd1 vccd1 vccd1 _15079_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_45_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06921_ _06921_/A _06921_/B _06916_/X _06911_/X vssd1 vssd1 vccd1 vccd1 _06922_/C
+ sky130_fd_sc_hd__or4bb_1
XFILLER_84_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09640_ _14013_/Q _13072_/B2 _09660_/S vssd1 vssd1 vccd1 vccd1 _14013_/D sky130_fd_sc_hd__mux2_1
X_06852_ _12904_/S _06997_/A vssd1 vssd1 vccd1 vccd1 _06852_/Y sky130_fd_sc_hd__nand2_2
XFILLER_110_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09571_ _13947_/Q _13327_/A0 _09589_/S vssd1 vssd1 vccd1 vccd1 _13947_/D sky130_fd_sc_hd__mux2_1
X_06783_ _14584_/Q _14583_/Q _14585_/Q vssd1 vssd1 vccd1 vccd1 _06987_/D sky130_fd_sc_hd__and3_1
XFILLER_48_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_47_clk clkbuf_5_8_0_clk/X vssd1 vssd1 vccd1 vccd1 _15558_/CLK sky130_fd_sc_hd__clkbuf_16
X_08522_ _14608_/Q _14610_/Q _08536_/C _13127_/C vssd1 vssd1 vccd1 vccd1 _08532_/B
+ sky130_fd_sc_hd__or4_4
XFILLER_70_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08453_ _08453_/A _08773_/B vssd1 vssd1 vccd1 vccd1 _08453_/X sky130_fd_sc_hd__and2_1
XFILLER_63_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07404_ _14741_/Q _07403_/X _07500_/S vssd1 vssd1 vccd1 vccd1 _07404_/X sky130_fd_sc_hd__mux2_4
X_08384_ _07278_/B _10523_/A2 _08383_/X vssd1 vssd1 vccd1 vccd1 _13202_/B sky130_fd_sc_hd__a21o_4
XFILLER_51_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07335_ _15308_/Q _15464_/Q _07335_/S vssd1 vssd1 vccd1 vccd1 _07336_/A sky130_fd_sc_hd__mux2_8
XFILLER_91_1084 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07266_ _07263_/X _07264_/X _07273_/B _07274_/A vssd1 vssd1 vccd1 vccd1 _07268_/A
+ sky130_fd_sc_hd__a31o_1
X_09005_ _14008_/Q _13976_/Q _09005_/S vssd1 vssd1 vccd1 vccd1 _09005_/X sky130_fd_sc_hd__mux2_1
XFILLER_117_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07197_ _07197_/A _07197_/B vssd1 vssd1 vccd1 vccd1 _07197_/X sky130_fd_sc_hd__xor2_1
XFILLER_3_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout510 _14710_/Q vssd1 vssd1 vccd1 vccd1 _07498_/C sky130_fd_sc_hd__buf_12
Xfanout521 _14605_/Q vssd1 vssd1 vccd1 vccd1 _09435_/A sky130_fd_sc_hd__buf_12
X_09907_ _11860_/A1 _14268_/Q _09925_/S vssd1 vssd1 vccd1 vccd1 _14268_/D sky130_fd_sc_hd__mux2_1
Xfanout532 _09448_/S1 vssd1 vssd1 vccd1 vccd1 _09446_/A1 sky130_fd_sc_hd__buf_12
Xfanout543 _14604_/Q vssd1 vssd1 vccd1 vccd1 _08487_/A sky130_fd_sc_hd__buf_12
Xfanout554 _08490_/A1 vssd1 vssd1 vccd1 vccd1 _09438_/S0 sky130_fd_sc_hd__buf_8
XFILLER_101_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout565 _08490_/A1 vssd1 vssd1 vccd1 vccd1 _08910_/S sky130_fd_sc_hd__buf_12
XFILLER_47_906 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout576 _12468_/A1 vssd1 vssd1 vccd1 vccd1 _12500_/B1 sky130_fd_sc_hd__buf_12
X_09838_ _14202_/Q _11858_/A1 _09858_/S vssd1 vssd1 vccd1 vccd1 _14202_/D sky130_fd_sc_hd__mux2_1
XTAP_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout587 _12061_/A vssd1 vssd1 vccd1 vccd1 _12080_/A sky130_fd_sc_hd__buf_6
Xfanout598 fanout600/X vssd1 vssd1 vccd1 vccd1 _12383_/A sky130_fd_sc_hd__buf_12
XFILLER_86_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09769_ _14136_/Q _11649_/A0 _09795_/S vssd1 vssd1 vccd1 vccd1 _14136_/D sky130_fd_sc_hd__mux2_1
XFILLER_6_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_38_clk clkbuf_5_9_0_clk/X vssd1 vssd1 vccd1 vccd1 _15462_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_27_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11800_ _15223_/Q _13080_/B2 _11816_/S vssd1 vssd1 vccd1 vccd1 _15223_/D sky130_fd_sc_hd__mux2_1
XTAP_2224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12780_ _13436_/Q _12647_/B _08030_/Y _13603_/Q _12737_/A vssd1 vssd1 vccd1 vccd1
+ _12780_/X sky130_fd_sc_hd__a221o_2
XTAP_1501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11731_ _15160_/Q _11872_/A1 _11742_/S vssd1 vssd1 vccd1 vccd1 _15160_/D sky130_fd_sc_hd__mux2_1
XTAP_1534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14450_ _15200_/CLK _14450_/D vssd1 vssd1 vccd1 vccd1 _14450_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11662_ _13337_/A0 _15094_/Q _11675_/S vssd1 vssd1 vccd1 vccd1 _15094_/D sky130_fd_sc_hd__mux2_1
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13401_ _15667_/CLK _13401_/D vssd1 vssd1 vccd1 vccd1 _13401_/Q sky130_fd_sc_hd__dfxtp_1
X_10613_ _13720_/Q _10602_/B _10612_/X vssd1 vssd1 vccd1 vccd1 _10613_/X sky130_fd_sc_hd__a21o_1
X_11593_ _13233_/B _11593_/B vssd1 vssd1 vccd1 vccd1 _11604_/A sky130_fd_sc_hd__nor2_1
X_14381_ _15286_/CLK _14381_/D vssd1 vssd1 vccd1 vccd1 _14381_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10544_ _11563_/A _11561_/A vssd1 vssd1 vccd1 vccd1 _10544_/X sky130_fd_sc_hd__and2b_1
X_13332_ _13332_/A0 _15662_/Q _13345_/S vssd1 vssd1 vccd1 vccd1 _15662_/D sky130_fd_sc_hd__mux2_1
XFILLER_6_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13263_ _15347_/Q _15594_/Q _13300_/S vssd1 vssd1 vccd1 vccd1 _15594_/D sky130_fd_sc_hd__mux2_1
X_10475_ _07235_/B _10481_/B _10474_/X vssd1 vssd1 vccd1 vccd1 _13226_/B sky130_fd_sc_hd__a21o_4
XFILLER_182_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15002_ _15006_/CLK _15002_/D vssd1 vssd1 vccd1 vccd1 _15002_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_157_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_996 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12214_ _12502_/S _12214_/B vssd1 vssd1 vccd1 vccd1 _12214_/X sky130_fd_sc_hd__or2_1
X_13194_ _15565_/Q _13214_/B _13193_/X vssd1 vssd1 vccd1 vccd1 _15565_/D sky130_fd_sc_hd__a21o_1
XFILLER_124_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12145_ _12168_/A _12145_/B vssd1 vssd1 vccd1 vccd1 _12145_/X sky130_fd_sc_hd__or2_1
XFILLER_155_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12076_ _12582_/A _12076_/B vssd1 vssd1 vccd1 vccd1 _12076_/X sky130_fd_sc_hd__or2_1
XFILLER_96_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11027_ _11027_/A _11294_/B vssd1 vssd1 vccd1 vccd1 _11027_/X sky130_fd_sc_hd__and2_1
XFILLER_49_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_29_clk clkbuf_opt_2_0_clk/X vssd1 vssd1 vccd1 vccd1 _15520_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_64_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12978_ _10634_/X _14873_/Q _13029_/S vssd1 vssd1 vccd1 vccd1 _12978_/X sky130_fd_sc_hd__mux2_4
XFILLER_45_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14717_ _15543_/CLK _14717_/D vssd1 vssd1 vccd1 vccd1 _14717_/Q sky130_fd_sc_hd__dfxtp_4
X_11929_ _13134_/A _11929_/B _11929_/C vssd1 vssd1 vccd1 vccd1 _11929_/X sky130_fd_sc_hd__and3_2
XFILLER_61_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14648_ _15619_/CLK _14648_/D vssd1 vssd1 vccd1 vccd1 _14648_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_162_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_17 _15071_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_28 _14747_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_39 input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14579_ _15335_/CLK _14579_/D vssd1 vssd1 vccd1 vccd1 _14579_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_174_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07120_ _14840_/Q _14832_/Q _07146_/S vssd1 vssd1 vccd1 vccd1 _07121_/B sky130_fd_sc_hd__mux2_1
XFILLER_119_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_855 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07051_ _14629_/Q _14661_/Q _07078_/S vssd1 vssd1 vccd1 vccd1 _07051_/X sky130_fd_sc_hd__mux2_1
XFILLER_118_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput102 _07107_/X vssd1 vssd1 vccd1 vccd1 ext_write_strobe[3] sky130_fd_sc_hd__clkbuf_2
XFILLER_161_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_270 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07953_ _13554_/Q _13553_/Q vssd1 vssd1 vccd1 vccd1 _07961_/D sky130_fd_sc_hd__and2_1
XFILLER_141_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06904_ _15378_/Q _06733_/Y _15377_/Q _07571_/A _06903_/X vssd1 vssd1 vccd1 vccd1
+ _06904_/X sky130_fd_sc_hd__a221o_1
X_07884_ _13536_/Q _13535_/Q _07884_/C _07884_/D vssd1 vssd1 vccd1 vccd1 _07900_/C
+ sky130_fd_sc_hd__and4_4
XFILLER_56_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09623_ _13997_/Q _13104_/B2 _09627_/S vssd1 vssd1 vccd1 vccd1 _13997_/D sky130_fd_sc_hd__mux2_1
X_06835_ _08668_/B _14906_/Q _14909_/Q _08501_/A _06834_/Y vssd1 vssd1 vccd1 vccd1
+ _06835_/X sky130_fd_sc_hd__o221a_1
XFILLER_95_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09554_ _09554_/A _09554_/B _09554_/C vssd1 vssd1 vccd1 vccd1 _09554_/X sky130_fd_sc_hd__and3_1
XFILLER_102_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06766_ _14929_/Q vssd1 vssd1 vccd1 vccd1 _10581_/A sky130_fd_sc_hd__inv_2
XFILLER_83_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08505_ _14613_/Q _14614_/Q _13131_/C vssd1 vssd1 vccd1 vccd1 _13127_/C sky130_fd_sc_hd__or3_4
X_06697_ _14513_/Q vssd1 vssd1 vccd1 vccd1 _06697_/Y sky130_fd_sc_hd__inv_2
X_09485_ _14095_/Q _09522_/A2 _09519_/B1 _14063_/Q _09543_/A vssd1 vssd1 vccd1 vccd1
+ _09485_/X sky130_fd_sc_hd__a221o_1
XFILLER_52_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08436_ _13748_/Q _12906_/S _08426_/B _08435_/X vssd1 vssd1 vccd1 vccd1 _13748_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_24_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08367_ _08346_/X _08366_/Y _11318_/S vssd1 vssd1 vccd1 vccd1 _08367_/X sky130_fd_sc_hd__mux2_1
XFILLER_11_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07318_ _07312_/X _07314_/Y _07352_/A _07352_/B vssd1 vssd1 vccd1 vccd1 _07360_/A
+ sky130_fd_sc_hd__a22o_1
X_08298_ _11297_/S _08298_/B vssd1 vssd1 vccd1 vccd1 _08299_/C sky130_fd_sc_hd__nand2_1
X_07249_ _13926_/Q _15513_/Q _07334_/S vssd1 vssd1 vccd1 vccd1 _07264_/A sky130_fd_sc_hd__mux2_8
XFILLER_164_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10260_ _14645_/Q _14798_/Q _10730_/S vssd1 vssd1 vccd1 vccd1 _14645_/D sky130_fd_sc_hd__mux2_1
XFILLER_11_76 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10191_ _11877_/A1 _14575_/Q _10192_/S vssd1 vssd1 vccd1 vccd1 _14575_/D sky130_fd_sc_hd__mux2_1
XFILLER_105_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout340 _11681_/A0 vssd1 vssd1 vccd1 vccd1 _13323_/A0 sky130_fd_sc_hd__buf_6
XFILLER_143_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout351 _06857_/X vssd1 vssd1 vccd1 vccd1 _12834_/B sky130_fd_sc_hd__buf_12
Xfanout362 _08519_/X vssd1 vssd1 vccd1 vccd1 _13130_/C1 sky130_fd_sc_hd__buf_12
X_13950_ _15212_/CLK _13950_/D vssd1 vssd1 vccd1 vccd1 _13950_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout373 _11349_/B vssd1 vssd1 vccd1 vccd1 _11013_/A sky130_fd_sc_hd__buf_6
XFILLER_74_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout384 _08236_/X vssd1 vssd1 vccd1 vccd1 _11362_/B sky130_fd_sc_hd__buf_12
XFILLER_4_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout395 _08228_/X vssd1 vssd1 vccd1 vccd1 _11371_/A sky130_fd_sc_hd__buf_12
XFILLER_46_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12901_ _15429_/Q _15614_/Q _12932_/S vssd1 vssd1 vccd1 vccd1 _15429_/D sky130_fd_sc_hd__mux2_1
XFILLER_74_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13881_ _15655_/CLK _13881_/D vssd1 vssd1 vccd1 vccd1 _13881_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_74_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15620_ _15620_/CLK _15620_/D vssd1 vssd1 vccd1 vccd1 _15620_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_46_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12832_ _15366_/Q _12759_/B _12831_/X _12832_/C1 vssd1 vssd1 vccd1 vccd1 _15366_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_185_1038 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_994 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15551_ _15676_/CLK _15551_/D vssd1 vssd1 vccd1 vccd1 _15551_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12763_ _13601_/Q _12762_/X _12763_/S vssd1 vssd1 vccd1 vccd1 _12763_/X sky130_fd_sc_hd__mux2_1
XFILLER_43_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14502_ _15386_/CLK _14502_/D vssd1 vssd1 vccd1 vccd1 _14502_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11714_ _15143_/Q _13322_/A0 _11741_/S vssd1 vssd1 vccd1 vccd1 _15143_/D sky130_fd_sc_hd__mux2_1
XTAP_1364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15482_ _15523_/CLK _15482_/D vssd1 vssd1 vccd1 vccd1 _15482_/Q sky130_fd_sc_hd__dfxtp_1
X_12694_ _15347_/Q _12765_/B _12693_/X _12809_/C1 vssd1 vssd1 vccd1 vccd1 _15347_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_14_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_148 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14433_ _15663_/CLK _14433_/D vssd1 vssd1 vccd1 vccd1 _14433_/Q sky130_fd_sc_hd__dfxtp_1
X_11645_ _11853_/A1 _15077_/Q _11675_/S vssd1 vssd1 vccd1 vccd1 _15077_/D sky130_fd_sc_hd__mux2_1
XFILLER_168_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_1071 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput15 ext_read_data[22] vssd1 vssd1 vccd1 vccd1 input15/X sky130_fd_sc_hd__buf_4
X_14364_ _15279_/CLK _14364_/D vssd1 vssd1 vccd1 vccd1 _14364_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_168_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11576_ _11576_/A _11576_/B _11576_/C _11576_/D vssd1 vssd1 vccd1 vccd1 _11576_/Y
+ sky130_fd_sc_hd__nor4_1
Xinput26 ext_read_data[3] vssd1 vssd1 vccd1 vccd1 input26/X sky130_fd_sc_hd__buf_6
XFILLER_167_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13315_ _15646_/Q _12828_/B _13316_/S vssd1 vssd1 vccd1 vccd1 _15646_/D sky130_fd_sc_hd__mux2_1
X_10527_ _10527_/A _10527_/B _10527_/C _10527_/D vssd1 vssd1 vccd1 vccd1 _10529_/A
+ sky130_fd_sc_hd__or4_1
XFILLER_143_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14295_ _15276_/CLK _14295_/D vssd1 vssd1 vccd1 vccd1 _14295_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_171_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10458_ _08244_/A _13747_/Q _15425_/Q _08244_/B vssd1 vssd1 vccd1 vccd1 _10458_/X
+ sky130_fd_sc_hd__a22o_1
X_13246_ _13217_/A _11626_/A _13214_/B vssd1 vssd1 vccd1 vccd1 _13246_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_182_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10389_ _10387_/X _10389_/B vssd1 vssd1 vccd1 vccd1 _10390_/C sky130_fd_sc_hd__nand2b_1
XFILLER_97_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13177_ _13177_/A _13252_/B vssd1 vssd1 vccd1 vccd1 _13177_/Y sky130_fd_sc_hd__nor2_1
XFILLER_97_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12128_ _12477_/A1 _12127_/X _12490_/A vssd1 vssd1 vccd1 vccd1 _12128_/X sky130_fd_sc_hd__a21o_1
XFILLER_111_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12059_ _12500_/A1 _12058_/X _12582_/A vssd1 vssd1 vccd1 vccd1 _12059_/X sky130_fd_sc_hd__a21o_1
XFILLER_42_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09270_ _13893_/Q _09522_/A2 _08512_/B _14408_/Q _08507_/A vssd1 vssd1 vccd1 vccd1
+ _09270_/X sky130_fd_sc_hd__a221o_1
XFILLER_33_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08221_ _13712_/Q _13350_/A0 _08221_/S vssd1 vssd1 vccd1 vccd1 _13712_/D sky130_fd_sc_hd__mux2_1
XFILLER_159_660 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08152_ _08121_/X _08151_/X _08119_/X vssd1 vssd1 vccd1 vccd1 _08152_/X sky130_fd_sc_hd__a21o_1
X_07103_ _07131_/A _07103_/B vssd1 vssd1 vccd1 vccd1 _07103_/X sky130_fd_sc_hd__and2_4
XFILLER_119_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08083_ _08083_/A _08083_/B vssd1 vssd1 vccd1 vccd1 _08083_/Y sky130_fd_sc_hd__nand2_1
XFILLER_146_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_9_clk clkbuf_5_2_0_clk/X vssd1 vssd1 vccd1 vccd1 _15659_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_134_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07034_ _07033_/X _13590_/Q _12728_/S vssd1 vssd1 vccd1 vccd1 _07034_/X sky130_fd_sc_hd__mux2_1
XFILLER_162_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08985_ _09130_/A _08985_/B _08985_/C vssd1 vssd1 vccd1 vccd1 _08985_/X sky130_fd_sc_hd__and3_1
XFILLER_29_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07936_ _13548_/Q _13547_/Q _07935_/D _13549_/Q vssd1 vssd1 vccd1 vccd1 _07936_/Y
+ sky130_fd_sc_hd__a31oi_1
XFILLER_180_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07867_ _07874_/A _07866_/X input35/X vssd1 vssd1 vccd1 vccd1 _07867_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_29_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09606_ _13980_/Q _13328_/A0 _09627_/S vssd1 vssd1 vccd1 vccd1 _13980_/D sky130_fd_sc_hd__mux2_1
XFILLER_16_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06818_ _06806_/X _06815_/X _06817_/X _15540_/Q vssd1 vssd1 vccd1 vccd1 _06851_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_43_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07798_ _13513_/Q _07798_/B vssd1 vssd1 vccd1 vccd1 _07799_/B sky130_fd_sc_hd__xnor2_1
XFILLER_25_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09537_ _08668_/D _09534_/X _09536_/X vssd1 vssd1 vccd1 vccd1 _09537_/X sky130_fd_sc_hd__a21o_1
XFILLER_25_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06749_ _13448_/Q vssd1 vssd1 vccd1 vccd1 _06749_/Y sky130_fd_sc_hd__inv_2
XFILLER_25_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09468_ _14255_/Q _14287_/Q _14319_/Q _14351_/Q _09342_/S _13144_/A0 vssd1 vssd1
+ vccd1 vccd1 _09468_/X sky130_fd_sc_hd__mux4_1
XFILLER_184_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08419_ _14596_/Q _14595_/Q _08777_/A _13120_/S _14927_/D vssd1 vssd1 vccd1 vccd1
+ _08419_/X sky130_fd_sc_hd__a32o_1
XFILLER_185_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09399_ _13963_/Q _13705_/Q _09535_/S vssd1 vssd1 vccd1 vccd1 _09399_/X sky130_fd_sc_hd__mux2_1
XFILLER_40_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11430_ _11431_/A _11431_/B vssd1 vssd1 vccd1 vccd1 _11430_/X sky130_fd_sc_hd__or2_1
XFILLER_137_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11361_ _11360_/Y _07104_/C _11641_/S vssd1 vssd1 vccd1 vccd1 _15044_/D sky130_fd_sc_hd__mux2_1
XFILLER_180_600 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10312_ _14697_/Q _14882_/Q _10715_/S vssd1 vssd1 vccd1 vccd1 _14697_/D sky130_fd_sc_hd__mux2_1
X_13100_ _13017_/X _13104_/A2 _13104_/B1 _13343_/A0 vssd1 vssd1 vccd1 vccd1 _13100_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_164_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11292_ _08233_/B _08299_/X _11290_/Y _11291_/Y wire438/X vssd1 vssd1 vccd1 vccd1
+ _11292_/X sky130_fd_sc_hd__o221a_1
X_14080_ _15331_/CLK _14080_/D vssd1 vssd1 vccd1 vccd1 _14080_/Q sky130_fd_sc_hd__dfxtp_1
X_10243_ _14628_/Q _14781_/Q _10650_/S vssd1 vssd1 vccd1 vccd1 _14628_/D sky130_fd_sc_hd__mux2_1
XFILLER_180_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13031_ _15490_/Q _13093_/A2 _13116_/C _13030_/X vssd1 vssd1 vccd1 vccd1 _15490_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_98_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10174_ _11860_/A1 _14558_/Q _10192_/S vssd1 vssd1 vccd1 vccd1 _14558_/D sky130_fd_sc_hd__mux2_1
XFILLER_160_390 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_96 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14982_ _15017_/CLK _14982_/D vssd1 vssd1 vccd1 vccd1 _14982_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout170 _11818_/Y vssd1 vssd1 vccd1 vccd1 _11850_/S sky130_fd_sc_hd__buf_12
Xfanout181 _10132_/Y vssd1 vssd1 vccd1 vccd1 _10159_/S sky130_fd_sc_hd__buf_12
XFILLER_19_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout192 _09964_/Y vssd1 vssd1 vccd1 vccd1 _09996_/S sky130_fd_sc_hd__buf_12
XFILLER_59_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13933_ _15315_/CLK _13933_/D vssd1 vssd1 vccd1 vccd1 _13933_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13864_ _14485_/CLK _13864_/D vssd1 vssd1 vccd1 vccd1 _13864_/Q sky130_fd_sc_hd__dfxtp_1
X_15603_ _15637_/CLK _15603_/D vssd1 vssd1 vccd1 vccd1 _15603_/Q sky130_fd_sc_hd__dfxtp_1
X_12815_ _13441_/Q _12647_/B _08030_/Y _13608_/Q _12743_/A vssd1 vssd1 vccd1 vccd1
+ _12815_/X sky130_fd_sc_hd__a221o_1
X_13795_ _14493_/CLK _13795_/D vssd1 vssd1 vccd1 vccd1 _13795_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15534_ _15534_/CLK _15534_/D vssd1 vssd1 vccd1 vccd1 _15534_/Q sky130_fd_sc_hd__dfxtp_1
X_12746_ _15354_/Q _12745_/C _15355_/Q vssd1 vssd1 vccd1 vccd1 _12747_/B sky130_fd_sc_hd__a21oi_1
XFILLER_31_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15465_ _15497_/CLK _15465_/D vssd1 vssd1 vccd1 vccd1 _15465_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_179_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12677_ _12737_/A _12677_/B vssd1 vssd1 vccd1 vccd1 _12677_/X sky130_fd_sc_hd__or2_1
XFILLER_30_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14416_ _15315_/CLK _14416_/D vssd1 vssd1 vccd1 vccd1 _14416_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_175_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11628_ _11621_/A _11621_/B _13242_/B _11617_/Y vssd1 vssd1 vccd1 vccd1 _11629_/B
+ sky130_fd_sc_hd__a2bb2o_2
X_15396_ _15397_/CLK _15396_/D vssd1 vssd1 vccd1 vccd1 _15396_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14347_ _15527_/CLK _14347_/D vssd1 vssd1 vccd1 vccd1 _14347_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_183_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11559_ _11557_/Y _11558_/X _15064_/Q _11614_/S vssd1 vssd1 vccd1 vccd1 _15064_/D
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_10_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14278_ _15301_/CLK _14278_/D vssd1 vssd1 vccd1 vccd1 _14278_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13229_ _13229_/A _13229_/B vssd1 vssd1 vccd1 vccd1 _13229_/Y sky130_fd_sc_hd__nor2_1
XFILLER_98_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08770_ hold5/A _14592_/Q _08770_/C _12946_/B vssd1 vssd1 vccd1 vccd1 _08779_/A sky130_fd_sc_hd__or4b_2
XTAP_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07721_ _07750_/A _07721_/B vssd1 vssd1 vccd1 vccd1 _07721_/Y sky130_fd_sc_hd__nand2_1
XFILLER_38_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07652_ _14764_/Q _07651_/A _07651_/Y _08012_/C1 vssd1 vssd1 vccd1 vccd1 _13475_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_19_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07583_ _13457_/Q _07583_/B vssd1 vssd1 vccd1 vccd1 _07583_/Y sky130_fd_sc_hd__nor2_1
XFILLER_81_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09322_ _08510_/B _09318_/X _09319_/X _09321_/X vssd1 vssd1 vccd1 vccd1 _09322_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_90_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_5_13_0_clk clkbuf_4_6_0_clk/X vssd1 vssd1 vccd1 vccd1 clkbuf_5_13_0_clk/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_22_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09253_ _14535_/Q _14148_/Q _14180_/Q _14116_/Q _09557_/S _09550_/A1 vssd1 vssd1
+ vccd1 vccd1 _09253_/X sky130_fd_sc_hd__mux4_1
XFILLER_21_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08204_ _13695_/Q _13333_/A0 _08216_/S vssd1 vssd1 vccd1 vccd1 _13695_/D sky130_fd_sc_hd__mux2_1
X_09184_ _14468_/Q _14436_/Q _13857_/Q _14210_/Q _09438_/S0 _09448_/S1 vssd1 vssd1
+ vccd1 vccd1 _09184_/X sky130_fd_sc_hd__mux4_2
X_08135_ _08093_/B _08133_/X _08134_/Y _08121_/X vssd1 vssd1 vccd1 vccd1 _08135_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_88_1023 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_5_28_0_clk clkbuf_5_29_0_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_5_28_0_clk/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_161_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08066_ _14759_/Q _13637_/Q _08066_/S vssd1 vssd1 vccd1 vccd1 _13637_/D sky130_fd_sc_hd__mux2_1
XFILLER_134_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07017_ _07016_/X _14738_/Q _07098_/S vssd1 vssd1 vccd1 vccd1 _13584_/D sky130_fd_sc_hd__mux2_1
XFILLER_162_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_251_clk clkbuf_5_1_0_clk/X vssd1 vssd1 vccd1 vccd1 _15108_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_88_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1040 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08968_ _09419_/A2 _08966_/X _08967_/X _09421_/A1 vssd1 vssd1 vccd1 vccd1 _08968_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_57_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07919_ _07921_/B _07918_/X _08012_/A2 vssd1 vssd1 vccd1 vccd1 _07919_/X sky130_fd_sc_hd__a21bo_1
XFILLER_112_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_1092 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08899_ _15108_/Q _15076_/Q _15649_/Q _13383_/Q _09132_/S _08988_/A1 vssd1 vssd1
+ vccd1 vccd1 _08899_/X sky130_fd_sc_hd__mux4_1
XFILLER_1_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10930_ _14948_/Q _10929_/B _10929_/Y _11521_/A vssd1 vssd1 vccd1 vccd1 _14948_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_95_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_64 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10861_ _14893_/Q _13775_/Q _12932_/S vssd1 vssd1 vccd1 vccd1 _14893_/D sky130_fd_sc_hd__mux2_1
XFILLER_13_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12600_ _14549_/Q _14162_/Q _14194_/Q _14130_/Q _12612_/S _12613_/A vssd1 vssd1 vccd1
+ vccd1 _12600_/X sky130_fd_sc_hd__mux4_1
XPHY_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13580_ _15620_/CLK _13580_/D vssd1 vssd1 vccd1 vccd1 _13580_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10792_ _14824_/Q _15456_/Q _12928_/S vssd1 vssd1 vccd1 vccd1 _14824_/D sky130_fd_sc_hd__mux2_1
XPHY_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12531_ _14546_/Q _14159_/Q _14191_/Q _14127_/Q _12612_/S _12613_/A vssd1 vssd1 vccd1
+ vccd1 _12531_/X sky130_fd_sc_hd__mux4_1
XPHY_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_74 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15250_ _15674_/CLK _15250_/D vssd1 vssd1 vccd1 vccd1 _15250_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_157_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12462_ _14543_/Q _14156_/Q _14188_/Q _14124_/Q _12472_/S _12465_/S1 vssd1 vssd1
+ vccd1 vccd1 _12462_/X sky130_fd_sc_hd__mux4_1
XFILLER_173_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14201_ _15211_/CLK _14201_/D vssd1 vssd1 vccd1 vccd1 _14201_/Q sky130_fd_sc_hd__dfxtp_1
X_11413_ _11412_/Y _15050_/Q _11641_/S vssd1 vssd1 vccd1 vccd1 _15050_/D sky130_fd_sc_hd__mux2_1
XFILLER_137_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15181_ _15181_/CLK _15181_/D vssd1 vssd1 vccd1 vccd1 _15181_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_166_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12393_ _14540_/Q _14153_/Q _14185_/Q _14121_/Q _12591_/S _12590_/A vssd1 vssd1 vccd1
+ vccd1 _12393_/X sky130_fd_sc_hd__mux4_1
X_14132_ _15650_/CLK _14132_/D vssd1 vssd1 vccd1 vccd1 _14132_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_181_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11344_ _11344_/A _11344_/B _11343_/X vssd1 vssd1 vccd1 vccd1 _11344_/X sky130_fd_sc_hd__or3b_1
XFILLER_125_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14063_ _15677_/CLK _14063_/D vssd1 vssd1 vccd1 vccd1 _14063_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_165_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11275_ _11329_/A _11329_/B vssd1 vssd1 vccd1 vccd1 _11275_/Y sky130_fd_sc_hd__nand2_1
X_13014_ _10694_/X _14885_/Q _13038_/S vssd1 vssd1 vccd1 vccd1 _13014_/X sky130_fd_sc_hd__mux2_4
X_10226_ input21/X _14611_/Q _13291_/S vssd1 vssd1 vccd1 vccd1 _14611_/D sky130_fd_sc_hd__mux2_1
XFILLER_79_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_242_clk clkbuf_5_5_0_clk/X vssd1 vssd1 vccd1 vccd1 _15657_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_67_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10157_ _14542_/Q _11876_/A1 _10159_/S vssd1 vssd1 vccd1 vccd1 _14542_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4 hold4/A vssd1 vssd1 vccd1 vccd1 hold4/X sky130_fd_sc_hd__bufbuf_16
XFILLER_66_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10088_ _14444_/Q _11874_/A1 _10097_/S vssd1 vssd1 vccd1 vccd1 _14444_/D sky130_fd_sc_hd__mux2_1
X_14965_ _15000_/CLK _14965_/D vssd1 vssd1 vccd1 vccd1 _14965_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13916_ _15497_/CLK _13916_/D vssd1 vssd1 vccd1 vccd1 _13916_/Q sky130_fd_sc_hd__dfxtp_1
X_14896_ _15208_/CLK _14896_/D vssd1 vssd1 vccd1 vccd1 _14896_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13847_ _15176_/CLK _13847_/D vssd1 vssd1 vccd1 vccd1 _13847_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_74_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13778_ _15398_/CLK _13778_/D vssd1 vssd1 vccd1 vccd1 _13778_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_188_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15517_ _15517_/CLK _15517_/D vssd1 vssd1 vccd1 vccd1 _15517_/Q sky130_fd_sc_hd__dfxtp_1
X_12729_ _12737_/A _12729_/B vssd1 vssd1 vccd1 vccd1 _12729_/X sky130_fd_sc_hd__or2_1
XFILLER_88_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15448_ _15634_/CLK _15448_/D vssd1 vssd1 vccd1 vccd1 _15448_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15379_ _15379_/CLK _15379_/D vssd1 vssd1 vccd1 vccd1 _15379_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_128_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_346 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09940_ _11860_/A1 _14300_/Q _09958_/S vssd1 vssd1 vccd1 vccd1 _14300_/D sky130_fd_sc_hd__mux2_1
XFILLER_131_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09871_ _11857_/A1 _14233_/Q _09897_/S vssd1 vssd1 vccd1 vccd1 _14233_/D sky130_fd_sc_hd__mux2_1
XFILLER_48_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_233_clk clkbuf_5_4_0_clk/X vssd1 vssd1 vccd1 vccd1 _14525_/CLK sky130_fd_sc_hd__clkbuf_16
X_08822_ _13845_/Q _13321_/A0 _08851_/S vssd1 vssd1 vccd1 vccd1 _13845_/D sky130_fd_sc_hd__mux2_1
XTAP_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_458 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08753_ _14589_/Q _14588_/Q _14587_/Q _08753_/D vssd1 vssd1 vccd1 vccd1 _08753_/X
+ sky130_fd_sc_hd__or4_1
X_07704_ _14745_/Q _07713_/A _07703_/Y _07949_/C1 vssd1 vssd1 vccd1 vccd1 _13488_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_94_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08684_ _13454_/Q _08684_/A2 _08693_/B1 _13621_/Q _08683_/X vssd1 vssd1 vccd1 vccd1
+ _08688_/B sky130_fd_sc_hd__a221o_1
XFILLER_38_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07635_ _13471_/Q _07635_/B vssd1 vssd1 vccd1 vccd1 _07636_/B sky130_fd_sc_hd__xnor2_1
XTAP_1908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07566_ _14741_/Q _07644_/A _07565_/X _12832_/C1 vssd1 vssd1 vccd1 vccd1 _13452_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_107_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09305_ _14376_/Q _15192_/Q _13831_/Q _14570_/Q _09481_/S _08519_/A vssd1 vssd1 vccd1
+ vccd1 _09306_/B sky130_fd_sc_hd__mux4_1
XFILLER_94_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07497_ _13349_/A0 _13413_/Q _07501_/S vssd1 vssd1 vccd1 vccd1 _13413_/D sky130_fd_sc_hd__mux2_1
XFILLER_10_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09236_ _09405_/A _09229_/X _09232_/X _09450_/B1 vssd1 vssd1 vccd1 vccd1 _09236_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_103_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09167_ _13888_/Q _09445_/A2 _09522_/B1 _14403_/Q _09437_/A1 vssd1 vssd1 vccd1 vccd1
+ _09167_/X sky130_fd_sc_hd__a221o_1
XFILLER_107_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08118_ _13656_/Q _10344_/S _08096_/X _08117_/X vssd1 vssd1 vccd1 vccd1 _13656_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_181_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09098_ _14366_/Q _15182_/Q _13821_/Q _14560_/Q _09444_/S _09446_/A1 vssd1 vssd1
+ vccd1 vccd1 _09099_/B sky130_fd_sc_hd__mux4_1
XFILLER_108_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08049_ _14742_/Q _13620_/Q _08066_/S vssd1 vssd1 vccd1 vccd1 _13620_/D sky130_fd_sc_hd__mux2_1
XFILLER_123_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11060_ _10958_/Y _10979_/B _11349_/A vssd1 vssd1 vccd1 vccd1 _11061_/A sky130_fd_sc_hd__mux2_1
XFILLER_27_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10011_ _13332_/A0 _14369_/Q _10028_/S vssd1 vssd1 vccd1 vccd1 _14369_/D sky130_fd_sc_hd__mux2_1
XFILLER_49_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_224_clk clkbuf_5_7_0_clk/X vssd1 vssd1 vccd1 vccd1 _15500_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_114_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14750_ _15608_/CLK _14750_/D vssd1 vssd1 vccd1 vccd1 _14750_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_3844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11962_ _12468_/A1 _11959_/X _12455_/C1 vssd1 vssd1 vccd1 vccd1 _11962_/X sky130_fd_sc_hd__o21a_1
XFILLER_28_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_86 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13701_ _15293_/CLK _13701_/D vssd1 vssd1 vccd1 vccd1 _13701_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10913_ _14939_/Q _10944_/B _10912_/Y _13183_/B vssd1 vssd1 vccd1 vccd1 _14939_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_56_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14681_ _15589_/CLK _14681_/D vssd1 vssd1 vccd1 vccd1 _14681_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11893_ _12500_/B1 _11890_/X _12501_/C1 vssd1 vssd1 vccd1 vccd1 _11893_/X sky130_fd_sc_hd__o21a_1
X_13632_ _13632_/CLK _13632_/D vssd1 vssd1 vccd1 vccd1 _13632_/Q sky130_fd_sc_hd__dfxtp_1
X_10844_ _14876_/Q _13792_/Q _12917_/S vssd1 vssd1 vccd1 vccd1 _14876_/D sky130_fd_sc_hd__mux2_1
X_13563_ _13565_/CLK _13563_/D vssd1 vssd1 vccd1 vccd1 _13563_/Q sky130_fd_sc_hd__dfxtp_2
X_10775_ _14807_/Q _15439_/Q _12918_/S vssd1 vssd1 vccd1 vccd1 _14807_/D sky130_fd_sc_hd__mux2_1
X_15302_ _15666_/CLK _15302_/D vssd1 vssd1 vccd1 vccd1 _15302_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12514_ _08405_/B _12511_/X _08405_/C vssd1 vssd1 vccd1 vccd1 _12514_/X sky130_fd_sc_hd__o21a_1
XFILLER_13_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13494_ _13632_/CLK _13494_/D vssd1 vssd1 vccd1 vccd1 _13494_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_158_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15233_ _15233_/CLK _15233_/D vssd1 vssd1 vccd1 vccd1 _15233_/Q sky130_fd_sc_hd__dfxtp_1
X_12445_ _12468_/A1 _12442_/X _12455_/C1 vssd1 vssd1 vccd1 vccd1 _12445_/X sky130_fd_sc_hd__o21a_1
XFILLER_173_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_72 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15164_ _15233_/CLK _15164_/D vssd1 vssd1 vccd1 vccd1 _15164_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_176_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12376_ _08405_/B _12373_/X _08405_/C vssd1 vssd1 vccd1 vccd1 _12376_/X sky130_fd_sc_hd__o21a_1
XFILLER_125_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14115_ _15665_/CLK _14115_/D vssd1 vssd1 vccd1 vccd1 _14115_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_125_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11327_ _11327_/A _11327_/B vssd1 vssd1 vccd1 vccd1 _11327_/X sky130_fd_sc_hd__or2_1
XFILLER_114_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15095_ _15668_/CLK _15095_/D vssd1 vssd1 vccd1 vccd1 _15095_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_125_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14046_ _15285_/CLK _14046_/D vssd1 vssd1 vccd1 vccd1 _14046_/Q sky130_fd_sc_hd__dfxtp_1
X_11258_ _11258_/A _11258_/B vssd1 vssd1 vccd1 vccd1 _11258_/Y sky130_fd_sc_hd__nor2_1
XFILLER_79_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_215_clk clkbuf_5_19_0_clk/X vssd1 vssd1 vccd1 vccd1 _15526_/CLK sky130_fd_sc_hd__clkbuf_16
X_10209_ input3/X hold8/A _13282_/S vssd1 vssd1 vccd1 vccd1 _14594_/D sky130_fd_sc_hd__mux2_1
XFILLER_39_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11189_ _11199_/A _11189_/B vssd1 vssd1 vccd1 vccd1 _11189_/Y sky130_fd_sc_hd__nor2_1
XFILLER_122_894 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14948_ _15577_/CLK _14948_/D vssd1 vssd1 vccd1 vccd1 _14948_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_480 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14879_ _15643_/CLK _14879_/D vssd1 vssd1 vccd1 vccd1 _14879_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07420_ _14745_/Q _07419_/X _07500_/S vssd1 vssd1 vccd1 vccd1 _07420_/X sky130_fd_sc_hd__mux2_8
XFILLER_63_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07351_ _07351_/A _07351_/B _07351_/C _07350_/X vssd1 vssd1 vccd1 vccd1 _07363_/B
+ sky130_fd_sc_hd__or4b_2
XFILLER_148_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07282_ _07278_/A _07278_/B _07280_/Y _07281_/X vssd1 vssd1 vccd1 vccd1 _07350_/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_148_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09021_ _13849_/Q _14202_/Q _09073_/S vssd1 vssd1 vccd1 vccd1 _09021_/X sky130_fd_sc_hd__mux2_1
XFILLER_117_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09923_ _11876_/A1 _14284_/Q _09925_/S vssd1 vssd1 vccd1 vccd1 _14284_/D sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_206_clk clkbuf_5_16_0_clk/X vssd1 vssd1 vccd1 vccd1 _15655_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_86_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09854_ _14218_/Q _11874_/A1 _09863_/S vssd1 vssd1 vccd1 vccd1 _14218_/D sky130_fd_sc_hd__mux2_1
XTAP_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08805_ _13339_/A0 _13831_/Q _08816_/S vssd1 vssd1 vccd1 vccd1 _13831_/D sky130_fd_sc_hd__mux2_1
XTAP_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09785_ _14152_/Q _13340_/A0 _09795_/S vssd1 vssd1 vccd1 vccd1 _14152_/D sky130_fd_sc_hd__mux2_1
XTAP_3107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06997_ _06997_/A _06997_/B _06997_/C vssd1 vssd1 vccd1 vccd1 _15540_/D sky130_fd_sc_hd__and3_1
XTAP_3118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08736_ _13415_/Q _08736_/A2 _08733_/X _08735_/X vssd1 vssd1 vccd1 vccd1 _08736_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_27_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_107 _15031_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_118 _07123_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_344 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_129 _08405_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08667_ _13123_/B _08724_/C _08668_/D vssd1 vssd1 vccd1 vccd1 _08667_/X sky130_fd_sc_hd__and3_2
XFILLER_121_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07618_ _07616_/X _07621_/B _07629_/A vssd1 vssd1 vccd1 vccd1 _07618_/X sky130_fd_sc_hd__a21bo_1
XFILLER_53_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08598_ _08722_/A _08598_/B _08598_/C vssd1 vssd1 vccd1 vccd1 _08598_/X sky130_fd_sc_hd__or3_1
XFILLER_26_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07549_ _13448_/Q _07549_/B vssd1 vssd1 vccd1 vccd1 _07549_/Y sky130_fd_sc_hd__nor2_1
XFILLER_139_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10560_ _14731_/Q _10559_/Y _10560_/S vssd1 vssd1 vccd1 vccd1 _14731_/D sky130_fd_sc_hd__mux2_1
X_09219_ _13922_/Q _09218_/X _12504_/A vssd1 vssd1 vccd1 vccd1 _13922_/D sky130_fd_sc_hd__mux2_1
XFILLER_127_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10491_ _10491_/A _13223_/B vssd1 vssd1 vccd1 vccd1 _10527_/B sky130_fd_sc_hd__and2_1
XFILLER_182_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12230_ _14243_/Q _14275_/Q _14307_/Q _14339_/Q _12499_/S _12486_/S1 vssd1 vssd1
+ vccd1 vccd1 _12230_/X sky130_fd_sc_hd__mux4_1
XFILLER_107_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_248 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12161_ _14240_/Q _14272_/Q _14304_/Q _14336_/Q _12246_/S _12268_/A vssd1 vssd1 vccd1
+ vccd1 _12161_/X sky130_fd_sc_hd__mux4_1
XFILLER_108_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11112_ _11053_/X _11061_/Y _11297_/S vssd1 vssd1 vccd1 vccd1 _11112_/X sky130_fd_sc_hd__mux2_1
XFILLER_2_955 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12092_ _14237_/Q _14269_/Q _14301_/Q _14333_/Q _12472_/S _12465_/S1 vssd1 vssd1
+ vccd1 vccd1 _12092_/X sky130_fd_sc_hd__mux4_1
XFILLER_89_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11043_ _11356_/B _11041_/Y _11042_/Y _11307_/A vssd1 vssd1 vccd1 vccd1 _11043_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_118_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_4_3_0_clk clkbuf_4_3_0_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_5_7_0_clk/A sky130_fd_sc_hd__clkbuf_8
XFILLER_76_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14802_ _15434_/CLK _14802_/D vssd1 vssd1 vccd1 vccd1 _14802_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12994_ _07440_/X _13024_/A2 _12993_/X _13024_/B2 vssd1 vssd1 vccd1 vccd1 _12994_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_91_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14733_ _15619_/CLK _14733_/D vssd1 vssd1 vccd1 vccd1 _14733_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11945_ _14005_/Q _13973_/Q _12543_/S vssd1 vssd1 vccd1 vccd1 _11946_/B sky130_fd_sc_hd__mux2_1
XFILLER_44_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14664_ _15635_/CLK _14664_/D vssd1 vssd1 vccd1 vccd1 _14664_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11876_ _15297_/Q _11876_/A1 _11878_/S vssd1 vssd1 vccd1 vccd1 _15297_/D sky130_fd_sc_hd__mux2_1
XTAP_2984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13615_ _13803_/CLK _13615_/D vssd1 vssd1 vccd1 vccd1 _13615_/Q sky130_fd_sc_hd__dfxtp_1
X_10827_ _14859_/Q _07228_/A _12906_/S vssd1 vssd1 vccd1 vccd1 _14859_/D sky130_fd_sc_hd__mux2_1
X_14595_ _15536_/CLK _14595_/D vssd1 vssd1 vccd1 vccd1 _14595_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_186_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_1080 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13546_ _15399_/CLK _13546_/D vssd1 vssd1 vccd1 vccd1 _13546_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_186_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_555 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10758_ _15422_/Q _14790_/Q _10759_/S vssd1 vssd1 vccd1 vccd1 _14790_/D sky130_fd_sc_hd__mux2_1
XFILLER_186_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13477_ _15542_/CLK _13477_/D vssd1 vssd1 vccd1 vccd1 _13477_/Q sky130_fd_sc_hd__dfxtp_2
X_10689_ _15065_/Q _10714_/A2 _10686_/X _10688_/X vssd1 vssd1 vccd1 vccd1 _10689_/X
+ sky130_fd_sc_hd__o22a_2
X_15216_ _15220_/CLK _15216_/D vssd1 vssd1 vccd1 vccd1 _15216_/Q sky130_fd_sc_hd__dfxtp_1
X_12428_ _14026_/Q _13994_/Q _12430_/S vssd1 vssd1 vccd1 vccd1 _12429_/B sky130_fd_sc_hd__mux2_1
XFILLER_127_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15147_ _15220_/CLK _15147_/D vssd1 vssd1 vccd1 vccd1 _15147_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12359_ _14023_/Q _13991_/Q _12541_/S vssd1 vssd1 vccd1 vccd1 _12360_/B sky130_fd_sc_hd__mux2_1
XFILLER_153_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15078_ _15651_/CLK _15078_/D vssd1 vssd1 vccd1 vccd1 _15078_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06920_ _06920_/A _06920_/B _06918_/X vssd1 vssd1 vccd1 vccd1 _06922_/B sky130_fd_sc_hd__or3b_2
XFILLER_141_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14029_ _15088_/CLK _14029_/D vssd1 vssd1 vccd1 vccd1 _14029_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06851_ _06851_/A _06851_/B vssd1 vssd1 vccd1 vccd1 _06997_/A sky130_fd_sc_hd__nor2_1
XFILLER_68_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09570_ _13946_/Q _13326_/A0 _09589_/S vssd1 vssd1 vccd1 vccd1 _13946_/D sky130_fd_sc_hd__mux2_1
X_06782_ _06782_/A _10735_/S _06782_/C vssd1 vssd1 vccd1 vccd1 _06782_/Y sky130_fd_sc_hd__nand3_2
XFILLER_36_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08521_ _08521_/A _08529_/B vssd1 vssd1 vccd1 vccd1 _08521_/Y sky130_fd_sc_hd__nor2_8
XFILLER_36_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08452_ _13756_/Q _12910_/S _08426_/X _08451_/X vssd1 vssd1 vccd1 vccd1 _13756_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_51_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07403_ _13656_/Q _07499_/A2 _07499_/B1 _14684_/Q _07402_/X vssd1 vssd1 vccd1 vccd1
+ _07403_/X sky130_fd_sc_hd__a221o_1
XFILLER_168_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08383_ _08244_/A _13759_/Q _15413_/Q _08244_/B vssd1 vssd1 vccd1 vccd1 _08383_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_32_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07334_ _13909_/Q _15496_/Q _07334_/S vssd1 vssd1 vccd1 vccd1 _07337_/A sky130_fd_sc_hd__mux2_8
XFILLER_91_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_1096 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07265_ _07265_/A _07265_/B vssd1 vssd1 vccd1 vccd1 _07273_/B sky130_fd_sc_hd__or2_1
X_09004_ _09523_/A1 _09002_/X _09003_/X vssd1 vssd1 vccd1 vccd1 _09008_/B sky130_fd_sc_hd__a21o_1
X_07196_ _15337_/Q _15493_/Q _07335_/S vssd1 vssd1 vccd1 vccd1 _07197_/B sky130_fd_sc_hd__mux2_8
XFILLER_105_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout500 _08240_/A vssd1 vssd1 vccd1 vccd1 _10520_/A1 sky130_fd_sc_hd__buf_6
XFILLER_133_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout511 _14607_/Q vssd1 vssd1 vccd1 vccd1 _06676_/A sky130_fd_sc_hd__buf_12
XFILLER_132_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09906_ _12967_/A1 _14267_/Q _09925_/S vssd1 vssd1 vccd1 vccd1 _14267_/D sky130_fd_sc_hd__mux2_1
Xfanout522 _09466_/A vssd1 vssd1 vccd1 vccd1 _09532_/A sky130_fd_sc_hd__buf_12
Xfanout533 _08487_/A vssd1 vssd1 vccd1 vccd1 _09448_/S1 sky130_fd_sc_hd__buf_12
XFILLER_24_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout544 _09425_/S vssd1 vssd1 vccd1 vccd1 _09225_/S0 sky130_fd_sc_hd__buf_12
XFILLER_76_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout555 _08490_/A1 vssd1 vssd1 vccd1 vccd1 _09521_/S sky130_fd_sc_hd__buf_12
XFILLER_58_222 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout566 _14603_/Q vssd1 vssd1 vccd1 vccd1 _08490_/A1 sky130_fd_sc_hd__buf_12
X_09837_ _14201_/Q _11649_/A0 _09863_/S vssd1 vssd1 vccd1 vccd1 _14201_/D sky130_fd_sc_hd__mux2_1
XTAP_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout577 _08453_/A vssd1 vssd1 vccd1 vccd1 _12468_/A1 sky130_fd_sc_hd__buf_12
XFILLER_47_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout588 _12061_/A vssd1 vssd1 vccd1 vccd1 _12452_/A sky130_fd_sc_hd__clkbuf_16
XTAP_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout599 fanout600/X vssd1 vssd1 vccd1 vccd1 _12613_/A sky130_fd_sc_hd__buf_6
XFILLER_86_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09768_ _14135_/Q _11681_/A0 _09790_/S vssd1 vssd1 vccd1 vccd1 _14135_/D sky130_fd_sc_hd__mux2_1
XFILLER_73_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08719_ _13545_/Q _08747_/A2 _08747_/B1 _13481_/Q vssd1 vssd1 vccd1 vccd1 _08719_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_2225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09699_ _11854_/A1 _14069_/Q _09728_/S vssd1 vssd1 vccd1 vccd1 _14069_/D sky130_fd_sc_hd__mux2_1
XTAP_2236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_826 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11730_ _15159_/Q _11838_/A1 _11742_/S vssd1 vssd1 vccd1 vccd1 _15159_/D sky130_fd_sc_hd__mux2_1
XTAP_1524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_656 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11661_ _13336_/A0 _15093_/Q _11675_/S vssd1 vssd1 vccd1 vccd1 _15093_/D sky130_fd_sc_hd__mux2_1
XTAP_1579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13400_ _15666_/CLK _13400_/D vssd1 vssd1 vccd1 vccd1 _13400_/Q sky130_fd_sc_hd__dfxtp_1
X_10612_ _15560_/Q _10731_/B _10733_/B1 _14937_/Q vssd1 vssd1 vccd1 vccd1 _10612_/X
+ sky130_fd_sc_hd__a22o_1
X_14380_ _15303_/CLK _14380_/D vssd1 vssd1 vccd1 vccd1 _14380_/Q sky130_fd_sc_hd__dfxtp_1
X_11592_ _13233_/B _11593_/B vssd1 vssd1 vccd1 vccd1 _11606_/A sky130_fd_sc_hd__and2_1
XFILLER_167_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13331_ _13331_/A0 _15661_/Q _13345_/S vssd1 vssd1 vccd1 vccd1 _15661_/D sky130_fd_sc_hd__mux2_1
X_10543_ _10527_/B _10543_/B _10543_/C vssd1 vssd1 vccd1 vccd1 _10543_/X sky130_fd_sc_hd__and3b_1
XFILLER_167_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13262_ _15346_/Q _15593_/Q _13300_/S vssd1 vssd1 vccd1 vccd1 _15593_/D sky130_fd_sc_hd__mux2_1
XFILLER_109_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10474_ _10507_/A1 _13751_/Q _15421_/Q _08244_/B vssd1 vssd1 vccd1 vccd1 _10474_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_109_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15001_ _15584_/CLK _15001_/D vssd1 vssd1 vccd1 vccd1 _15001_/Q sky130_fd_sc_hd__dfxtp_1
X_12213_ _15287_/Q _15255_/Q _15223_/Q _15154_/Q _12489_/S0 _12489_/S1 vssd1 vssd1
+ vccd1 vccd1 _12214_/B sky130_fd_sc_hd__mux4_1
XFILLER_182_388 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13193_ _06769_/Y _11457_/A _11475_/B _13192_/Y vssd1 vssd1 vccd1 vccd1 _13193_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_29_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12144_ _15284_/Q _15252_/Q _15220_/Q _15151_/Q _12154_/S _12253_/S1 vssd1 vssd1
+ vccd1 vccd1 _12145_/B sky130_fd_sc_hd__mux4_1
XFILLER_124_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12075_ _15281_/Q _15249_/Q _15217_/Q _15148_/Q _12470_/S _12080_/A vssd1 vssd1 vccd1
+ vccd1 _12076_/B sky130_fd_sc_hd__mux4_1
XFILLER_1_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11026_ _11037_/A _11563_/A vssd1 vssd1 vccd1 vccd1 _11294_/B sky130_fd_sc_hd__nand2_1
XFILLER_38_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12977_ _15472_/Q _13105_/A2 _13025_/B1 _12976_/X vssd1 vssd1 vccd1 vccd1 _15472_/D
+ sky130_fd_sc_hd__a22o_1
XTAP_3471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11928_ _12618_/A1 _11927_/X _11926_/X _12618_/C1 vssd1 vssd1 vccd1 vccd1 _11929_/C
+ sky130_fd_sc_hd__a211o_1
X_14716_ _15525_/CLK _14716_/D vssd1 vssd1 vccd1 vccd1 _14716_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_2770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14647_ _15618_/CLK _14647_/D vssd1 vssd1 vccd1 vccd1 _14647_/Q sky130_fd_sc_hd__dfxtp_1
X_11859_ _15280_/Q _12967_/A1 _11878_/S vssd1 vssd1 vccd1 vccd1 _15280_/D sky130_fd_sc_hd__mux2_1
XFILLER_159_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_18 _15073_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_29 _14748_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14578_ _15200_/CLK _14578_/D vssd1 vssd1 vccd1 vccd1 _14578_/Q sky130_fd_sc_hd__dfxtp_1
X_13529_ _13632_/CLK _13529_/D vssd1 vssd1 vccd1 vccd1 _13529_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_159_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07050_ _07049_/X _14749_/Q _07077_/S vssd1 vssd1 vccd1 vccd1 _13595_/D sky130_fd_sc_hd__mux2_1
XFILLER_174_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07952_ _14746_/Q _07964_/A _07951_/Y _07965_/C1 vssd1 vssd1 vccd1 vccd1 _13553_/D
+ sky130_fd_sc_hd__o211a_1
X_06903_ _15377_/Q _07571_/A _15376_/Q _07571_/B _06902_/X vssd1 vssd1 vccd1 vccd1
+ _06903_/X sky130_fd_sc_hd__o221a_1
X_07883_ _14760_/Q _07903_/A _07882_/Y _08012_/C1 vssd1 vssd1 vccd1 vccd1 _13535_/D
+ sky130_fd_sc_hd__o211a_1
X_09622_ _13996_/Q _13344_/A0 _09627_/S vssd1 vssd1 vccd1 vccd1 _13996_/D sky130_fd_sc_hd__mux2_1
XFILLER_83_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06834_ _09382_/A _06834_/B vssd1 vssd1 vccd1 vccd1 _06834_/Y sky130_fd_sc_hd__nand2_1
XFILLER_55_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09553_ _09553_/A1 _09551_/X _09552_/X vssd1 vssd1 vccd1 vccd1 _09554_/C sky130_fd_sc_hd__a21o_1
X_06765_ input24/X vssd1 vssd1 vccd1 vccd1 _06765_/Y sky130_fd_sc_hd__inv_2
XFILLER_71_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08504_ _13125_/B _14608_/Q _14610_/Q _14609_/Q vssd1 vssd1 vccd1 vccd1 _08517_/A
+ sky130_fd_sc_hd__or4_4
XFILLER_24_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09484_ _14031_/Q _13999_/Q _09484_/S vssd1 vssd1 vccd1 vccd1 _09484_/X sky130_fd_sc_hd__mux2_1
XFILLER_23_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06696_ _13473_/Q vssd1 vssd1 vccd1 vccd1 _06696_/Y sky130_fd_sc_hd__inv_2
XFILLER_24_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_628 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_144 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08435_ _14609_/Q _08390_/C _08425_/X _10764_/S vssd1 vssd1 vccd1 vccd1 _08435_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_178_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08366_ _08366_/A vssd1 vssd1 vccd1 vccd1 _08366_/Y sky130_fd_sc_hd__inv_2
XFILLER_149_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07317_ _07317_/A vssd1 vssd1 vccd1 vccd1 _07352_/B sky130_fd_sc_hd__inv_2
XFILLER_177_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08297_ _11088_/S _08280_/Y _08296_/X vssd1 vssd1 vccd1 vccd1 _08298_/B sky130_fd_sc_hd__o21ai_2
XFILLER_137_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07248_ _07248_/A vssd1 vssd1 vccd1 vccd1 _07260_/B sky130_fd_sc_hd__inv_2
XFILLER_178_1046 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07179_ _15353_/Q _15060_/Q _07188_/S vssd1 vssd1 vccd1 vccd1 _07179_/X sky130_fd_sc_hd__mux2_8
XFILLER_127_44 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_88 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10190_ _11876_/A1 _14574_/Q _10192_/S vssd1 vssd1 vccd1 vccd1 _14574_/D sky130_fd_sc_hd__mux2_1
XFILLER_87_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout330 _07412_/X vssd1 vssd1 vccd1 vccd1 _13328_/A0 sky130_fd_sc_hd__buf_8
Xfanout341 _07392_/X vssd1 vssd1 vccd1 vccd1 _11681_/A0 sky130_fd_sc_hd__buf_6
Xfanout352 _10602_/B vssd1 vssd1 vccd1 vccd1 _10652_/B sky130_fd_sc_hd__buf_8
XFILLER_120_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout363 _09522_/B1 vssd1 vssd1 vccd1 vccd1 _09403_/B1 sky130_fd_sc_hd__buf_12
XFILLER_143_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout374 _08242_/X vssd1 vssd1 vccd1 vccd1 _11349_/B sky130_fd_sc_hd__buf_8
XFILLER_115_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout385 _08236_/X vssd1 vssd1 vccd1 vccd1 _11252_/A sky130_fd_sc_hd__buf_8
XFILLER_4_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12900_ _15428_/Q _15613_/Q _12900_/S vssd1 vssd1 vccd1 vccd1 _15428_/D sky130_fd_sc_hd__mux2_1
Xfanout396 _11129_/A vssd1 vssd1 vccd1 vccd1 _11283_/A sky130_fd_sc_hd__buf_8
XFILLER_74_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13880_ _15081_/CLK _13880_/D vssd1 vssd1 vccd1 vccd1 _13880_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12831_ _06861_/Y _12828_/X _12829_/X _12830_/X vssd1 vssd1 vccd1 vccd1 _12831_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_36_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15550_ _15648_/CLK _15550_/D vssd1 vssd1 vccd1 vccd1 _15550_/Q sky130_fd_sc_hd__dfxtp_1
X_12762_ _15064_/Q _12761_/X _12792_/B vssd1 vssd1 vccd1 vccd1 _12762_/X sky130_fd_sc_hd__mux2_1
XFILLER_36_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14501_ _15383_/CLK _14501_/D vssd1 vssd1 vccd1 vccd1 _14501_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11713_ _15142_/Q _11854_/A1 _11742_/S vssd1 vssd1 vccd1 vccd1 _15142_/D sky130_fd_sc_hd__mux2_1
XTAP_1354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15481_ _15525_/CLK _15481_/D vssd1 vssd1 vccd1 vccd1 _15481_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12693_ _12737_/A _12693_/B vssd1 vssd1 vccd1 vccd1 _12693_/X sky130_fd_sc_hd__or2_1
XTAP_1365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_436 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14432_ _15556_/CLK _14432_/D vssd1 vssd1 vccd1 vccd1 _14432_/Q sky130_fd_sc_hd__dfxtp_1
X_11644_ _13319_/A0 _15076_/Q _11670_/S vssd1 vssd1 vccd1 vccd1 _15076_/D sky130_fd_sc_hd__mux2_1
XFILLER_52_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14363_ _15220_/CLK _14363_/D vssd1 vssd1 vccd1 vccd1 _14363_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_122_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_1083 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11575_ _11573_/Y _11574_/X _15066_/Q _11614_/S vssd1 vssd1 vccd1 vccd1 _15066_/D
+ sky130_fd_sc_hd__a2bb2o_1
Xinput16 ext_read_data[23] vssd1 vssd1 vccd1 vccd1 input16/X sky130_fd_sc_hd__buf_8
XFILLER_122_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput27 ext_read_data[4] vssd1 vssd1 vccd1 vccd1 input27/X sky130_fd_sc_hd__clkbuf_8
XFILLER_155_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_884 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13314_ _15645_/Q _12821_/B _13316_/S vssd1 vssd1 vccd1 vccd1 _15645_/D sky130_fd_sc_hd__mux2_1
X_10526_ _10524_/X _10526_/B vssd1 vssd1 vccd1 vccd1 _10527_/D sky130_fd_sc_hd__nand2b_1
XFILLER_182_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14294_ _15211_/CLK _14294_/D vssd1 vssd1 vccd1 vccd1 _14294_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13245_ _13217_/A _11626_/A _11624_/A vssd1 vssd1 vccd1 vccd1 _13245_/X sky130_fd_sc_hd__o21a_1
X_10457_ _07213_/X _10457_/A2 _10456_/X vssd1 vssd1 vccd1 vccd1 _11610_/A sky130_fd_sc_hd__a21o_4
XFILLER_184_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13176_ _15559_/Q _13252_/B _13174_/Y _13175_/X vssd1 vssd1 vccd1 vccd1 _15559_/D
+ sky130_fd_sc_hd__a22o_1
X_10388_ _11440_/A _11476_/B vssd1 vssd1 vccd1 vccd1 _10389_/B sky130_fd_sc_hd__or2_1
XFILLER_151_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12127_ _13885_/Q _14400_/Q _12476_/S vssd1 vssd1 vccd1 vccd1 _12127_/X sky130_fd_sc_hd__mux2_1
XFILLER_96_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12058_ _13882_/Q _14397_/Q _12246_/S vssd1 vssd1 vccd1 vccd1 _12058_/X sky130_fd_sc_hd__mux2_1
XFILLER_84_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_203 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11009_ _11013_/A _13236_/B vssd1 vssd1 vccd1 vccd1 _11324_/B sky130_fd_sc_hd__nand2_1
XFILLER_93_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15679_ _15679_/CLK _15679_/D vssd1 vssd1 vccd1 vccd1 _15679_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08220_ _13711_/Q _11816_/A1 _08221_/S vssd1 vssd1 vccd1 vccd1 _13711_/D sky130_fd_sc_hd__mux2_1
X_08151_ _08150_/X _08185_/B _08151_/S vssd1 vssd1 vccd1 vccd1 _08151_/X sky130_fd_sc_hd__mux2_2
XFILLER_158_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_631 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07102_ _15043_/Q _08121_/A vssd1 vssd1 vccd1 vccd1 _07103_/B sky130_fd_sc_hd__or2_1
XFILLER_173_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08082_ _13646_/Q _12647_/B _08081_/X vssd1 vssd1 vccd1 vccd1 _08083_/B sky130_fd_sc_hd__o21ai_1
XFILLER_134_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07033_ _14623_/Q _14655_/Q _07078_/S vssd1 vssd1 vccd1 vccd1 _07033_/X sky130_fd_sc_hd__mux2_1
XFILLER_161_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08984_ _08988_/A1 _08982_/X _08983_/X vssd1 vssd1 vccd1 vccd1 _08985_/C sky130_fd_sc_hd__a21o_1
XFILLER_87_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07935_ _13549_/Q _13548_/Q _13547_/Q _07935_/D vssd1 vssd1 vccd1 vccd1 _07946_/D
+ sky130_fd_sc_hd__and4_2
XFILLER_87_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07866_ _13531_/Q _07866_/B vssd1 vssd1 vccd1 vccd1 _07866_/X sky130_fd_sc_hd__xor2_1
XFILLER_29_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09605_ _13979_/Q _13327_/A0 _09627_/S vssd1 vssd1 vccd1 vccd1 _13979_/D sky130_fd_sc_hd__mux2_1
X_06817_ _13732_/Q _06817_/B vssd1 vssd1 vccd1 vccd1 _06817_/X sky130_fd_sc_hd__or2_1
XFILLER_113_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07797_ _14737_/Q _07816_/A _07796_/Y _08084_/C1 vssd1 vssd1 vccd1 vccd1 _13512_/D
+ sky130_fd_sc_hd__o211a_1
X_09536_ _14484_/Q _09536_/A2 _13130_/B1 _14452_/Q _06676_/A vssd1 vssd1 vccd1 vccd1
+ _09536_/X sky130_fd_sc_hd__a221o_1
XFILLER_71_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06748_ _13480_/Q vssd1 vssd1 vccd1 vccd1 _06748_/Y sky130_fd_sc_hd__inv_2
XFILLER_145_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09467_ _13123_/A _09464_/X _09466_/X _09382_/A vssd1 vssd1 vccd1 vccd1 _09467_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_52_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06679_ _14908_/Q vssd1 vssd1 vccd1 vccd1 _06834_/B sky130_fd_sc_hd__inv_2
XFILLER_12_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08418_ _14928_/D _08417_/X _12504_/A vssd1 vssd1 vccd1 vccd1 _13741_/D sky130_fd_sc_hd__mux2_1
X_09398_ _09421_/A1 _09394_/X _09397_/X _09393_/X vssd1 vssd1 vccd1 vccd1 _09411_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_178_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08349_ _08274_/X _08320_/Y _08348_/X _11283_/A vssd1 vssd1 vccd1 vccd1 _08349_/X
+ sky130_fd_sc_hd__a22o_2
XFILLER_149_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11360_ _11360_/A _11360_/B vssd1 vssd1 vccd1 vccd1 _11360_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_164_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10311_ _14696_/Q _14881_/Q _10715_/S vssd1 vssd1 vccd1 vccd1 _14696_/D sky130_fd_sc_hd__mux2_1
X_11291_ _11347_/A _11289_/X _08233_/B vssd1 vssd1 vccd1 vccd1 _11291_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_180_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_47 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13030_ _07488_/X _13039_/A2 _13029_/X _12944_/A vssd1 vssd1 vccd1 vccd1 _13030_/X
+ sky130_fd_sc_hd__a22o_1
X_10242_ _14627_/Q _14780_/Q _10630_/S vssd1 vssd1 vccd1 vccd1 _14627_/D sky130_fd_sc_hd__mux2_1
XFILLER_106_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10173_ _12967_/A1 _14557_/Q _10192_/S vssd1 vssd1 vccd1 vccd1 _14557_/D sky130_fd_sc_hd__mux2_1
XFILLER_66_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout160 _08626_/S vssd1 vssd1 vccd1 vccd1 _12929_/S sky130_fd_sc_hd__buf_12
XFILLER_102_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14981_ _15581_/CLK _14981_/D vssd1 vssd1 vccd1 vccd1 _14981_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout171 _11785_/Y vssd1 vssd1 vccd1 vccd1 _11816_/S sky130_fd_sc_hd__buf_12
XFILLER_47_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout182 _10132_/Y vssd1 vssd1 vccd1 vccd1 _10164_/S sky130_fd_sc_hd__buf_12
XFILLER_102_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout193 _09931_/Y vssd1 vssd1 vccd1 vccd1 _09958_/S sky130_fd_sc_hd__buf_12
X_13932_ _15315_/CLK _13932_/D vssd1 vssd1 vccd1 vccd1 _13932_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_19_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13863_ _15669_/CLK _13863_/D vssd1 vssd1 vccd1 vccd1 _13863_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15602_ _15643_/CLK _15602_/D vssd1 vssd1 vccd1 vccd1 _15602_/Q sky130_fd_sc_hd__dfxtp_1
X_12814_ _15071_/Q _12834_/B vssd1 vssd1 vccd1 vccd1 _12814_/X sky130_fd_sc_hd__or2_1
X_13794_ _15592_/CLK _13794_/D vssd1 vssd1 vccd1 vccd1 _13794_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_188_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12745_ _15355_/Q _15354_/Q _12745_/C vssd1 vssd1 vccd1 vccd1 _12754_/B sky130_fd_sc_hd__and3_1
XTAP_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15533_ _15648_/CLK _15533_/D vssd1 vssd1 vccd1 vccd1 _15533_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_767 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_907 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15464_ _15527_/CLK _15464_/D vssd1 vssd1 vccd1 vccd1 _15464_/Q sky130_fd_sc_hd__dfxtp_1
X_12676_ _13422_/Q _12675_/X _12728_/S vssd1 vssd1 vccd1 vccd1 _12677_/B sky130_fd_sc_hd__mux2_1
XFILLER_30_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14415_ _14415_/CLK _14415_/D vssd1 vssd1 vccd1 vccd1 _14415_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11627_ _11625_/Y _11627_/B vssd1 vssd1 vccd1 vccd1 _11629_/A sky130_fd_sc_hd__nand2b_1
X_15395_ _15397_/CLK _15395_/D vssd1 vssd1 vccd1 vccd1 _15395_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14346_ _15295_/CLK _14346_/D vssd1 vssd1 vccd1 vccd1 _14346_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_184_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11558_ _11542_/A _11548_/Y _11576_/B _11614_/S vssd1 vssd1 vccd1 vccd1 _11558_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_144_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10509_ _13218_/A _13217_/B vssd1 vssd1 vccd1 vccd1 _10541_/A sky130_fd_sc_hd__and2b_1
X_14277_ _15125_/CLK _14277_/D vssd1 vssd1 vccd1 vccd1 _14277_/Q sky130_fd_sc_hd__dfxtp_1
X_11489_ _11491_/B _11491_/C _13202_/B vssd1 vssd1 vccd1 vccd1 _11492_/A sky130_fd_sc_hd__a21oi_1
XFILLER_6_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_1102 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13228_ _13226_/Y _13227_/X _15576_/Q _13252_/B vssd1 vssd1 vccd1 vccd1 _15576_/D
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_112_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13159_ _13251_/A _13159_/B vssd1 vssd1 vccd1 vccd1 _13159_/Y sky130_fd_sc_hd__nand2_1
XFILLER_33_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07720_ _13493_/Q _07724_/C vssd1 vssd1 vccd1 vccd1 _07721_/B sky130_fd_sc_hd__xnor2_1
X_07651_ _07651_/A _07651_/B vssd1 vssd1 vccd1 vccd1 _07651_/Y sky130_fd_sc_hd__nand2_1
XFILLER_65_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07582_ _14745_/Q _07607_/A _07581_/Y _12809_/C1 vssd1 vssd1 vccd1 vccd1 _13456_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_92_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09321_ _15128_/Q _09558_/A2 _13130_/C1 _09320_/X vssd1 vssd1 vccd1 vccd1 _09321_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_40_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_570 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09252_ _09524_/A _09252_/B _09252_/C vssd1 vssd1 vccd1 vccd1 _09252_/X sky130_fd_sc_hd__and3_1
X_08203_ _13694_/Q _13078_/B2 _08216_/S vssd1 vssd1 vccd1 vccd1 _13694_/D sky130_fd_sc_hd__mux2_1
XFILLER_18_1070 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09183_ _09437_/A1 _09182_/X _09181_/X _09405_/A vssd1 vssd1 vccd1 vccd1 _09183_/X
+ sky130_fd_sc_hd__o211a_1
X_08134_ _08133_/S _06762_/Y _08151_/S vssd1 vssd1 vccd1 vccd1 _08134_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_146_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08065_ _14758_/Q _13636_/Q _08066_/S vssd1 vssd1 vccd1 vccd1 _13636_/D sky130_fd_sc_hd__mux2_1
XFILLER_174_494 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_859 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07016_ _07015_/X _13584_/Q _12640_/S vssd1 vssd1 vccd1 vccd1 _07016_/X sky130_fd_sc_hd__mux2_1
XFILLER_89_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08967_ _14521_/Q _14134_/Q _14166_/Q _14102_/Q _09047_/S _09530_/S1 vssd1 vssd1
+ vccd1 vccd1 _08967_/X sky130_fd_sc_hd__mux4_1
XFILLER_48_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_1052 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07918_ _13544_/Q _07924_/D vssd1 vssd1 vccd1 vccd1 _07918_/X sky130_fd_sc_hd__or2_1
XFILLER_25_1074 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08898_ _09234_/S1 _08896_/X _08897_/X vssd1 vssd1 vccd1 vccd1 _08898_/X sky130_fd_sc_hd__a21o_1
XFILLER_56_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07849_ _07858_/D _07848_/Y _07830_/A vssd1 vssd1 vccd1 vccd1 _07849_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_72_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10860_ _14892_/Q _13776_/Q _12885_/S vssd1 vssd1 vccd1 vccd1 _14892_/D sky130_fd_sc_hd__mux2_1
XFILLER_17_76 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_66 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09519_ _13905_/Q _09522_/A2 _09519_/B1 _14420_/Q _08507_/A vssd1 vssd1 vccd1 vccd1
+ _09519_/X sky130_fd_sc_hd__a221o_1
XPHY_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10791_ _14823_/Q hold9/X _12927_/S vssd1 vssd1 vccd1 vccd1 _14823_/D sky130_fd_sc_hd__mux2_1
XFILLER_24_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12530_ _14482_/Q _14450_/Q _13871_/Q _14224_/Q _12612_/S _12613_/A vssd1 vssd1 vccd1
+ vccd1 _12530_/X sky130_fd_sc_hd__mux4_1
XPHY_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12461_ _14479_/Q _14447_/Q _13868_/Q _14221_/Q _12489_/S0 _12489_/S1 vssd1 vssd1
+ vccd1 vccd1 _12461_/X sky130_fd_sc_hd__mux4_1
XFILLER_33_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14200_ _15176_/CLK _14200_/D vssd1 vssd1 vccd1 vccd1 _14200_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11412_ _11423_/D _11412_/B vssd1 vssd1 vccd1 vccd1 _11412_/Y sky130_fd_sc_hd__xnor2_1
X_15180_ _15279_/CLK _15180_/D vssd1 vssd1 vccd1 vccd1 _15180_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_126_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12392_ _14476_/Q _14444_/Q _13865_/Q _14218_/Q _12591_/S _12590_/A vssd1 vssd1 vccd1
+ vccd1 _12392_/X sky130_fd_sc_hd__mux4_1
XFILLER_165_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14131_ _15108_/CLK _14131_/D vssd1 vssd1 vccd1 vccd1 _14131_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_165_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11343_ _11329_/A _11289_/X _11318_/X _11048_/Y vssd1 vssd1 vccd1 vccd1 _11343_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_4_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14062_ _15676_/CLK _14062_/D vssd1 vssd1 vccd1 vccd1 _14062_/Q sky130_fd_sc_hd__dfxtp_1
X_11274_ _11243_/X _11273_/X _11297_/S vssd1 vssd1 vccd1 vccd1 _11329_/B sky130_fd_sc_hd__mux2_1
XFILLER_98_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13013_ _15484_/Q _10877_/S _13116_/C _13012_/X vssd1 vssd1 vccd1 vccd1 _15484_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_134_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10225_ input20/X _14610_/Q _13284_/S vssd1 vssd1 vccd1 vccd1 _14610_/D sky130_fd_sc_hd__mux2_1
XFILLER_67_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10156_ _14541_/Q _13342_/A0 _10164_/S vssd1 vssd1 vccd1 vccd1 _14541_/D sky130_fd_sc_hd__mux2_1
XFILLER_94_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5 hold5/A vssd1 vssd1 vccd1 vccd1 hold5/X sky130_fd_sc_hd__bufbuf_16
X_10087_ _14443_/Q _13340_/A0 _10097_/S vssd1 vssd1 vccd1 vccd1 _14443_/D sky130_fd_sc_hd__mux2_1
X_14964_ _14966_/CLK _14964_/D vssd1 vssd1 vccd1 vccd1 _14964_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13915_ _15510_/CLK _13915_/D vssd1 vssd1 vccd1 vccd1 _13915_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14895_ _15530_/CLK _14895_/D vssd1 vssd1 vccd1 vccd1 _14895_/Q sky130_fd_sc_hd__dfxtp_1
X_13846_ _15244_/CLK _13846_/D vssd1 vssd1 vccd1 vccd1 _13846_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13777_ _15397_/CLK _13777_/D vssd1 vssd1 vccd1 vccd1 _13777_/Q sky130_fd_sc_hd__dfxtp_4
X_10989_ _11037_/A _13202_/B vssd1 vssd1 vccd1 vccd1 _11242_/B sky130_fd_sc_hd__and2_1
XFILLER_43_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15516_ _15517_/CLK _15516_/D vssd1 vssd1 vccd1 vccd1 _15516_/Q sky130_fd_sc_hd__dfxtp_1
X_12728_ _13429_/Q _12727_/X _12728_/S vssd1 vssd1 vccd1 vccd1 _12729_/B sky130_fd_sc_hd__mux2_1
XFILLER_175_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15447_ _15447_/CLK _15447_/D vssd1 vssd1 vccd1 vccd1 hold2/A sky130_fd_sc_hd__dfxtp_1
XFILLER_175_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12659_ _12666_/B _12659_/B vssd1 vssd1 vccd1 vccd1 _12659_/Y sky130_fd_sc_hd__nor2_1
XFILLER_157_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15378_ _15378_/CLK _15378_/D vssd1 vssd1 vccd1 vccd1 _15378_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_184_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14329_ _15278_/CLK _14329_/D vssd1 vssd1 vccd1 vccd1 _14329_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09870_ _13323_/A0 _14232_/Q _09892_/S vssd1 vssd1 vccd1 vccd1 _14232_/D sky130_fd_sc_hd__mux2_1
XTAP_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08821_ _13844_/Q _13320_/A0 _08851_/S vssd1 vssd1 vccd1 vccd1 _13844_/D sky130_fd_sc_hd__mux2_1
XTAP_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08752_ _13806_/Q _12900_/S _08751_/X vssd1 vssd1 vccd1 vccd1 _13806_/D sky130_fd_sc_hd__o21a_1
X_07703_ _07700_/Y _07732_/A _07713_/A vssd1 vssd1 vccd1 vccd1 _07703_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_66_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08683_ _13518_/Q _08683_/A2 _08691_/A2 _13589_/Q vssd1 vssd1 vccd1 vccd1 _08683_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_26_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07634_ _14759_/Q _07629_/A _07633_/Y _08002_/C1 vssd1 vssd1 vccd1 vccd1 _13470_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_81_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07565_ _07567_/B _07564_/X _07644_/A vssd1 vssd1 vccd1 vccd1 _07565_/X sky130_fd_sc_hd__a21bo_1
XFILLER_0_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09304_ _15293_/Q _15261_/Q _15229_/Q _15160_/Q _09481_/S _09553_/A1 vssd1 vssd1
+ vccd1 vccd1 _09304_/X sky130_fd_sc_hd__mux4_1
XFILLER_94_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07496_ _14764_/Q _07495_/X _07500_/S vssd1 vssd1 vccd1 vccd1 _07496_/X sky130_fd_sc_hd__mux2_8
XFILLER_167_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09235_ _09419_/A2 _09233_/X _09234_/X _09421_/A1 vssd1 vssd1 vccd1 vccd1 _09235_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_142_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09166_ _13952_/Q _13694_/Q _09441_/S vssd1 vssd1 vccd1 vccd1 _09166_/X sky130_fd_sc_hd__mux2_1
XFILLER_119_34 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08117_ input30/X input7/X input16/X input25/X _08150_/S _08151_/S vssd1 vssd1 vccd1
+ vccd1 _08117_/X sky130_fd_sc_hd__mux4_2
X_09097_ _13916_/Q _09096_/X _12481_/A vssd1 vssd1 vccd1 vccd1 _13916_/D sky130_fd_sc_hd__mux2_1
XFILLER_134_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08048_ _14741_/Q _13619_/Q _08072_/S vssd1 vssd1 vccd1 vccd1 _13619_/D sky130_fd_sc_hd__mux2_1
XFILLER_134_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10010_ _13331_/A0 _14368_/Q _10028_/S vssd1 vssd1 vccd1 vccd1 _14368_/D sky130_fd_sc_hd__mux2_1
XFILLER_88_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09999_ _13320_/A0 _14357_/Q _10029_/S vssd1 vssd1 vccd1 vccd1 _14357_/D sky130_fd_sc_hd__mux2_1
XFILLER_88_275 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11961_ _12582_/A _11961_/B vssd1 vssd1 vccd1 vccd1 _11961_/X sky130_fd_sc_hd__or2_1
XFILLER_57_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10912_ _11436_/B _10944_/B vssd1 vssd1 vccd1 vccd1 _10912_/Y sky130_fd_sc_hd__nand2_1
X_13700_ _15127_/CLK _13700_/D vssd1 vssd1 vccd1 vccd1 _13700_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14680_ _15588_/CLK _14680_/D vssd1 vssd1 vccd1 vccd1 _14680_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_151_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11892_ _12260_/A _11892_/B vssd1 vssd1 vccd1 vccd1 _11892_/X sky130_fd_sc_hd__or2_1
XTAP_3889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13631_ _15389_/CLK _13631_/D vssd1 vssd1 vccd1 vccd1 _13631_/Q sky130_fd_sc_hd__dfxtp_1
X_10843_ _14875_/Q _13793_/Q _12917_/S vssd1 vssd1 vccd1 vccd1 _14875_/D sky130_fd_sc_hd__mux2_1
XFILLER_44_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13562_ _13632_/CLK _13562_/D vssd1 vssd1 vccd1 vccd1 _13562_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10774_ hold7/A _15438_/Q _12910_/S vssd1 vssd1 vccd1 vccd1 _14806_/D sky130_fd_sc_hd__mux2_1
XFILLER_44_96 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15301_ _15301_/CLK _15301_/D vssd1 vssd1 vccd1 vccd1 _15301_/Q sky130_fd_sc_hd__dfxtp_1
X_12513_ _12617_/S _12513_/B vssd1 vssd1 vccd1 vccd1 _12513_/X sky130_fd_sc_hd__or2_1
XFILLER_157_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13493_ _15385_/CLK _13493_/D vssd1 vssd1 vccd1 vccd1 _13493_/Q sky130_fd_sc_hd__dfxtp_2
Xclkbuf_leaf_160_clk clkbuf_5_19_0_clk/X vssd1 vssd1 vccd1 vccd1 _14197_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_100_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12444_ _12582_/A _12444_/B vssd1 vssd1 vccd1 vccd1 _12444_/X sky130_fd_sc_hd__or2_1
X_15232_ _15336_/CLK _15232_/D vssd1 vssd1 vccd1 vccd1 _15232_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_173_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15163_ _15336_/CLK _15163_/D vssd1 vssd1 vccd1 vccd1 _15163_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_125_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12375_ _12617_/S _12375_/B vssd1 vssd1 vccd1 vccd1 _12375_/X sky130_fd_sc_hd__or2_1
XFILLER_181_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14114_ _15315_/CLK _14114_/D vssd1 vssd1 vccd1 vccd1 _14114_/Q sky130_fd_sc_hd__dfxtp_1
X_11326_ _11048_/Y _11296_/A _11325_/X _11307_/A _11323_/Y vssd1 vssd1 vccd1 vccd1
+ _11327_/B sky130_fd_sc_hd__o221a_1
XFILLER_158_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15094_ _15094_/CLK _15094_/D vssd1 vssd1 vccd1 vccd1 _15094_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_180_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14045_ _15133_/CLK _14045_/D vssd1 vssd1 vccd1 vccd1 _14045_/Q sky130_fd_sc_hd__dfxtp_1
X_11257_ _15028_/Q _11302_/A _11255_/X _11256_/X vssd1 vssd1 vccd1 vccd1 _15028_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_80_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10208_ input2/X hold4/A _13284_/S vssd1 vssd1 vccd1 vccd1 _14593_/D sky130_fd_sc_hd__mux2_1
XFILLER_67_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_5_12_0_clk clkbuf_4_6_0_clk/X vssd1 vssd1 vccd1 vccd1 clkbuf_5_12_0_clk/X
+ sky130_fd_sc_hd__clkbuf_8
X_11188_ _14986_/Q _11164_/S _11170_/X _11187_/Y vssd1 vssd1 vccd1 vccd1 _14986_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_94_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10139_ _14524_/Q _13325_/A0 _10159_/S vssd1 vssd1 vccd1 vccd1 _14524_/D sky130_fd_sc_hd__mux2_1
XFILLER_39_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14947_ _15570_/CLK _14947_/D vssd1 vssd1 vccd1 vccd1 _14947_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_5_27_0_clk clkbuf_5_27_0_clk/A vssd1 vssd1 vccd1 vccd1 _15447_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_78_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_120 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14878_ _15592_/CLK _14878_/D vssd1 vssd1 vccd1 vccd1 _14878_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_78_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13829_ _15291_/CLK _13829_/D vssd1 vssd1 vccd1 vccd1 _13829_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07350_ _07350_/A _07350_/B _07350_/C _07350_/D vssd1 vssd1 vccd1 vccd1 _07350_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_188_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07281_ _15320_/Q _15476_/Q _07340_/S vssd1 vssd1 vccd1 vccd1 _07281_/X sky130_fd_sc_hd__mux2_8
XFILLER_176_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_151_clk clkbuf_5_24_0_clk/X vssd1 vssd1 vccd1 vccd1 _15619_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_15_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09020_ _14234_/Q _14266_/Q _14298_/Q _14330_/Q _09073_/S _09234_/S1 vssd1 vssd1
+ vccd1 vccd1 _09020_/X sky130_fd_sc_hd__mux4_1
XFILLER_176_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_1027 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09922_ _13098_/B2 _14283_/Q _09930_/S vssd1 vssd1 vccd1 vccd1 _14283_/D sky130_fd_sc_hd__mux2_1
X_09853_ _14217_/Q _11873_/A1 _09863_/S vssd1 vssd1 vccd1 vccd1 _14217_/D sky130_fd_sc_hd__mux2_1
XFILLER_131_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08804_ _11838_/A1 _13830_/Q _08816_/S vssd1 vssd1 vccd1 vccd1 _13830_/D sky130_fd_sc_hd__mux2_1
XFILLER_86_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09784_ _14151_/Q _11872_/A1 _09795_/S vssd1 vssd1 vccd1 vccd1 _14151_/D sky130_fd_sc_hd__mux2_1
XTAP_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_640 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06996_ _15540_/Q _15615_/Q _12904_/S vssd1 vssd1 vccd1 vccd1 _06997_/C sky130_fd_sc_hd__mux2_1
XTAP_3108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08735_ _13447_/Q _08746_/A2 _08749_/A2 _13582_/Q _08734_/X vssd1 vssd1 vccd1 vccd1
+ _08735_/X sky130_fd_sc_hd__a221o_1
XFILLER_39_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_108 _15344_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08666_ _13794_/Q _08665_/X _12917_/S vssd1 vssd1 vccd1 vccd1 _13794_/D sky130_fd_sc_hd__mux2_1
XFILLER_38_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_119 _07137_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07617_ _13466_/Q _13465_/Q _07617_/C vssd1 vssd1 vccd1 vccd1 _07621_/B sky130_fd_sc_hd__nand3_2
XFILLER_54_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08597_ _14508_/Q _08748_/B1 _08595_/X _08596_/X vssd1 vssd1 vccd1 vccd1 _08598_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_42_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07548_ _13448_/Q _13447_/Q _13446_/Q _13445_/Q vssd1 vssd1 vccd1 vccd1 _07559_/D
+ sky130_fd_sc_hd__and4_2
XFILLER_22_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07479_ _13675_/Q _07483_/A2 _07483_/B1 _14703_/Q _07478_/X vssd1 vssd1 vccd1 vccd1
+ _07479_/X sky130_fd_sc_hd__a221o_1
Xclkbuf_leaf_142_clk clkbuf_5_28_0_clk/X vssd1 vssd1 vccd1 vccd1 _15372_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_167_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09218_ _09202_/X _09205_/X _09212_/X _09217_/X vssd1 vssd1 vccd1 vccd1 _09218_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_10_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10490_ _11561_/A _11563_/A vssd1 vssd1 vccd1 vccd1 _13223_/B sky130_fd_sc_hd__nand2_1
XFILLER_148_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09149_ _09406_/S1 _09147_/X _09148_/X vssd1 vssd1 vccd1 vccd1 _09149_/X sky130_fd_sc_hd__a21o_1
XFILLER_108_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12160_ _15317_/Q _13081_/A2 _12159_/X vssd1 vssd1 vccd1 vccd1 _15317_/D sky130_fd_sc_hd__a21o_1
XFILLER_135_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11111_ _14967_/Q _10984_/Y _11109_/Y _11110_/Y vssd1 vssd1 vccd1 vccd1 _14967_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_122_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12091_ _15314_/Q _13119_/S _12090_/X vssd1 vssd1 vccd1 vccd1 _15314_/D sky130_fd_sc_hd__a21o_1
XFILLER_150_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_967 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11042_ _11356_/C _13159_/B _08273_/A _11356_/B vssd1 vssd1 vccd1 vccd1 _11042_/Y
+ sky130_fd_sc_hd__a211oi_1
XFILLER_77_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14801_ _15619_/CLK _14801_/D vssd1 vssd1 vccd1 vccd1 _14801_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_188_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12993_ _10659_/X _14878_/Q _13029_/S vssd1 vssd1 vccd1 vccd1 _12993_/X sky130_fd_sc_hd__mux2_8
XTAP_3642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_194 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14732_ _15615_/CLK _14732_/D vssd1 vssd1 vccd1 vccd1 _14732_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_3664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11944_ _12615_/A1 _11943_/X _12594_/S vssd1 vssd1 vccd1 vccd1 _11944_/X sky130_fd_sc_hd__a21o_1
XFILLER_44_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14663_ _15634_/CLK _14663_/D vssd1 vssd1 vccd1 vccd1 _14663_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11875_ _15296_/Q _13342_/A0 _11883_/S vssd1 vssd1 vccd1 vccd1 _15296_/D sky130_fd_sc_hd__mux2_1
XTAP_2974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10826_ _14858_/Q _07202_/X _10868_/S vssd1 vssd1 vccd1 vccd1 _14858_/D sky130_fd_sc_hd__mux2_1
X_13614_ _15543_/CLK _13614_/D vssd1 vssd1 vccd1 vccd1 _13614_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14594_ _15620_/CLK _14594_/D vssd1 vssd1 vccd1 vccd1 hold8/A sky130_fd_sc_hd__dfxtp_2
XFILLER_111_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10757_ _15421_/Q _14789_/Q _10759_/S vssd1 vssd1 vccd1 vccd1 _14789_/D sky130_fd_sc_hd__mux2_1
XFILLER_13_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13545_ _15399_/CLK _13545_/D vssd1 vssd1 vccd1 vccd1 _13545_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_133_clk clkbuf_5_29_0_clk/X vssd1 vssd1 vccd1 vccd1 _15398_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_125_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13476_ _14517_/CLK _13476_/D vssd1 vssd1 vccd1 vccd1 _13476_/Q sky130_fd_sc_hd__dfxtp_2
X_10688_ _14984_/Q _10718_/A2 _10722_/B1 _14952_/Q _10687_/X vssd1 vssd1 vccd1 vccd1
+ _10688_/X sky130_fd_sc_hd__a221o_1
XFILLER_9_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15215_ _15279_/CLK _15215_/D vssd1 vssd1 vccd1 vccd1 _15215_/Q sky130_fd_sc_hd__dfxtp_1
X_12427_ _12615_/A1 _12426_/X _12559_/A vssd1 vssd1 vccd1 vccd1 _12427_/X sky130_fd_sc_hd__a21o_1
XFILLER_173_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12358_ _12592_/A1 _12357_/X _12536_/A vssd1 vssd1 vccd1 vccd1 _12358_/X sky130_fd_sc_hd__a21o_1
X_15146_ _15279_/CLK _15146_/D vssd1 vssd1 vccd1 vccd1 _15146_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_486 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11309_ _11309_/A _11309_/B vssd1 vssd1 vccd1 vccd1 _11309_/Y sky130_fd_sc_hd__nand2_1
XFILLER_99_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15077_ _15077_/CLK _15077_/D vssd1 vssd1 vccd1 vccd1 _15077_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12289_ _12592_/A1 _12288_/X _12536_/A vssd1 vssd1 vccd1 vccd1 _12289_/X sky130_fd_sc_hd__a21o_1
XFILLER_84_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14028_ _14405_/CLK _14028_/D vssd1 vssd1 vccd1 vccd1 _14028_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_1071 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_1074 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06850_ _15615_/Q _06830_/X _08390_/B _06833_/X _06849_/X vssd1 vssd1 vccd1 vccd1
+ _06851_/B sky130_fd_sc_hd__a41o_1
XFILLER_132_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06781_ _06782_/A _10735_/S _06782_/C vssd1 vssd1 vccd1 vccd1 _06781_/X sky130_fd_sc_hd__and3_4
XFILLER_82_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08520_ _08668_/C _08520_/B vssd1 vssd1 vccd1 vccd1 _08529_/B sky130_fd_sc_hd__nand2_4
X_08451_ _08451_/A _08773_/B vssd1 vssd1 vccd1 vccd1 _08451_/X sky130_fd_sc_hd__and2_1
XFILLER_24_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07402_ _14652_/Q _07498_/B _07498_/C vssd1 vssd1 vccd1 vccd1 _07402_/X sky130_fd_sc_hd__and3_1
XFILLER_168_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08382_ _11025_/A _13199_/B vssd1 vssd1 vccd1 vccd1 _11036_/B sky130_fd_sc_hd__nor2_1
XFILLER_91_1042 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07333_ _07331_/Y _07332_/X _07327_/A _07329_/Y vssd1 vssd1 vccd1 vccd1 _07333_/X
+ sky130_fd_sc_hd__o2bb2a_1
Xclkbuf_leaf_124_clk clkbuf_5_31_0_clk/X vssd1 vssd1 vccd1 vccd1 _15386_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_52_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07264_ _07264_/A _07264_/B vssd1 vssd1 vccd1 vccd1 _07264_/X sky130_fd_sc_hd__or2_1
XFILLER_137_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09003_ _13880_/Q _09522_/A2 _09519_/B1 _14395_/Q _08507_/A vssd1 vssd1 vccd1 vccd1
+ _09003_/X sky130_fd_sc_hd__a221o_1
X_07195_ _07197_/A vssd1 vssd1 vccd1 vccd1 _07195_/Y sky130_fd_sc_hd__inv_2
XFILLER_132_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout501 _14767_/Q vssd1 vssd1 vccd1 vccd1 _08240_/A sky130_fd_sc_hd__buf_12
X_09905_ _11858_/A1 _14266_/Q _09925_/S vssd1 vssd1 vccd1 vccd1 _14266_/D sky130_fd_sc_hd__mux2_1
Xfanout512 _14607_/Q vssd1 vssd1 vccd1 vccd1 _13049_/A1 sky130_fd_sc_hd__buf_12
Xfanout523 _09466_/A vssd1 vssd1 vccd1 vccd1 _09543_/A sky130_fd_sc_hd__buf_12
Xfanout534 _09511_/S1 vssd1 vssd1 vccd1 vccd1 _09523_/A1 sky130_fd_sc_hd__buf_12
XFILLER_59_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_990 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout545 _09425_/S vssd1 vssd1 vccd1 vccd1 _09132_/S sky130_fd_sc_hd__buf_8
Xfanout556 _08490_/A1 vssd1 vssd1 vccd1 vccd1 _09005_/S sky130_fd_sc_hd__buf_6
X_09836_ _14200_/Q _13323_/A0 _09858_/S vssd1 vssd1 vccd1 vccd1 _14200_/D sky130_fd_sc_hd__mux2_1
XFILLER_58_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout567 _12515_/C1 vssd1 vssd1 vccd1 vccd1 _08449_/A sky130_fd_sc_hd__buf_12
XTAP_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout578 _14600_/Q vssd1 vssd1 vccd1 vccd1 _08453_/A sky130_fd_sc_hd__buf_12
XTAP_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout589 _14599_/Q vssd1 vssd1 vccd1 vccd1 _12061_/A sky130_fd_sc_hd__buf_12
XFILLER_74_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06979_ _06971_/X _06978_/Y _06975_/Y _06974_/B vssd1 vssd1 vccd1 vccd1 _06979_/X
+ sky130_fd_sc_hd__a211o_1
X_09767_ _14134_/Q _11680_/A0 _09790_/S vssd1 vssd1 vccd1 vccd1 _14134_/D sky130_fd_sc_hd__mux2_1
XFILLER_86_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08718_ _13449_/Q _08746_/A2 _08749_/A2 _13584_/Q _08717_/X vssd1 vssd1 vccd1 vccd1
+ _08722_/B sky130_fd_sc_hd__a221o_1
XFILLER_132_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09698_ _11853_/A1 _14068_/Q _09728_/S vssd1 vssd1 vccd1 vccd1 _14068_/D sky130_fd_sc_hd__mux2_1
XFILLER_92_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08649_ _15382_/Q _08690_/A2 _08690_/B1 _13427_/Q vssd1 vssd1 vccd1 vccd1 _08649_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_1514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_1076 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11660_ _13335_/A0 _15092_/Q _11670_/S vssd1 vssd1 vccd1 vccd1 _15092_/D sky130_fd_sc_hd__mux2_1
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_668 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10611_ _15001_/Q _10569_/B _10733_/A2 _14969_/Q _10732_/C1 vssd1 vssd1 vccd1 vccd1
+ _10611_/X sky130_fd_sc_hd__a221o_1
XFILLER_186_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_115_clk _15447_/CLK vssd1 vssd1 vccd1 vccd1 _15636_/CLK sky130_fd_sc_hd__clkbuf_16
X_11591_ _11598_/A _11591_/B vssd1 vssd1 vccd1 vccd1 _11593_/B sky130_fd_sc_hd__xnor2_1
XFILLER_168_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13330_ _13330_/A0 _15660_/Q _13345_/S vssd1 vssd1 vccd1 vccd1 _15660_/D sky130_fd_sc_hd__mux2_1
XFILLER_167_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10542_ _10542_/A _10542_/B vssd1 vssd1 vccd1 vccd1 _10543_/C sky130_fd_sc_hd__nand2_1
XFILLER_127_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13261_ _15345_/Q _15592_/Q _13288_/S vssd1 vssd1 vccd1 vccd1 _15592_/D sky130_fd_sc_hd__mux2_1
X_10473_ _07233_/A _10360_/B _10472_/X vssd1 vssd1 vccd1 vccd1 _11589_/B sky130_fd_sc_hd__a21oi_4
X_12212_ _14370_/Q _15186_/Q _13825_/Q _14564_/Q _12489_/S0 _12489_/S1 vssd1 vssd1
+ vccd1 vccd1 _12212_/X sky130_fd_sc_hd__mux4_1
X_15000_ _15000_/CLK _15000_/D vssd1 vssd1 vccd1 vccd1 _15000_/Q sky130_fd_sc_hd__dfxtp_1
X_13192_ _06769_/Y _11457_/A _13214_/B vssd1 vssd1 vccd1 vccd1 _13192_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_68_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12143_ _14367_/Q _15183_/Q _13822_/Q _14561_/Q _12154_/S _12253_/S1 vssd1 vssd1
+ vccd1 vccd1 _12143_/X sky130_fd_sc_hd__mux4_1
XFILLER_124_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12074_ _14364_/Q _15180_/Q _13819_/Q _14558_/Q _12079_/S _12080_/A vssd1 vssd1 vccd1
+ vccd1 _12074_/X sky130_fd_sc_hd__mux4_1
XFILLER_150_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11025_ _11025_/A _13220_/B vssd1 vssd1 vccd1 vccd1 _11027_/A sky130_fd_sc_hd__nand2_1
XFILLER_77_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12976_ _13072_/B2 _13024_/A2 _12975_/X _13024_/B2 vssd1 vssd1 vccd1 vccd1 _12976_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_3472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14715_ _15525_/CLK _14715_/D vssd1 vssd1 vccd1 vccd1 _14715_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_3494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11927_ _11910_/X _11911_/X _12617_/S vssd1 vssd1 vccd1 vccd1 _11927_/X sky130_fd_sc_hd__mux2_1
XTAP_2760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14646_ _15534_/CLK _14646_/D vssd1 vssd1 vccd1 vccd1 _14646_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11858_ _15279_/Q _11858_/A1 _11878_/S vssd1 vssd1 vccd1 vccd1 _15279_/D sky130_fd_sc_hd__mux2_1
XFILLER_82_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_106_clk clkbuf_5_26_0_clk/X vssd1 vssd1 vccd1 vccd1 _15643_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_158_320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10809_ _14841_/Q _07297_/A _12481_/A vssd1 vssd1 vccd1 vccd1 _14841_/D sky130_fd_sc_hd__mux2_1
XANTENNA_19 _15046_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11789_ _15212_/Q _13322_/A0 _11816_/S vssd1 vssd1 vccd1 vccd1 _15212_/D sky130_fd_sc_hd__mux2_1
X_14577_ _15542_/CLK _14577_/D vssd1 vssd1 vccd1 vccd1 _14577_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_174_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13528_ _13632_/CLK _13528_/D vssd1 vssd1 vccd1 vccd1 _13528_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_9_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13459_ _15381_/CLK _13459_/D vssd1 vssd1 vccd1 vccd1 _13459_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_63_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15129_ _15544_/CLK _15129_/D vssd1 vssd1 vccd1 vccd1 _15129_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_142_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07951_ _07964_/A _07951_/B vssd1 vssd1 vccd1 vccd1 _07951_/Y sky130_fd_sc_hd__nand2_1
XFILLER_114_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06902_ _15376_/Q _07571_/B _15375_/Q _06739_/Y _06901_/X vssd1 vssd1 vccd1 vccd1
+ _06902_/X sky130_fd_sc_hd__a221o_1
X_07882_ _07903_/A _07882_/B vssd1 vssd1 vccd1 vccd1 _07882_/Y sky130_fd_sc_hd__nand2_1
XFILLER_96_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09621_ _13995_/Q _11876_/A1 _09627_/S vssd1 vssd1 vccd1 vccd1 _13995_/D sky130_fd_sc_hd__mux2_1
XFILLER_83_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06833_ _14596_/Q hold5/A _14592_/Q _08770_/C vssd1 vssd1 vccd1 vccd1 _06833_/X sky130_fd_sc_hd__or4_1
XFILLER_56_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09552_ _14098_/Q _08494_/Y _08512_/B _14066_/Q _09543_/A vssd1 vssd1 vccd1 vccd1
+ _09552_/X sky130_fd_sc_hd__a221o_1
X_06764_ input22/X vssd1 vssd1 vccd1 vccd1 _06764_/Y sky130_fd_sc_hd__inv_2
X_08503_ _08538_/A _08513_/A vssd1 vssd1 vccd1 vccd1 _08503_/Y sky130_fd_sc_hd__nor2_4
XFILLER_102_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09483_ _09553_/A1 _09481_/X _09482_/X vssd1 vssd1 vccd1 vccd1 _09487_/B sky130_fd_sc_hd__a21o_1
XFILLER_93_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06695_ _13505_/Q vssd1 vssd1 vccd1 vccd1 _06873_/B sky130_fd_sc_hd__inv_2
XFILLER_36_495 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08434_ _13747_/Q _12906_/S _08426_/B _08433_/X vssd1 vssd1 vccd1 vccd1 _13747_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_52_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08365_ _11034_/B _11036_/A vssd1 vssd1 vccd1 vccd1 _08366_/A sky130_fd_sc_hd__nor2_1
XFILLER_32_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07316_ _15313_/Q _15469_/Q _07340_/S vssd1 vssd1 vccd1 vccd1 _07317_/A sky130_fd_sc_hd__mux2_4
XFILLER_177_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08296_ _11356_/C _11399_/A _10999_/B _11356_/B vssd1 vssd1 vccd1 vccd1 _08296_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_178_1003 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07247_ _15324_/Q _15480_/Q _07335_/S vssd1 vssd1 vccd1 vccd1 _07248_/A sky130_fd_sc_hd__mux2_8
XFILLER_178_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_4_2_0_clk clkbuf_4_3_0_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_5_5_0_clk/A sky130_fd_sc_hd__clkbuf_8
XFILLER_178_1058 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07178_ _15352_/Q _15059_/Q _07188_/S vssd1 vssd1 vccd1 vccd1 _07178_/X sky130_fd_sc_hd__mux2_8
XFILLER_3_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout320 _07432_/X vssd1 vssd1 vccd1 vccd1 _13080_/B2 sky130_fd_sc_hd__buf_8
Xfanout331 _07408_/X vssd1 vssd1 vccd1 vccd1 _13327_/A0 sky130_fd_sc_hd__buf_6
Xfanout342 _13322_/A0 vssd1 vssd1 vccd1 vccd1 _11680_/A0 sky130_fd_sc_hd__buf_6
XFILLER_87_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout353 _10581_/X vssd1 vssd1 vccd1 vccd1 _10602_/B sky130_fd_sc_hd__buf_12
Xfanout364 _08508_/Y vssd1 vssd1 vccd1 vccd1 _09522_/B1 sky130_fd_sc_hd__buf_12
XFILLER_59_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout375 _11023_/A vssd1 vssd1 vccd1 vccd1 _11025_/A sky130_fd_sc_hd__buf_6
XFILLER_86_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout386 _11047_/B vssd1 vssd1 vccd1 vccd1 _11297_/S sky130_fd_sc_hd__buf_12
Xfanout397 _11129_/A vssd1 vssd1 vccd1 vccd1 _11329_/A sky130_fd_sc_hd__clkbuf_4
X_09819_ _14185_/Q _13341_/A0 _09828_/S vssd1 vssd1 vccd1 vccd1 _14185_/D sky130_fd_sc_hd__mux2_1
XFILLER_59_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12830_ _13443_/Q _12647_/B _08030_/Y _13610_/Q _12743_/A vssd1 vssd1 vccd1 vccd1
+ _12830_/X sky130_fd_sc_hd__a221o_1
XTAP_2012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12761_ _15357_/Q _12767_/C vssd1 vssd1 vccd1 vccd1 _12761_/X sky130_fd_sc_hd__xor2_1
XFILLER_43_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14500_ _15383_/CLK _14500_/D vssd1 vssd1 vccd1 vccd1 _14500_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11712_ _15141_/Q _13320_/A0 _11742_/S vssd1 vssd1 vccd1 vccd1 _15141_/D sky130_fd_sc_hd__mux2_1
XTAP_2089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12692_ _13424_/Q _12691_/X _12728_/S vssd1 vssd1 vccd1 vccd1 _12693_/B sky130_fd_sc_hd__mux2_1
XTAP_1355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15480_ _15489_/CLK _15480_/D vssd1 vssd1 vccd1 vccd1 _15480_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_43_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14431_ _15663_/CLK _14431_/D vssd1 vssd1 vccd1 vccd1 _14431_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11643_ _14714_/Q _14715_/Q _13318_/C _11818_/A vssd1 vssd1 vccd1 vccd1 _11643_/X
+ sky130_fd_sc_hd__or4_4
XFILLER_14_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11574_ _11564_/A _11566_/X _11576_/D _11614_/S vssd1 vssd1 vccd1 vccd1 _11574_/X
+ sky130_fd_sc_hd__a31o_1
X_14362_ _15178_/CLK _14362_/D vssd1 vssd1 vccd1 vccd1 _14362_/Q sky130_fd_sc_hd__dfxtp_1
Xinput17 ext_read_data[24] vssd1 vssd1 vccd1 vccd1 input17/X sky130_fd_sc_hd__buf_6
XFILLER_168_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_1095 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput28 ext_read_data[5] vssd1 vssd1 vccd1 vccd1 input28/X sky130_fd_sc_hd__buf_6
XFILLER_122_1046 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_96 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10525_ _13215_/B _13214_/A vssd1 vssd1 vccd1 vccd1 _10526_/B sky130_fd_sc_hd__nand2b_1
XFILLER_10_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13313_ _15644_/Q _12813_/B _13316_/S vssd1 vssd1 vccd1 vccd1 _15644_/D sky130_fd_sc_hd__mux2_1
X_14293_ _14606_/CLK _14293_/D vssd1 vssd1 vccd1 vccd1 _14293_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_156_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13244_ _13242_/Y _13243_/X _15581_/Q _13252_/B vssd1 vssd1 vccd1 vccd1 _15581_/D
+ sky130_fd_sc_hd__a2bb2o_1
X_10456_ _10520_/A1 _13779_/Q _13747_/Q _10520_/B2 vssd1 vssd1 vccd1 vccd1 _10456_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_108_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13175_ _13242_/A _11399_/A _13219_/S vssd1 vssd1 vccd1 vccd1 _13175_/X sky130_fd_sc_hd__o21a_1
X_10387_ _11440_/A _11476_/B vssd1 vssd1 vccd1 vccd1 _10387_/X sky130_fd_sc_hd__and2_1
X_12126_ _12498_/A _12126_/B vssd1 vssd1 vccd1 vccd1 _12126_/X sky130_fd_sc_hd__and2_1
XFILLER_69_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12057_ _12452_/A _12057_/B vssd1 vssd1 vccd1 vccd1 _12057_/X sky130_fd_sc_hd__and2_1
X_11008_ _11023_/A _13233_/B vssd1 vssd1 vccd1 vccd1 _11312_/A sky130_fd_sc_hd__nand2_1
XFILLER_81_1096 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_398 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12959_ _15466_/Q _13081_/A2 _13025_/B1 _12958_/X vssd1 vssd1 vccd1 vccd1 _15466_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_45_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15678_ _15678_/CLK _15678_/D vssd1 vssd1 vccd1 vccd1 _15678_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14629_ _15596_/CLK _14629_/D vssd1 vssd1 vccd1 vccd1 _14629_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_159_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08150_ input7/X input16/X _08150_/S vssd1 vssd1 vccd1 vccd1 _08150_/X sky130_fd_sc_hd__mux2_1
XFILLER_20_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07101_ _07115_/B _07163_/A vssd1 vssd1 vccd1 vccd1 _07101_/X sky130_fd_sc_hd__and2_4
XFILLER_174_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08081_ _06825_/C _08080_/X _12640_/S vssd1 vssd1 vccd1 vccd1 _08081_/X sky130_fd_sc_hd__a21o_1
XFILLER_173_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07032_ _07031_/X _14743_/Q _07077_/S vssd1 vssd1 vccd1 vccd1 _13589_/D sky130_fd_sc_hd__mux2_1
XFILLER_146_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08983_ _14071_/Q _09231_/A2 _09403_/B1 _14039_/Q _09221_/A vssd1 vssd1 vccd1 vccd1
+ _08983_/X sky130_fd_sc_hd__a221o_1
XFILLER_88_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07934_ _14741_/Q _08012_/A2 _07933_/Y vssd1 vssd1 vccd1 vccd1 _13548_/D sky130_fd_sc_hd__o21a_1
XFILLER_102_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07865_ _14755_/Q _07874_/A _07864_/X _08002_/C1 vssd1 vssd1 vccd1 vccd1 _13530_/D
+ sky130_fd_sc_hd__o211a_1
X_09604_ _13978_/Q _13326_/A0 _09627_/S vssd1 vssd1 vccd1 vccd1 _13978_/D sky130_fd_sc_hd__mux2_1
X_06816_ _13733_/Q _13730_/Q _13731_/Q _13729_/Q vssd1 vssd1 vccd1 vccd1 _06817_/B
+ sky130_fd_sc_hd__or4_1
X_07796_ _07798_/B _07795_/Y _07816_/A vssd1 vssd1 vccd1 vccd1 _07796_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_71_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09535_ _13873_/Q _14226_/Q _09535_/S vssd1 vssd1 vccd1 vccd1 _09535_/X sky130_fd_sc_hd__mux2_1
X_06747_ _13449_/Q vssd1 vssd1 vccd1 vccd1 _06747_/Y sky130_fd_sc_hd__inv_2
XFILLER_25_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09466_ _09466_/A _09466_/B vssd1 vssd1 vccd1 vccd1 _09466_/X sky130_fd_sc_hd__or2_1
XFILLER_184_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1027 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06678_ _14905_/Q vssd1 vssd1 vccd1 vccd1 _06678_/Y sky130_fd_sc_hd__inv_2
XFILLER_40_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08417_ _14596_/Q _08390_/A _06991_/B _08477_/C vssd1 vssd1 vccd1 vccd1 _08417_/X
+ sky130_fd_sc_hd__a211o_1
X_09397_ _14478_/Q _09536_/A2 _13130_/B1 _14446_/Q _09396_/X vssd1 vssd1 vccd1 vccd1
+ _09397_/X sky130_fd_sc_hd__a221o_1
XFILLER_185_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08348_ _08307_/B _08381_/B _11047_/B vssd1 vssd1 vccd1 vccd1 _08348_/X sky130_fd_sc_hd__mux2_1
XFILLER_164_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08279_ _11349_/B _11383_/A vssd1 vssd1 vccd1 vccd1 _10999_/A sky130_fd_sc_hd__nor2_1
X_10310_ _14695_/Q _14880_/Q _10715_/S vssd1 vssd1 vccd1 vccd1 _14695_/D sky130_fd_sc_hd__mux2_1
XFILLER_152_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11290_ _11329_/A _11290_/B vssd1 vssd1 vccd1 vccd1 _11290_/Y sky130_fd_sc_hd__nor2_1
XFILLER_138_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10241_ _14626_/Q _14779_/Q _10650_/S vssd1 vssd1 vccd1 vccd1 _14626_/D sky130_fd_sc_hd__mux2_1
XFILLER_98_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10172_ _11858_/A1 _14556_/Q _10192_/S vssd1 vssd1 vccd1 vccd1 _14556_/D sky130_fd_sc_hd__mux2_1
XFILLER_79_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14980_ _14988_/CLK _14980_/D vssd1 vssd1 vccd1 vccd1 _14980_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout150 _12910_/S vssd1 vssd1 vccd1 vccd1 _12878_/S sky130_fd_sc_hd__buf_8
Xfanout161 _08626_/S vssd1 vssd1 vccd1 vccd1 _12928_/S sky130_fd_sc_hd__buf_8
Xfanout172 _11785_/Y vssd1 vssd1 vccd1 vccd1 _11817_/S sky130_fd_sc_hd__buf_12
XFILLER_87_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13931_ _15518_/CLK _13931_/D vssd1 vssd1 vccd1 vccd1 _13931_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout183 _10099_/X vssd1 vssd1 vccd1 vccd1 _10131_/S sky130_fd_sc_hd__buf_12
Xfanout194 _09931_/Y vssd1 vssd1 vccd1 vccd1 _09963_/S sky130_fd_sc_hd__buf_12
XFILLER_93_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13862_ _15275_/CLK _13862_/D vssd1 vssd1 vccd1 vccd1 _13862_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_74_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15601_ _15635_/CLK _15601_/D vssd1 vssd1 vccd1 vccd1 _15601_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12813_ _12828_/A _12813_/B vssd1 vssd1 vccd1 vccd1 _12813_/X sky130_fd_sc_hd__or2_1
X_13793_ _15596_/CLK _13793_/D vssd1 vssd1 vccd1 vccd1 _13793_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_27_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_40 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15532_ _15648_/CLK _15532_/D vssd1 vssd1 vccd1 vccd1 _15532_/Q sky130_fd_sc_hd__dfxtp_1
X_12744_ _15354_/Q _12759_/B _12743_/X _12788_/C1 vssd1 vssd1 vccd1 vccd1 _15354_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_37_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15463_ _15499_/CLK _15463_/D vssd1 vssd1 vccd1 vccd1 _15463_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_188_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12675_ _13589_/Q _12674_/X _12785_/B vssd1 vssd1 vccd1 vccd1 _12675_/X sky130_fd_sc_hd__mux2_1
XTAP_1196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14414_ _15673_/CLK _14414_/D vssd1 vssd1 vccd1 vccd1 _14414_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_169_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11626_ _11626_/A _11626_/B vssd1 vssd1 vccd1 vccd1 _11627_/B sky130_fd_sc_hd__nand2_1
X_15394_ _15397_/CLK _15394_/D vssd1 vssd1 vccd1 vccd1 _15394_/Q sky130_fd_sc_hd__dfxtp_1
X_14345_ _15544_/CLK _14345_/D vssd1 vssd1 vccd1 vccd1 _14345_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_183_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11557_ _11542_/A _11548_/Y _11576_/B vssd1 vssd1 vccd1 vccd1 _11557_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_156_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10508_ _07241_/A _10523_/A2 _10507_/X vssd1 vssd1 vccd1 vccd1 _13217_/B sky130_fd_sc_hd__a21oi_4
X_11488_ _13233_/A _11496_/A _10362_/X _11478_/B vssd1 vssd1 vccd1 vccd1 _11491_/C
+ sky130_fd_sc_hd__o211ai_2
XFILLER_6_163 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14276_ _15289_/CLK _14276_/D vssd1 vssd1 vccd1 vccd1 _14276_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_137_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10439_ _07201_/A _10481_/B _10438_/X vssd1 vssd1 vccd1 vccd1 _11626_/A sky130_fd_sc_hd__a21oi_4
X_13227_ _13242_/A _13226_/B _13252_/B _11589_/B vssd1 vssd1 vccd1 vccd1 _13227_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_83_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_170_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13158_ _15553_/Q _13252_/B _13157_/X vssd1 vssd1 vccd1 vccd1 _15553_/D sky130_fd_sc_hd__a21o_1
XTAP_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12109_ _12500_/A1 _12108_/X _12500_/B1 vssd1 vssd1 vccd1 vccd1 _12109_/X sky130_fd_sc_hd__a21o_1
XFILLER_97_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13089_ _15512_/Q _13129_/A _13042_/A _13088_/X vssd1 vssd1 vccd1 vccd1 _15512_/D
+ sky130_fd_sc_hd__a22o_1
XTAP_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07650_ _13475_/Q _07650_/B vssd1 vssd1 vccd1 vccd1 _07651_/B sky130_fd_sc_hd__xnor2_1
XFILLER_65_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07581_ _07579_/Y _07583_/B _07607_/A vssd1 vssd1 vccd1 vccd1 _07581_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_53_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09320_ _15669_/Q _13403_/Q _09481_/S vssd1 vssd1 vccd1 vccd1 _09320_/X sky130_fd_sc_hd__mux2_1
XFILLER_22_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09251_ _09550_/A1 _09249_/X _09250_/X vssd1 vssd1 vccd1 vccd1 _09252_/C sky130_fd_sc_hd__a21o_1
XFILLER_61_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08202_ _13693_/Q _11689_/A0 _08216_/S vssd1 vssd1 vccd1 vccd1 _13693_/D sky130_fd_sc_hd__mux2_1
X_09182_ _15287_/Q _15255_/Q _15223_/Q _15154_/Q _09444_/S _09448_/S1 vssd1 vssd1
+ vccd1 vccd1 _09182_/X sky130_fd_sc_hd__mux4_1
XFILLER_147_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08133_ input3/X input11/X _08133_/S vssd1 vssd1 vccd1 vccd1 _08133_/X sky130_fd_sc_hd__mux2_1
XFILLER_174_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08064_ _14757_/Q _13635_/Q _08066_/S vssd1 vssd1 vccd1 vccd1 _13635_/D sky130_fd_sc_hd__mux2_1
XFILLER_135_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07015_ _14617_/Q _14649_/Q _07096_/S vssd1 vssd1 vccd1 vccd1 _07015_/X sky130_fd_sc_hd__mux2_1
XFILLER_134_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08966_ _15111_/Q _15079_/Q _15652_/Q _13386_/Q _09047_/S _09530_/S1 vssd1 vssd1
+ vccd1 vccd1 _08966_/X sky130_fd_sc_hd__mux4_1
XFILLER_29_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07917_ _13544_/Q _07924_/D vssd1 vssd1 vccd1 vccd1 _07921_/B sky130_fd_sc_hd__nand2_1
XFILLER_112_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08897_ _13875_/Q _09231_/A2 _09403_/B1 _14390_/Q _09445_/C1 vssd1 vssd1 vccd1 vccd1
+ _08897_/X sky130_fd_sc_hd__a221o_1
XFILLER_25_1086 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_95_clk clkbuf_5_24_0_clk/X vssd1 vssd1 vccd1 vccd1 _15622_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_29_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07848_ _13525_/Q _13524_/Q _07847_/D _13526_/Q vssd1 vssd1 vccd1 vccd1 _07848_/Y
+ sky130_fd_sc_hd__a31oi_1
XFILLER_72_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_590 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07779_ _07787_/A _13509_/Q _08817_/B vssd1 vssd1 vccd1 vccd1 _07779_/X sky130_fd_sc_hd__and3_1
XFILLER_72_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_88 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09518_ _13969_/Q _13711_/Q _09521_/S vssd1 vssd1 vccd1 vccd1 _09518_/X sky130_fd_sc_hd__mux2_1
X_10790_ _14822_/Q _15454_/Q _12927_/S vssd1 vssd1 vccd1 vccd1 _14822_/D sky130_fd_sc_hd__mux2_1
XFILLER_140_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09449_ _09449_/A1 _09447_/X _09448_/X _09449_/B2 vssd1 vssd1 vccd1 vccd1 _09449_/X
+ sky130_fd_sc_hd__a22o_1
XPHY_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12460_ _14253_/Q _14285_/Q _14317_/Q _14349_/Q _12489_/S0 _12465_/S1 vssd1 vssd1
+ vccd1 vccd1 _12460_/X sky130_fd_sc_hd__mux4_1
XFILLER_71_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11411_ _11400_/B _11404_/B _11421_/A vssd1 vssd1 vccd1 vccd1 _11412_/B sky130_fd_sc_hd__o21ba_1
XFILLER_138_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12391_ _14250_/Q _14282_/Q _14314_/Q _14346_/Q _12591_/S _12590_/A vssd1 vssd1 vccd1
+ vccd1 _12391_/X sky130_fd_sc_hd__mux4_1
XFILLER_137_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11342_ _11259_/S _11331_/Y _11341_/Y _08249_/Y vssd1 vssd1 vccd1 vccd1 _11344_/B
+ sky130_fd_sc_hd__o211a_1
X_14130_ _15680_/CLK _14130_/D vssd1 vssd1 vccd1 vccd1 _14130_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_181_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11273_ _11258_/Y _11272_/Y _11318_/S vssd1 vssd1 vccd1 vccd1 _11273_/X sky130_fd_sc_hd__mux2_1
XFILLER_4_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14061_ _14093_/CLK _14061_/D vssd1 vssd1 vccd1 vccd1 _14061_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_125_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13012_ _07464_/X _13039_/A2 _13011_/X _12944_/A vssd1 vssd1 vccd1 vccd1 _13012_/X
+ sky130_fd_sc_hd__a22o_1
X_10224_ input19/X _14609_/Q _13291_/S vssd1 vssd1 vccd1 vccd1 _14609_/D sky130_fd_sc_hd__mux2_1
XFILLER_79_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10155_ _14540_/Q _13341_/A0 _10164_/S vssd1 vssd1 vccd1 vccd1 _14540_/D sky130_fd_sc_hd__mux2_1
X_10086_ _14442_/Q _11872_/A1 _10097_/S vssd1 vssd1 vccd1 vccd1 _14442_/D sky130_fd_sc_hd__mux2_1
X_14963_ _14966_/CLK _14963_/D vssd1 vssd1 vccd1 vccd1 _14963_/Q sky130_fd_sc_hd__dfxtp_1
Xhold6 hold6/A vssd1 vssd1 vccd1 vccd1 hold6/X sky130_fd_sc_hd__bufbuf_16
Xclkbuf_leaf_86_clk clkbuf_5_13_0_clk/X vssd1 vssd1 vccd1 vccd1 _14703_/CLK sky130_fd_sc_hd__clkbuf_16
X_13914_ _15501_/CLK _13914_/D vssd1 vssd1 vccd1 vccd1 _13914_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14894_ _15530_/CLK _14894_/D vssd1 vssd1 vccd1 vccd1 _14894_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13845_ _15651_/CLK _13845_/D vssd1 vssd1 vccd1 vccd1 _13845_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13776_ _15398_/CLK _13776_/D vssd1 vssd1 vccd1 vccd1 _13776_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_15_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10988_ _11318_/S _10985_/Y _10987_/X vssd1 vssd1 vccd1 vccd1 _10988_/Y sky130_fd_sc_hd__o21ai_1
X_15515_ _15525_/CLK _15515_/D vssd1 vssd1 vccd1 vccd1 _15515_/Q sky130_fd_sc_hd__dfxtp_1
X_12727_ _13596_/Q _12726_/X _12763_/S vssd1 vssd1 vccd1 vccd1 _12727_/X sky130_fd_sc_hd__mux2_1
X_15446_ _15446_/CLK _15446_/D vssd1 vssd1 vccd1 vccd1 _15446_/Q sky130_fd_sc_hd__dfxtp_1
X_12658_ _15342_/Q _12657_/C _15343_/Q vssd1 vssd1 vccd1 vccd1 _12659_/B sky130_fd_sc_hd__a21oi_1
XFILLER_30_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11609_ _11600_/A _11599_/B _13236_/A vssd1 vssd1 vccd1 vccd1 _11610_/B sky130_fd_sc_hd__a21o_2
X_15377_ _15377_/CLK _15377_/D vssd1 vssd1 vccd1 vccd1 _15377_/Q sky130_fd_sc_hd__dfxtp_1
X_12589_ _14033_/Q _14001_/Q _12591_/S vssd1 vssd1 vccd1 vccd1 _12590_/B sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_10_clk clkbuf_5_2_0_clk/X vssd1 vssd1 vccd1 vccd1 _15674_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_172_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14328_ _15284_/CLK _14328_/D vssd1 vssd1 vccd1 vccd1 _14328_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14259_ _15203_/CLK _14259_/D vssd1 vssd1 vccd1 vccd1 _14259_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_143_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08820_ _13843_/Q _11852_/A1 _08846_/S vssd1 vssd1 vccd1 vccd1 _13843_/D sky130_fd_sc_hd__mux2_1
XTAP_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08751_ _13129_/A _08751_/B _08751_/C vssd1 vssd1 vccd1 vccd1 _08751_/X sky130_fd_sc_hd__or3_4
XTAP_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_77_clk clkbuf_5_15_0_clk/X vssd1 vssd1 vccd1 vccd1 _15626_/CLK sky130_fd_sc_hd__clkbuf_16
X_07702_ _07717_/A _07717_/B vssd1 vssd1 vccd1 vccd1 _07732_/A sky130_fd_sc_hd__and2_2
XFILLER_38_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08682_ _13796_/Q _12927_/S _08681_/X vssd1 vssd1 vccd1 vccd1 _13796_/D sky130_fd_sc_hd__o21a_1
XFILLER_38_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07633_ _07631_/Y _07635_/B _07629_/A vssd1 vssd1 vccd1 vccd1 _07633_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_54_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07564_ _13452_/Q _07576_/C vssd1 vssd1 vccd1 vccd1 _07564_/X sky130_fd_sc_hd__or2_1
XFILLER_53_368 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09303_ _13926_/Q _13149_/S _09302_/X vssd1 vssd1 vccd1 vccd1 _13926_/D sky130_fd_sc_hd__a21o_1
X_07495_ _13679_/Q _07499_/A2 _07499_/B1 _14707_/Q _07494_/X vssd1 vssd1 vccd1 vccd1
+ _07495_/X sky130_fd_sc_hd__a221o_1
XFILLER_55_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09234_ _14534_/Q _14147_/Q _14179_/Q _14115_/Q _09230_/S _09234_/S1 vssd1 vssd1
+ vccd1 vccd1 _09234_/X sky130_fd_sc_hd__mux4_1
X_09165_ _09419_/A2 _09163_/X _09164_/X _09421_/A1 _14607_/Q vssd1 vssd1 vccd1 vccd1
+ _09165_/X sky130_fd_sc_hd__a221o_1
XFILLER_147_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08116_ input16/X input25/X _08133_/S vssd1 vssd1 vccd1 vccd1 _08169_/B sky130_fd_sc_hd__mux2_1
XFILLER_175_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09096_ _06676_/A _09085_/X _09094_/X _09095_/X vssd1 vssd1 vccd1 vccd1 _09096_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_119_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08047_ _14740_/Q _13618_/Q _08072_/S vssd1 vssd1 vccd1 vccd1 _13618_/D sky130_fd_sc_hd__mux2_1
XFILLER_150_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_874 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09998_ _11852_/A1 _14356_/Q _10028_/S vssd1 vssd1 vccd1 vccd1 _14356_/D sky130_fd_sc_hd__mux2_1
XFILLER_95_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08949_ _12573_/A _08949_/B _08949_/C vssd1 vssd1 vccd1 vccd1 _08949_/X sky130_fd_sc_hd__and3_2
Xclkbuf_leaf_68_clk clkbuf_5_14_0_clk/X vssd1 vssd1 vccd1 vccd1 _15572_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_85_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11960_ _15276_/Q _15244_/Q _15212_/Q _15143_/Q _12079_/S _12268_/A vssd1 vssd1 vccd1
+ vccd1 _11961_/B sky130_fd_sc_hd__mux4_1
XFILLER_57_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10911_ _14938_/Q _10944_/B _10910_/Y _08313_/Y vssd1 vssd1 vccd1 vccd1 _14938_/D
+ sky130_fd_sc_hd__o22a_1
XTAP_3868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11891_ _15273_/Q _15241_/Q _15209_/Q _15140_/Q _12154_/S _12253_/S1 vssd1 vssd1
+ vccd1 vccd1 _11892_/B sky130_fd_sc_hd__mux4_1
X_13630_ _15386_/CLK _13630_/D vssd1 vssd1 vccd1 vccd1 _13630_/Q sky130_fd_sc_hd__dfxtp_1
X_10842_ _14874_/Q _13794_/Q _12917_/S vssd1 vssd1 vccd1 vccd1 _14874_/D sky130_fd_sc_hd__mux2_1
XFILLER_53_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13561_ _13632_/CLK _13561_/D vssd1 vssd1 vccd1 vccd1 _13561_/Q sky130_fd_sc_hd__dfxtp_2
X_10773_ _14805_/Q _15437_/Q _12933_/S vssd1 vssd1 vccd1 vccd1 _14805_/D sky130_fd_sc_hd__mux2_1
XFILLER_185_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15300_ _15300_/CLK _15300_/D vssd1 vssd1 vccd1 vccd1 _15300_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12512_ _15300_/Q _15268_/Q _15236_/Q _15167_/Q _12522_/S _12521_/A vssd1 vssd1 vccd1
+ vccd1 _12513_/B sky130_fd_sc_hd__mux4_1
X_13492_ _15389_/CLK _13492_/D vssd1 vssd1 vccd1 vccd1 _13492_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_139_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15231_ _15295_/CLK _15231_/D vssd1 vssd1 vccd1 vccd1 _15231_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12443_ _15297_/Q _15265_/Q _15233_/Q _15164_/Q _12453_/S _12452_/A vssd1 vssd1 vccd1
+ vccd1 _12444_/B sky130_fd_sc_hd__mux4_1
XFILLER_60_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_207 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15162_ _15295_/CLK _15162_/D vssd1 vssd1 vccd1 vccd1 _15162_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12374_ _15294_/Q _15262_/Q _15230_/Q _15161_/Q _12522_/S _12379_/A vssd1 vssd1 vccd1
+ vccd1 _12375_/B sky130_fd_sc_hd__mux4_1
XFILLER_126_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14113_ _15663_/CLK _14113_/D vssd1 vssd1 vccd1 vccd1 _14113_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11325_ _11312_/Y _11324_/Y _11349_/A vssd1 vssd1 vccd1 vccd1 _11325_/X sky130_fd_sc_hd__mux2_2
X_15093_ _15666_/CLK _15093_/D vssd1 vssd1 vccd1 vccd1 _15093_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11256_ _11344_/A _08249_/Y _08259_/Y _11346_/A2 vssd1 vssd1 vccd1 vccd1 _11256_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_140_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14044_ _14415_/CLK _14044_/D vssd1 vssd1 vccd1 vccd1 _14044_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_140_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10207_ input32/X _14592_/Q _13291_/S vssd1 vssd1 vccd1 vccd1 _14592_/D sky130_fd_sc_hd__mux2_1
X_11187_ _11199_/A _11187_/B vssd1 vssd1 vccd1 vccd1 _11187_/Y sky130_fd_sc_hd__nor2_1
XFILLER_121_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10138_ _14523_/Q _11649_/A0 _10164_/S vssd1 vssd1 vccd1 vccd1 _14523_/D sky130_fd_sc_hd__mux2_1
XFILLER_67_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_59_clk _15031_/CLK vssd1 vssd1 vccd1 vccd1 _15041_/CLK sky130_fd_sc_hd__clkbuf_16
X_14946_ _15570_/CLK _14946_/D vssd1 vssd1 vccd1 vccd1 _14946_/Q sky130_fd_sc_hd__dfxtp_1
X_10069_ _14425_/Q _11680_/A0 _10092_/S vssd1 vssd1 vccd1 vccd1 _14425_/D sky130_fd_sc_hd__mux2_1
XFILLER_36_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14877_ _15422_/CLK _14877_/D vssd1 vssd1 vccd1 vccd1 _14877_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13828_ _14373_/CLK _13828_/D vssd1 vssd1 vccd1 vccd1 _13828_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13759_ _14888_/CLK _13759_/D vssd1 vssd1 vccd1 vccd1 _13759_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_43_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07280_ _07280_/A vssd1 vssd1 vccd1 vccd1 _07280_/Y sky130_fd_sc_hd__inv_2
XFILLER_54_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15429_ _15429_/CLK _15429_/D vssd1 vssd1 vccd1 vccd1 _15429_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_163_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_792 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_1055 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_1039 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09921_ _11874_/A1 _14282_/Q _09930_/S vssd1 vssd1 vccd1 vccd1 _14282_/D sky130_fd_sc_hd__mux2_1
XFILLER_113_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_690 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09852_ _14216_/Q _11872_/A1 _09863_/S vssd1 vssd1 vccd1 vccd1 _14216_/D sky130_fd_sc_hd__mux2_1
XTAP_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08803_ _11870_/A1 _13829_/Q _08816_/S vssd1 vssd1 vccd1 vccd1 _13829_/D sky130_fd_sc_hd__mux2_1
XTAP_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09783_ _14150_/Q _13338_/A0 _09795_/S vssd1 vssd1 vccd1 vccd1 _14150_/D sky130_fd_sc_hd__mux2_1
XTAP_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06995_ _15540_/Q _10892_/B _06997_/B _06994_/X vssd1 vssd1 vccd1 vccd1 _14923_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_3109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_1083 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08734_ _13511_/Q _08750_/A2 _08747_/A2 _13543_/Q vssd1 vssd1 vccd1 vccd1 _08734_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_2408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08665_ _14498_/Q _08693_/A2 _08662_/X _08663_/X _08664_/X vssd1 vssd1 vccd1 vccd1
+ _08665_/X sky130_fd_sc_hd__a2111o_4
XANTENNA_109 input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07616_ _13465_/Q _07617_/C _13466_/Q vssd1 vssd1 vccd1 vccd1 _07616_/X sky130_fd_sc_hd__a21o_1
XTAP_1718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08596_ _13602_/Q _08749_/A2 _08685_/A2 _13563_/Q vssd1 vssd1 vccd1 vccd1 _08596_/X
+ sky130_fd_sc_hd__a22o_1
X_07547_ _14736_/Q _07644_/A _07546_/Y _08084_/C1 vssd1 vssd1 vccd1 vccd1 _13447_/D
+ sky130_fd_sc_hd__o211a_1
X_07478_ _14671_/Q _07490_/B _14710_/Q vssd1 vssd1 vccd1 vccd1 _07478_/X sky130_fd_sc_hd__and3_1
XFILLER_139_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09217_ _09449_/B2 _09213_/X _09214_/X _09216_/X vssd1 vssd1 vccd1 vccd1 _09217_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_182_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09148_ _14079_/Q _09231_/A2 _09403_/B1 _14047_/Q _09391_/A vssd1 vssd1 vccd1 vccd1
+ _09148_/X sky130_fd_sc_hd__a221o_1
XFILLER_108_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09079_ _14365_/Q _15181_/Q _13820_/Q _14559_/Q _09190_/S _09429_/S1 vssd1 vssd1
+ vccd1 vccd1 _09080_/B sky130_fd_sc_hd__mux4_1
XFILLER_163_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11110_ _11380_/A _11181_/B _10984_/Y vssd1 vssd1 vccd1 vccd1 _11110_/Y sky130_fd_sc_hd__a21oi_1
X_12090_ _12596_/A _12090_/B _12090_/C vssd1 vssd1 vccd1 vccd1 _12090_/X sky130_fd_sc_hd__and3_1
XFILLER_146_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11041_ _11041_/A _11041_/B vssd1 vssd1 vccd1 vccd1 _11041_/Y sky130_fd_sc_hd__nor2_1
XFILLER_2_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_54 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14800_ _15618_/CLK _14800_/D vssd1 vssd1 vccd1 vccd1 _14800_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12992_ _15477_/Q _13105_/A2 _13025_/B1 _12991_/X vssd1 vssd1 vccd1 vccd1 _15477_/D
+ sky130_fd_sc_hd__a22o_1
XTAP_3621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14731_ _15584_/CLK _14731_/D vssd1 vssd1 vccd1 vccd1 _14731_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11943_ _13877_/Q _14392_/Q _12407_/S vssd1 vssd1 vccd1 vccd1 _11943_/X sky130_fd_sc_hd__mux2_1
XFILLER_55_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14662_ _15634_/CLK _14662_/D vssd1 vssd1 vccd1 vccd1 _14662_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11874_ _15295_/Q _11874_/A1 _11883_/S vssd1 vssd1 vccd1 vccd1 _15295_/D sky130_fd_sc_hd__mux2_1
XFILLER_55_96 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13613_ _15543_/CLK _13613_/D vssd1 vssd1 vccd1 vccd1 _13613_/Q sky130_fd_sc_hd__dfxtp_1
X_10825_ _14857_/Q _07213_/X _10868_/S vssd1 vssd1 vccd1 vccd1 _14857_/D sky130_fd_sc_hd__mux2_1
XTAP_2997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14593_ _15616_/CLK _14593_/D vssd1 vssd1 vccd1 vccd1 hold4/A sky130_fd_sc_hd__dfxtp_2
X_13544_ _15399_/CLK _13544_/D vssd1 vssd1 vccd1 vccd1 _13544_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_164_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10756_ _15420_/Q _14788_/Q _10765_/S vssd1 vssd1 vccd1 vccd1 _14788_/D sky130_fd_sc_hd__mux2_1
XFILLER_13_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13475_ _15398_/CLK _13475_/D vssd1 vssd1 vccd1 vccd1 _13475_/Q sky130_fd_sc_hd__dfxtp_2
X_10687_ _15016_/Q _10717_/A2 _10652_/B _15033_/Q _10717_/C1 vssd1 vssd1 vccd1 vccd1
+ _10687_/X sky130_fd_sc_hd__a221o_1
XFILLER_139_771 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15214_ _15278_/CLK _15214_/D vssd1 vssd1 vccd1 vccd1 _15214_/Q sky130_fd_sc_hd__dfxtp_1
X_12426_ _13898_/Q _14413_/Q _12430_/S vssd1 vssd1 vccd1 vccd1 _12426_/X sky130_fd_sc_hd__mux2_1
XFILLER_126_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15145_ _15278_/CLK _15145_/D vssd1 vssd1 vccd1 vccd1 _15145_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_126_454 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12357_ _13895_/Q _14410_/Q _12541_/S vssd1 vssd1 vccd1 vccd1 _12357_/X sky130_fd_sc_hd__mux2_1
XFILLER_142_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11308_ _11347_/A _11245_/B _11273_/X _11047_/Y _11307_/Y vssd1 vssd1 vccd1 vccd1
+ _11309_/B sky130_fd_sc_hd__a221o_1
XFILLER_141_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15076_ _15108_/CLK _15076_/D vssd1 vssd1 vccd1 vccd1 _15076_/Q sky130_fd_sc_hd__dfxtp_1
X_12288_ _13892_/Q _14407_/Q _12614_/S vssd1 vssd1 vccd1 vccd1 _12288_/X sky130_fd_sc_hd__mux2_1
XFILLER_141_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14027_ _15303_/CLK _14027_/D vssd1 vssd1 vccd1 vccd1 _14027_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11239_ _11639_/A _11239_/B vssd1 vssd1 vccd1 vccd1 _11239_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_95_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_1086 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06780_ _14923_/Q _14922_/Q vssd1 vssd1 vccd1 vccd1 _06782_/C sky130_fd_sc_hd__nand2_1
X_14929_ _15553_/CLK _14929_/D vssd1 vssd1 vccd1 vccd1 _14929_/Q sky130_fd_sc_hd__dfxtp_2
X_08450_ _13755_/Q _12878_/S _08426_/X _08449_/X vssd1 vssd1 vccd1 vccd1 _13755_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_36_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07401_ _13325_/A0 _13389_/Q _07501_/S vssd1 vssd1 vccd1 vccd1 _13389_/D sky130_fd_sc_hd__mux2_1
XFILLER_90_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08381_ _11252_/A _08381_/B vssd1 vssd1 vccd1 vccd1 _08381_/Y sky130_fd_sc_hd__nand2_1
XFILLER_23_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07332_ _15306_/Q _15462_/Q _07340_/S vssd1 vssd1 vccd1 vccd1 _07332_/X sky130_fd_sc_hd__mux2_2
XFILLER_50_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07263_ _07270_/A _07262_/Y _07274_/B vssd1 vssd1 vccd1 vccd1 _07263_/X sky130_fd_sc_hd__a21o_1
XFILLER_137_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09002_ _13944_/Q _13686_/Q _09005_/S vssd1 vssd1 vccd1 vccd1 _09002_/X sky130_fd_sc_hd__mux2_1
XFILLER_118_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_549 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07194_ _13938_/Q _15525_/Q _07334_/S vssd1 vssd1 vccd1 vccd1 _07197_/A sky130_fd_sc_hd__mux2_8
XFILLER_129_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_777 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09904_ _11857_/A1 _14265_/Q _09930_/S vssd1 vssd1 vccd1 vccd1 _14265_/D sky130_fd_sc_hd__mux2_1
Xfanout502 _08237_/A vssd1 vssd1 vccd1 vccd1 _10520_/B2 sky130_fd_sc_hd__buf_6
Xfanout513 _14607_/Q vssd1 vssd1 vccd1 vccd1 _13125_/B sky130_fd_sc_hd__buf_8
Xfanout524 _14605_/Q vssd1 vssd1 vccd1 vccd1 _09466_/A sky130_fd_sc_hd__buf_12
XFILLER_86_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout535 _09511_/S1 vssd1 vssd1 vccd1 vccd1 _08494_/B sky130_fd_sc_hd__buf_12
XFILLER_101_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout546 _09425_/S vssd1 vssd1 vccd1 vccd1 _09190_/S sky130_fd_sc_hd__buf_12
XFILLER_76_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09835_ _14199_/Q _11680_/A0 _09858_/S vssd1 vssd1 vccd1 vccd1 _14199_/D sky130_fd_sc_hd__mux2_1
Xfanout557 _08490_/A1 vssd1 vssd1 vccd1 vccd1 _09535_/S sky130_fd_sc_hd__buf_12
XFILLER_86_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout568 _12515_/C1 vssd1 vssd1 vccd1 vccd1 _08405_/D sky130_fd_sc_hd__buf_12
Xfanout579 _08405_/B vssd1 vssd1 vccd1 vccd1 _06670_/A sky130_fd_sc_hd__buf_12
XFILLER_101_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09766_ _14133_/Q _13321_/A0 _09795_/S vssd1 vssd1 vccd1 vccd1 _14133_/D sky130_fd_sc_hd__mux2_1
XFILLER_6_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06978_ _06969_/A _06977_/Y _06972_/X vssd1 vssd1 vccd1 vccd1 _06978_/Y sky130_fd_sc_hd__o21ai_1
XTAP_2205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08717_ _13513_/Q _08750_/A2 _08750_/B1 _13616_/Q vssd1 vssd1 vccd1 vccd1 _08717_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_73_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09697_ _13319_/A0 _14067_/Q _09723_/S vssd1 vssd1 vccd1 vccd1 _14067_/D sky130_fd_sc_hd__mux2_1
XFILLER_55_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08648_ _13594_/Q _08691_/A2 _08685_/A2 _13555_/Q _08647_/X vssd1 vssd1 vccd1 vccd1
+ _08652_/B sky130_fd_sc_hd__a221o_1
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1055 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08579_ _08722_/A _08579_/B _08579_/C vssd1 vssd1 vccd1 vccd1 _08579_/X sky130_fd_sc_hd__or3_1
XFILLER_30_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_833 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10610_ _14740_/Q _10609_/X _10610_/S vssd1 vssd1 vccd1 vccd1 _14740_/D sky130_fd_sc_hd__mux2_1
XFILLER_179_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11590_ _13217_/A _11598_/B vssd1 vssd1 vccd1 vccd1 _11591_/B sky130_fd_sc_hd__and2_1
Xclkbuf_5_11_0_clk clkbuf_4_5_0_clk/X vssd1 vssd1 vccd1 vccd1 clkbuf_5_11_0_clk/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_168_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10541_ _10541_/A _10541_/B vssd1 vssd1 vccd1 vccd1 _10542_/B sky130_fd_sc_hd__nor2_1
XFILLER_10_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13260_ _15344_/Q _15591_/Q _13300_/S vssd1 vssd1 vccd1 vccd1 _15591_/D sky130_fd_sc_hd__mux2_1
XFILLER_108_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10472_ _10520_/A1 _13783_/Q _13751_/Q _10520_/B2 vssd1 vssd1 vccd1 vccd1 _10472_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_157_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12211_ _12207_/X _12208_/X _12490_/A vssd1 vssd1 vccd1 vccd1 _12211_/X sky130_fd_sc_hd__mux2_1
XFILLER_136_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13191_ _13189_/Y _13190_/X _15564_/Q _13241_/A2 vssd1 vssd1 vccd1 vccd1 _15564_/D
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_157_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_5_26_0_clk clkbuf_5_27_0_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_5_26_0_clk/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_124_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_796 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12142_ _12138_/X _12139_/X _12168_/A vssd1 vssd1 vccd1 vccd1 _12142_/X sky130_fd_sc_hd__mux2_1
XFILLER_123_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12073_ _12069_/X _12070_/X _12582_/A vssd1 vssd1 vccd1 vccd1 _12073_/X sky130_fd_sc_hd__mux2_1
XFILLER_77_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11024_ _11312_/B _11294_/A vssd1 vssd1 vccd1 vccd1 _11024_/X sky130_fd_sc_hd__and2_1
XFILLER_89_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12975_ _10629_/X _14872_/Q _13029_/S vssd1 vssd1 vccd1 vccd1 _12975_/X sky130_fd_sc_hd__mux2_4
XTAP_3451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14714_ _15489_/CLK _14714_/D vssd1 vssd1 vccd1 vccd1 _14714_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_3484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11926_ _11919_/X _11921_/X _11923_/X _11925_/X _12616_/C1 vssd1 vssd1 vccd1 vccd1
+ _11926_/X sky130_fd_sc_hd__o221a_1
XTAP_2750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14645_ _14851_/CLK _14645_/D vssd1 vssd1 vccd1 vccd1 _14645_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11857_ _15278_/Q _11857_/A1 _11883_/S vssd1 vssd1 vccd1 vccd1 _15278_/D sky130_fd_sc_hd__mux2_1
XTAP_2794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10808_ _14840_/Q _07294_/A _12504_/A vssd1 vssd1 vccd1 vccd1 _14840_/D sky130_fd_sc_hd__mux2_1
XFILLER_60_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14576_ _15267_/CLK _14576_/D vssd1 vssd1 vccd1 vccd1 _14576_/Q sky130_fd_sc_hd__dfxtp_1
X_11788_ _15211_/Q _11854_/A1 _11817_/S vssd1 vssd1 vccd1 vccd1 _15211_/D sky130_fd_sc_hd__mux2_1
XFILLER_158_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13527_ _15386_/CLK _13527_/D vssd1 vssd1 vccd1 vccd1 _13527_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10739_ _15403_/Q _14771_/Q _13140_/S vssd1 vssd1 vccd1 vccd1 _14771_/D sky130_fd_sc_hd__mux2_1
XFILLER_173_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13458_ _15381_/CLK _13458_/D vssd1 vssd1 vccd1 vccd1 _13458_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_174_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12409_ _12402_/X _12404_/X _12406_/X _12408_/X _06671_/A vssd1 vssd1 vccd1 vccd1
+ _12409_/X sky130_fd_sc_hd__o221a_1
XFILLER_126_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13389_ _15655_/CLK _13389_/D vssd1 vssd1 vccd1 vccd1 _13389_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15128_ _15669_/CLK _15128_/D vssd1 vssd1 vccd1 vccd1 _15128_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_181_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07950_ _13553_/Q _07961_/C vssd1 vssd1 vccd1 vccd1 _07951_/B sky130_fd_sc_hd__xnor2_1
X_15059_ _15569_/CLK _15059_/D vssd1 vssd1 vccd1 vccd1 _15059_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_142_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06901_ _15375_/Q _06739_/Y _15374_/Q _06741_/Y _06900_/X vssd1 vssd1 vccd1 vccd1
+ _06901_/X sky130_fd_sc_hd__o221a_1
XFILLER_68_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07881_ _13535_/Q _07881_/B vssd1 vssd1 vccd1 vccd1 _07882_/B sky130_fd_sc_hd__xor2_1
XFILLER_29_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09620_ _13994_/Q _13098_/B2 _09628_/S vssd1 vssd1 vccd1 vccd1 _13994_/D sky130_fd_sc_hd__mux2_1
X_06832_ hold8/A _14591_/Q hold4/A vssd1 vssd1 vccd1 vccd1 _08770_/C sky130_fd_sc_hd__or3_1
X_09551_ _14034_/Q _14002_/Q _09551_/S vssd1 vssd1 vccd1 vccd1 _09551_/X sky130_fd_sc_hd__mux2_1
XFILLER_37_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06763_ input21/X vssd1 vssd1 vccd1 vccd1 _06763_/Y sky130_fd_sc_hd__inv_2
X_08502_ _08536_/A _08536_/B _08536_/C vssd1 vssd1 vccd1 vccd1 _08513_/A sky130_fd_sc_hd__or3_4
X_09482_ _13903_/Q _13123_/B _09519_/B1 _14418_/Q _13123_/A vssd1 vssd1 vccd1 vccd1
+ _09482_/X sky130_fd_sc_hd__a221o_1
XFILLER_52_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06694_ _13474_/Q vssd1 vssd1 vccd1 vccd1 _06694_/Y sky130_fd_sc_hd__inv_2
XFILLER_23_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08433_ _14610_/Q _08390_/C _08425_/X _13120_/S vssd1 vssd1 vccd1 vccd1 _08433_/X
+ sky130_fd_sc_hd__a211o_1
X_08364_ _11013_/A _13195_/B vssd1 vssd1 vccd1 vccd1 _11036_/A sky130_fd_sc_hd__nor2_1
XFILLER_20_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_354 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07315_ _13914_/Q _15501_/Q _07339_/S vssd1 vssd1 vccd1 vccd1 _07352_/A sky130_fd_sc_hd__mux2_8
XFILLER_165_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08295_ _07314_/A _10481_/B _08294_/X vssd1 vssd1 vccd1 vccd1 _11399_/A sky130_fd_sc_hd__a21o_4
XFILLER_137_527 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07246_ _13925_/Q _15512_/Q _07334_/S vssd1 vssd1 vccd1 vccd1 _07260_/A sky130_fd_sc_hd__mux2_8
XFILLER_176_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_13 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07177_ _15351_/Q _15058_/Q _07188_/S vssd1 vssd1 vccd1 vccd1 _07177_/X sky130_fd_sc_hd__mux2_8
XFILLER_11_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_232 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_906 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout310 _07448_/X vssd1 vssd1 vccd1 vccd1 _13337_/A0 sky130_fd_sc_hd__buf_6
Xfanout321 _13078_/B2 vssd1 vssd1 vccd1 vccd1 _13332_/A0 sky130_fd_sc_hd__buf_6
XFILLER_28_1062 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout332 _07408_/X vssd1 vssd1 vccd1 vccd1 _11860_/A1 sky130_fd_sc_hd__buf_4
Xfanout343 _07388_/X vssd1 vssd1 vccd1 vccd1 _13322_/A0 sky130_fd_sc_hd__buf_6
Xfanout354 _10733_/A2 vssd1 vssd1 vccd1 vccd1 _10718_/A2 sky130_fd_sc_hd__buf_12
Xfanout365 _08512_/B vssd1 vssd1 vccd1 vccd1 _09519_/B1 sky130_fd_sc_hd__buf_12
Xfanout376 _11356_/C vssd1 vssd1 vccd1 vccd1 _11023_/A sky130_fd_sc_hd__buf_6
XFILLER_143_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09818_ _14184_/Q _13340_/A0 _09828_/S vssd1 vssd1 vccd1 vccd1 _14184_/D sky130_fd_sc_hd__mux2_1
XFILLER_98_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout387 _11047_/B vssd1 vssd1 vccd1 vccd1 _11115_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_46_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout398 _11298_/A vssd1 vssd1 vccd1 vccd1 _11129_/A sky130_fd_sc_hd__buf_12
XFILLER_101_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_162 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09749_ _14117_/Q _13337_/A0 _09762_/S vssd1 vssd1 vccd1 vccd1 _14117_/D sky130_fd_sc_hd__mux2_1
XTAP_2002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12760_ _12743_/A _12758_/X _12759_/X _12788_/C1 vssd1 vssd1 vccd1 vccd1 _15356_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_2035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11711_ _15140_/Q _11852_/A1 _11741_/S vssd1 vssd1 vccd1 vccd1 _15140_/D sky130_fd_sc_hd__mux2_1
XTAP_1334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_282 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12691_ _13591_/Q _12690_/X _12763_/S vssd1 vssd1 vccd1 vccd1 _12691_/X sky130_fd_sc_hd__mux2_1
XTAP_1356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14430_ _15244_/CLK _14430_/D vssd1 vssd1 vccd1 vccd1 _14430_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_42_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11642_ _15075_/Q _15539_/Q _12904_/S vssd1 vssd1 vccd1 vccd1 _15075_/D sky130_fd_sc_hd__mux2_1
XFILLER_74_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_691 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14361_ _15142_/CLK _14361_/D vssd1 vssd1 vccd1 vccd1 _14361_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_168_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11573_ _11564_/A _11566_/X _11576_/D vssd1 vssd1 vccd1 vccd1 _11573_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_35_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput18 ext_read_data[25] vssd1 vssd1 vccd1 vccd1 input18/X sky130_fd_sc_hd__buf_6
XFILLER_167_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13312_ _15643_/Q _12805_/B _13316_/S vssd1 vssd1 vccd1 vccd1 _15643_/D sky130_fd_sc_hd__mux2_1
X_10524_ _13214_/A _13215_/B vssd1 vssd1 vccd1 vccd1 _10524_/X sky130_fd_sc_hd__and2b_1
XFILLER_10_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput29 ext_read_data[6] vssd1 vssd1 vccd1 vccd1 input29/X sky130_fd_sc_hd__buf_6
XFILLER_182_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14292_ _15172_/CLK _14292_/D vssd1 vssd1 vccd1 vccd1 _14292_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_122_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13243_ _13242_/A _13242_/B _13252_/B _11616_/A vssd1 vssd1 vccd1 vccd1 _13243_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_182_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10455_ _10455_/A _13229_/B vssd1 vssd1 vccd1 vccd1 _10470_/B sky130_fd_sc_hd__and2_1
XFILLER_155_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13174_ _13242_/A _11399_/A _11414_/C vssd1 vssd1 vccd1 vccd1 _13174_/Y sky130_fd_sc_hd__a21oi_1
X_10386_ _07294_/A _10360_/B _10385_/X vssd1 vssd1 vccd1 vccd1 _11476_/B sky130_fd_sc_hd__a21oi_4
XFILLER_124_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12125_ _13949_/Q _13691_/Q _12476_/S vssd1 vssd1 vccd1 vccd1 _12126_/B sky130_fd_sc_hd__mux2_1
XFILLER_97_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12056_ _13946_/Q _13688_/Q _12453_/S vssd1 vssd1 vccd1 vccd1 _12057_/B sky130_fd_sc_hd__mux2_1
XFILLER_111_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11007_ _11053_/S _11007_/B _11324_/A vssd1 vssd1 vccd1 vccd1 _11007_/X sky130_fd_sc_hd__and3_1
XFILLER_42_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12958_ _07392_/X _13024_/A2 _12957_/X _13024_/B2 vssd1 vssd1 vccd1 vccd1 _12958_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_3281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11909_ _14455_/Q _14423_/Q _13844_/Q _14197_/Q _08405_/A _12379_/A vssd1 vssd1 vccd1
+ vccd1 _11909_/X sky130_fd_sc_hd__mux4_1
X_15677_ _15677_/CLK _15677_/D vssd1 vssd1 vccd1 vccd1 _15677_/Q sky130_fd_sc_hd__dfxtp_1
X_12889_ _15417_/Q _15602_/Q _12928_/S vssd1 vssd1 vccd1 vccd1 _15417_/D sky130_fd_sc_hd__mux2_1
XTAP_2580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14628_ _15599_/CLK _14628_/D vssd1 vssd1 vccd1 vccd1 _14628_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14559_ _15218_/CLK _14559_/D vssd1 vssd1 vccd1 vccd1 _14559_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07100_ _07104_/C _07163_/A vssd1 vssd1 vccd1 vccd1 _07131_/A sky130_fd_sc_hd__and2b_4
XFILLER_173_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08080_ _14732_/Q _15205_/Q _06825_/B _06819_/X vssd1 vssd1 vccd1 vccd1 _08080_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_119_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07031_ _07030_/X _13589_/Q _12728_/S vssd1 vssd1 vccd1 vccd1 _07031_/X sky130_fd_sc_hd__mux2_1
XFILLER_162_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_582 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08982_ _14007_/Q _13975_/Q _09132_/S vssd1 vssd1 vccd1 vccd1 _08982_/X sky130_fd_sc_hd__mux2_1
XFILLER_130_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07933_ _08012_/A2 _07932_/X input35/X vssd1 vssd1 vccd1 vccd1 _07933_/Y sky130_fd_sc_hd__a21oi_1
X_07864_ _07866_/B _07863_/X _07874_/A vssd1 vssd1 vccd1 vccd1 _07864_/X sky130_fd_sc_hd__a21bo_1
XFILLER_69_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09603_ _13977_/Q _13325_/A0 _09628_/S vssd1 vssd1 vccd1 vccd1 _13977_/D sky130_fd_sc_hd__mux2_1
X_06815_ _06666_/Y _13049_/A1 _06809_/X _06812_/X _06814_/Y vssd1 vssd1 vccd1 vccd1
+ _06815_/X sky130_fd_sc_hd__o2111a_1
X_07795_ _13511_/Q _07802_/C _13512_/Q vssd1 vssd1 vccd1 vccd1 _07795_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_37_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09534_ _14258_/Q _14290_/Q _14322_/Q _14354_/Q _09535_/S _08494_/B vssd1 vssd1 vccd1
+ vccd1 _09534_/X sky130_fd_sc_hd__mux4_1
X_06746_ _13481_/Q vssd1 vssd1 vccd1 vccd1 _06746_/Y sky130_fd_sc_hd__inv_2
XFILLER_36_271 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09465_ _14383_/Q _15199_/Q _13838_/Q _14577_/Q _09469_/S _13144_/A0 vssd1 vssd1
+ vccd1 vccd1 _09466_/B sky130_fd_sc_hd__mux4_1
XFILLER_19_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06677_ _14906_/Q vssd1 vssd1 vccd1 vccd1 _06845_/B sky130_fd_sc_hd__inv_2
XFILLER_184_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_1039 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08416_ _08477_/C _06991_/B _08415_/X _13138_/S _14929_/D vssd1 vssd1 vccd1 vccd1
+ _13740_/D sky130_fd_sc_hd__o32a_1
XFILLER_169_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09396_ _09406_/S1 _09419_/A2 _09395_/X _06676_/A vssd1 vssd1 vccd1 vccd1 _09396_/X
+ sky130_fd_sc_hd__a31o_1
X_08347_ _08328_/X _08346_/X _11088_/S vssd1 vssd1 vccd1 vccd1 _08381_/B sky130_fd_sc_hd__mux2_1
XFILLER_138_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08278_ _13168_/B vssd1 vssd1 vccd1 vccd1 _11383_/A sky130_fd_sc_hd__inv_2
XFILLER_138_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07229_ _07219_/X _07221_/Y _07227_/A _07227_/B vssd1 vssd1 vccd1 vccd1 _07230_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_153_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_1091 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10240_ _14625_/Q _14778_/Q _10650_/S vssd1 vssd1 vccd1 vccd1 _14625_/D sky130_fd_sc_hd__mux2_1
XFILLER_3_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_254_clk clkbuf_5_0_0_clk/X vssd1 vssd1 vccd1 vccd1 _15273_/CLK sky130_fd_sc_hd__clkbuf_16
X_10171_ _11857_/A1 _14555_/Q _10197_/S vssd1 vssd1 vccd1 vccd1 _14555_/D sky130_fd_sc_hd__mux2_1
XFILLER_79_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout140 _12320_/A vssd1 vssd1 vccd1 vccd1 _12504_/A sky130_fd_sc_hd__clkbuf_8
Xfanout151 _12885_/S vssd1 vssd1 vccd1 vccd1 _12910_/S sky130_fd_sc_hd__buf_6
Xfanout162 _06781_/X vssd1 vssd1 vccd1 vccd1 _08626_/S sky130_fd_sc_hd__clkbuf_16
X_13930_ _15517_/CLK _13930_/D vssd1 vssd1 vccd1 vccd1 _13930_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout173 _11743_/X vssd1 vssd1 vccd1 vccd1 _11774_/S sky130_fd_sc_hd__buf_12
XFILLER_75_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout184 _10099_/X vssd1 vssd1 vccd1 vccd1 _10124_/S sky130_fd_sc_hd__buf_12
Xfanout195 _09898_/Y vssd1 vssd1 vccd1 vccd1 _09925_/S sky130_fd_sc_hd__buf_12
XFILLER_47_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13861_ _15301_/CLK _13861_/D vssd1 vssd1 vccd1 vccd1 _13861_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_170_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15600_ _15634_/CLK _15600_/D vssd1 vssd1 vccd1 vccd1 _15600_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12812_ _12819_/B _12812_/B vssd1 vssd1 vccd1 vccd1 _12813_/B sky130_fd_sc_hd__nor2_1
X_13792_ _15608_/CLK _13792_/D vssd1 vssd1 vccd1 vccd1 _13792_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_16_956 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15531_ _15537_/CLK _15531_/D vssd1 vssd1 vccd1 vccd1 hold1/A sky130_fd_sc_hd__dfxtp_1
X_12743_ _12743_/A _12743_/B vssd1 vssd1 vccd1 vccd1 _12743_/X sky130_fd_sc_hd__or2_1
XTAP_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15462_ _15462_/CLK _15462_/D vssd1 vssd1 vccd1 vccd1 _15462_/Q sky130_fd_sc_hd__dfxtp_1
X_12674_ _15052_/Q _12673_/X _12792_/B vssd1 vssd1 vccd1 vccd1 _12674_/X sky130_fd_sc_hd__mux2_1
XTAP_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14413_ _15527_/CLK _14413_/D vssd1 vssd1 vccd1 vccd1 _14413_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_187_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11625_ _11626_/A _11626_/B vssd1 vssd1 vccd1 vccd1 _11625_/Y sky130_fd_sc_hd__nor2_1
XFILLER_156_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15393_ _15393_/CLK _15393_/D vssd1 vssd1 vccd1 vccd1 _15393_/Q sky130_fd_sc_hd__dfxtp_1
X_14344_ _15293_/CLK _14344_/D vssd1 vssd1 vccd1 vccd1 _14344_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_184_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11556_ _11556_/A _11556_/B vssd1 vssd1 vccd1 vccd1 _11576_/B sky130_fd_sc_hd__nand2_1
XFILLER_155_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10507_ _10507_/A1 _13754_/Q _15418_/Q _10515_/B2 vssd1 vssd1 vccd1 vccd1 _10507_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_183_474 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14275_ _15306_/CLK _14275_/D vssd1 vssd1 vccd1 vccd1 _14275_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_171_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11487_ _11496_/A _11496_/C _10362_/X _13233_/A vssd1 vssd1 vccd1 vccd1 _11491_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_6_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13226_ _13242_/A _13226_/B vssd1 vssd1 vccd1 vccd1 _13226_/Y sky130_fd_sc_hd__nor2_1
XFILLER_6_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10438_ _08244_/A _13745_/Q _15427_/Q _14195_/Q vssd1 vssd1 vccd1 vccd1 _10438_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_152_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_245_clk clkbuf_5_4_0_clk/X vssd1 vssd1 vccd1 vccd1 _15665_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13157_ _13251_/A _10895_/B _11360_/A _11011_/Y _13219_/S vssd1 vssd1 vccd1 vccd1
+ _13157_/X sky130_fd_sc_hd__o221a_1
X_10369_ _11419_/A _11436_/A vssd1 vssd1 vccd1 vccd1 _10382_/A sky130_fd_sc_hd__xor2_1
XTAP_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12108_ _14076_/Q _14044_/Q _12476_/S vssd1 vssd1 vccd1 vccd1 _12108_/X sky130_fd_sc_hd__mux2_1
XTAP_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13088_ _12999_/X _13118_/A2 _13114_/B1 _07448_/X vssd1 vssd1 vccd1 vccd1 _13088_/X
+ sky130_fd_sc_hd__a22o_1
X_12039_ _14073_/Q _14041_/Q _12591_/S vssd1 vssd1 vccd1 vccd1 _12039_/X sky130_fd_sc_hd__mux2_1
XFILLER_111_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_4_1_0_clk clkbuf_4_1_0_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_5_3_0_clk/A sky130_fd_sc_hd__clkbuf_8
XFILLER_25_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07580_ _13456_/Q _07588_/D vssd1 vssd1 vccd1 vccd1 _07583_/B sky130_fd_sc_hd__and2_1
XFILLER_81_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09250_ _14084_/Q _09522_/A2 _09519_/B1 _14052_/Q _09532_/A vssd1 vssd1 vccd1 vccd1
+ _09250_/X sky130_fd_sc_hd__a221o_1
X_08201_ _13692_/Q _13074_/B2 _08216_/S vssd1 vssd1 vccd1 vccd1 _13692_/D sky130_fd_sc_hd__mux2_1
XFILLER_178_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09181_ _09435_/A _09181_/B vssd1 vssd1 vccd1 vccd1 _09181_/X sky130_fd_sc_hd__or2_1
XFILLER_144_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08132_ _13659_/Q _10285_/S _08119_/X _08131_/X vssd1 vssd1 vccd1 vccd1 _13659_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_30_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08063_ _14756_/Q _13634_/Q _08066_/S vssd1 vssd1 vccd1 vccd1 _13634_/D sky130_fd_sc_hd__mux2_1
XFILLER_88_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07014_ _07013_/X _14737_/Q _07098_/S vssd1 vssd1 vccd1 vccd1 _13583_/D sky130_fd_sc_hd__mux2_1
XFILLER_162_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_236_clk clkbuf_5_5_0_clk/X vssd1 vssd1 vccd1 vccd1 _15303_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_161_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08965_ _09530_/S1 _08963_/X _08964_/X vssd1 vssd1 vccd1 vccd1 _08965_/X sky130_fd_sc_hd__a21o_1
XFILLER_102_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07916_ _14736_/Q _08022_/B _07915_/Y _08016_/C1 vssd1 vssd1 vccd1 vccd1 _13543_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_25_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08896_ _13939_/Q _13681_/Q _09230_/S vssd1 vssd1 vccd1 vccd1 _08896_/X sky130_fd_sc_hd__mux2_1
XFILLER_84_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07847_ _13526_/Q _13525_/Q _13524_/Q _07847_/D vssd1 vssd1 vccd1 vccd1 _07858_/D
+ sky130_fd_sc_hd__and4_2
XFILLER_25_1098 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07778_ _14765_/Q _07777_/A _07777_/Y _08016_/C1 vssd1 vssd1 vccd1 vccd1 _13508_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_140_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09517_ _13936_/Q _13093_/A2 _09516_/X vssd1 vssd1 vccd1 vccd1 _13936_/D sky130_fd_sc_hd__a21o_1
X_06729_ _13457_/Q vssd1 vssd1 vccd1 vccd1 _06729_/Y sky130_fd_sc_hd__inv_2
XPHY_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09448_ _14544_/Q _14157_/Q _14189_/Q _14125_/Q _09441_/S _09448_/S1 vssd1 vssd1
+ vccd1 vccd1 _09448_/X sky130_fd_sc_hd__mux4_1
XPHY_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09379_ _14026_/Q _13994_/Q _09512_/S vssd1 vssd1 vccd1 vccd1 _09379_/X sky130_fd_sc_hd__mux2_1
X_11410_ _11421_/B _11410_/B vssd1 vssd1 vccd1 vccd1 _11423_/D sky130_fd_sc_hd__and2b_1
XFILLER_166_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12390_ _15327_/Q _13154_/S _12389_/X vssd1 vssd1 vccd1 vccd1 _15327_/D sky130_fd_sc_hd__a21o_1
XFILLER_123_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11341_ _11013_/A _11633_/A _10963_/A _11259_/S vssd1 vssd1 vccd1 vccd1 _11341_/Y
+ sky130_fd_sc_hd__o211ai_4
XFILLER_153_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14060_ _14405_/CLK _14060_/D vssd1 vssd1 vccd1 vccd1 _14060_/Q sky130_fd_sc_hd__dfxtp_1
X_11272_ _11272_/A _11272_/B vssd1 vssd1 vccd1 vccd1 _11272_/Y sky130_fd_sc_hd__nor2_1
XFILLER_118_390 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13011_ _10689_/X _14884_/Q _13029_/S vssd1 vssd1 vccd1 vccd1 _13011_/X sky130_fd_sc_hd__mux2_4
Xclkbuf_leaf_227_clk clkbuf_5_7_0_clk/X vssd1 vssd1 vccd1 vccd1 _15518_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_3_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10223_ input18/X _14608_/Q _13291_/S vssd1 vssd1 vccd1 vccd1 _14608_/D sky130_fd_sc_hd__mux2_1
XFILLER_180_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10154_ _14539_/Q _13340_/A0 _10164_/S vssd1 vssd1 vccd1 vccd1 _14539_/D sky130_fd_sc_hd__mux2_1
XFILLER_48_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14962_ _14966_/CLK _14962_/D vssd1 vssd1 vccd1 vccd1 _14962_/Q sky130_fd_sc_hd__dfxtp_1
Xhold7 hold7/A vssd1 vssd1 vccd1 vccd1 hold7/X sky130_fd_sc_hd__bufbuf_16
X_10085_ _14441_/Q _11838_/A1 _10097_/S vssd1 vssd1 vccd1 vccd1 _14441_/D sky130_fd_sc_hd__mux2_1
XFILLER_48_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13913_ _15673_/CLK _13913_/D vssd1 vssd1 vccd1 vccd1 _13913_/Q sky130_fd_sc_hd__dfxtp_1
X_14893_ _15646_/CLK _14893_/D vssd1 vssd1 vccd1 vccd1 _14893_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_74_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_40 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13844_ _14197_/CLK _13844_/D vssd1 vssd1 vccd1 vccd1 _13844_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13775_ _14517_/CLK _13775_/D vssd1 vssd1 vccd1 vccd1 _13775_/Q sky130_fd_sc_hd__dfxtp_4
X_10987_ _11330_/A _10987_/B vssd1 vssd1 vccd1 vccd1 _10987_/X sky130_fd_sc_hd__or2_1
XFILLER_43_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_786 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12726_ _15059_/Q _12725_/Y _12792_/B vssd1 vssd1 vccd1 vccd1 _12726_/X sky130_fd_sc_hd__mux2_1
X_15514_ _15523_/CLK _15514_/D vssd1 vssd1 vccd1 vccd1 _15514_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_90 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15445_ _15628_/CLK _15445_/D vssd1 vssd1 vccd1 vccd1 _15445_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_148_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12657_ _15343_/Q _15342_/Q _12657_/C vssd1 vssd1 vccd1 vccd1 _12666_/B sky130_fd_sc_hd__and3_2
XFILLER_90_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11608_ _15069_/Q _11614_/S _11607_/X vssd1 vssd1 vccd1 vccd1 _15069_/D sky130_fd_sc_hd__a21bo_1
XFILLER_12_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15376_ _15377_/CLK _15376_/D vssd1 vssd1 vccd1 vccd1 _15376_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12588_ _12592_/A1 _12587_/X _12548_/S vssd1 vssd1 vccd1 vccd1 _12588_/X sky130_fd_sc_hd__a21o_1
XFILLER_30_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xwire360 wire360/A vssd1 vssd1 vccd1 vccd1 wire360/X sky130_fd_sc_hd__buf_6
X_14327_ _15276_/CLK _14327_/D vssd1 vssd1 vccd1 vccd1 _14327_/Q sky130_fd_sc_hd__dfxtp_1
X_11539_ _13218_/A _11539_/B vssd1 vssd1 vccd1 vccd1 _11541_/B sky130_fd_sc_hd__xnor2_1
XFILLER_128_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14258_ _15672_/CLK _14258_/D vssd1 vssd1 vccd1 vccd1 _14258_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_218_clk clkbuf_5_18_0_clk/X vssd1 vssd1 vccd1 vccd1 _15336_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_98_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13209_ _13233_/A _13208_/B _13241_/A2 _11536_/A vssd1 vssd1 vccd1 vccd1 _13209_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_48_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14189_ _15675_/CLK _14189_/D vssd1 vssd1 vccd1 vccd1 _14189_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_112_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08750_ _13509_/Q _08750_/A2 _08750_/B1 _13612_/Q _08749_/X vssd1 vssd1 vccd1 vccd1
+ _08751_/C sky130_fd_sc_hd__a221o_1
XTAP_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07701_ _13488_/Q _13487_/Q _13486_/Q _13485_/Q vssd1 vssd1 vccd1 vccd1 _07717_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_78_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08681_ _10765_/S _08681_/B _08681_/C vssd1 vssd1 vccd1 vccd1 _08681_/X sky130_fd_sc_hd__or3_4
XFILLER_26_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07632_ _13470_/Q _13469_/Q _07655_/A vssd1 vssd1 vccd1 vccd1 _07635_/B sky130_fd_sc_hd__and3_1
XFILLER_0_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07563_ _13452_/Q _07576_/C vssd1 vssd1 vccd1 vccd1 _07567_/B sky130_fd_sc_hd__nand2_2
XFILLER_94_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09302_ _09300_/X _09301_/X _12573_/A _09291_/X vssd1 vssd1 vccd1 vccd1 _09302_/X
+ sky130_fd_sc_hd__o211a_2
XFILLER_22_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_712 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07494_ _14675_/Q _07498_/B _07498_/C vssd1 vssd1 vccd1 vccd1 _07494_/X sky130_fd_sc_hd__and3_1
XFILLER_167_706 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09233_ _15124_/Q _15092_/Q _15665_/Q _13399_/Q _09230_/S _09234_/S1 vssd1 vssd1
+ vccd1 vccd1 _09233_/X sky130_fd_sc_hd__mux4_1
XFILLER_181_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09164_ _14241_/Q _14273_/Q _14305_/Q _14337_/Q _09444_/S _09446_/A1 vssd1 vssd1
+ vccd1 vccd1 _09164_/X sky130_fd_sc_hd__mux4_1
XFILLER_119_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08115_ _13655_/Q _10344_/S _08096_/X _08114_/X vssd1 vssd1 vccd1 vccd1 _13655_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_175_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09095_ _09130_/A _09088_/X _09091_/X _09450_/B1 vssd1 vssd1 vccd1 vccd1 _09095_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_134_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08046_ _14739_/Q _13617_/Q _08072_/S vssd1 vssd1 vccd1 vccd1 _13617_/D sky130_fd_sc_hd__mux2_1
XFILLER_162_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_209_clk clkbuf_5_16_0_clk/X vssd1 vssd1 vccd1 vccd1 _15672_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_116_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09997_ _14714_/Q _14716_/Q _11743_/C _11851_/A vssd1 vssd1 vccd1 vccd1 _09997_/X
+ sky130_fd_sc_hd__or4_4
XFILLER_76_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08948_ _08668_/D _08944_/X _08947_/X _08943_/X vssd1 vssd1 vccd1 vccd1 _08949_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_85_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08879_ _13900_/Q _13344_/A0 _08880_/S vssd1 vssd1 vccd1 vccd1 _13900_/D sky130_fd_sc_hd__mux2_1
XTAP_3825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10910_ _11436_/A _10944_/B vssd1 vssd1 vccd1 vccd1 _10910_/Y sky130_fd_sc_hd__nand2_1
XFILLER_84_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11890_ _14356_/Q _15172_/Q _13811_/Q _14550_/Q _12154_/S _12253_/S1 vssd1 vssd1
+ vccd1 vccd1 _11890_/X sky130_fd_sc_hd__mux4_1
XFILLER_71_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10841_ _14873_/Q _13795_/Q _12900_/S vssd1 vssd1 vccd1 vccd1 _14873_/D sky130_fd_sc_hd__mux2_1
XFILLER_25_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_1103 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13560_ _13632_/CLK _13560_/D vssd1 vssd1 vccd1 vccd1 _13560_/Q sky130_fd_sc_hd__dfxtp_1
X_10772_ _14804_/Q _15436_/Q _12910_/S vssd1 vssd1 vccd1 vccd1 _14804_/D sky130_fd_sc_hd__mux2_1
XFILLER_40_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12511_ _14383_/Q _15199_/Q _13838_/Q _14577_/Q _12522_/S _12521_/A vssd1 vssd1 vccd1
+ vccd1 _12511_/X sky130_fd_sc_hd__mux4_1
X_13491_ _15383_/CLK _13491_/D vssd1 vssd1 vccd1 vccd1 _13491_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_9_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15230_ _15544_/CLK _15230_/D vssd1 vssd1 vccd1 vccd1 _15230_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_185_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12442_ _14380_/Q _15196_/Q _13835_/Q _14574_/Q _12453_/S _12061_/A vssd1 vssd1 vccd1
+ vccd1 _12442_/X sky130_fd_sc_hd__mux4_1
XFILLER_139_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15161_ _15161_/CLK _15161_/D vssd1 vssd1 vccd1 vccd1 _15161_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_176_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12373_ _14377_/Q _15193_/Q _13832_/Q _14571_/Q _12518_/S _12521_/A vssd1 vssd1 vccd1
+ vccd1 _12373_/X sky130_fd_sc_hd__mux4_1
XFILLER_138_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14112_ _15286_/CLK _14112_/D vssd1 vssd1 vccd1 vccd1 _14112_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_125_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11324_ _11324_/A _11324_/B vssd1 vssd1 vccd1 vccd1 _11324_/Y sky130_fd_sc_hd__nand2_1
XFILLER_176_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15092_ _15665_/CLK _15092_/D vssd1 vssd1 vccd1 vccd1 _15092_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_181_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14043_ _14083_/CLK _14043_/D vssd1 vssd1 vccd1 vccd1 _14043_/Q sky130_fd_sc_hd__dfxtp_1
X_11255_ _11283_/A _08330_/X _11254_/Y _08233_/B vssd1 vssd1 vccd1 vccd1 _11255_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_69_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10206_ input31/X _14591_/Q _13284_/S vssd1 vssd1 vccd1 vccd1 _14591_/D sky130_fd_sc_hd__mux2_1
XFILLER_68_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11186_ _14985_/Q _11202_/A _11170_/X _11185_/Y vssd1 vssd1 vccd1 vccd1 _14985_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_122_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10137_ _14522_/Q _11681_/A0 _10159_/S vssd1 vssd1 vccd1 vccd1 _14522_/D sky130_fd_sc_hd__mux2_1
X_14945_ _15570_/CLK _14945_/D vssd1 vssd1 vccd1 vccd1 _14945_/Q sky130_fd_sc_hd__dfxtp_1
X_10068_ _14424_/Q _13321_/A0 _10097_/S vssd1 vssd1 vccd1 vccd1 _14424_/D sky130_fd_sc_hd__mux2_1
XFILLER_78_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14876_ _15592_/CLK _14876_/D vssd1 vssd1 vccd1 vccd1 _14876_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_165_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_1069 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13827_ _15289_/CLK _13827_/D vssd1 vssd1 vccd1 vccd1 _13827_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13758_ _14888_/CLK _13758_/D vssd1 vssd1 vccd1 vccd1 _13758_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12709_ _15350_/Q _12710_/B vssd1 vssd1 vccd1 vccd1 _12723_/C sky130_fd_sc_hd__and2_1
XFILLER_188_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13689_ _15281_/CLK _13689_/D vssd1 vssd1 vccd1 vccd1 _13689_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15428_ _15589_/CLK _15428_/D vssd1 vssd1 vccd1 vccd1 _15428_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_157_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15359_ _15641_/CLK _15359_/D vssd1 vssd1 vccd1 vccd1 _15359_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_172_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_1067 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09920_ _13340_/A0 _14281_/Q _09930_/S vssd1 vssd1 vccd1 vccd1 _14281_/D sky130_fd_sc_hd__mux2_1
XFILLER_144_499 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09851_ _14215_/Q _11838_/A1 _09863_/S vssd1 vssd1 vccd1 vccd1 _14215_/D sky130_fd_sc_hd__mux2_1
XTAP_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08802_ _11761_/A0 _13828_/Q _08816_/S vssd1 vssd1 vccd1 vccd1 _13828_/D sky130_fd_sc_hd__mux2_1
XFILLER_98_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09782_ _14149_/Q _07448_/X _09795_/S vssd1 vssd1 vccd1 vccd1 _14149_/D sky130_fd_sc_hd__mux2_1
XFILLER_85_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06994_ _14923_/Q _12904_/S vssd1 vssd1 vccd1 vccd1 _06994_/X sky130_fd_sc_hd__or2_1
XTAP_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08733_ _15370_/Q _08748_/A2 _08748_/B1 _14488_/Q vssd1 vssd1 vccd1 vccd1 _08733_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_38_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_1095 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08664_ _13592_/Q _08691_/A2 _08693_/B1 _13624_/Q vssd1 vssd1 vccd1 vccd1 _08664_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_94_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07615_ _14754_/Q _07614_/A _07614_/Y _07987_/C1 vssd1 vssd1 vccd1 vccd1 _13465_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_42_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08595_ _15390_/Q _08748_/A2 _08736_/A2 _13435_/Q vssd1 vssd1 vccd1 vccd1 _08595_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_82_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07546_ _07549_/B _07545_/Y _07644_/A vssd1 vssd1 vccd1 vccd1 _07546_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_34_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07477_ _13344_/A0 _13408_/Q _07481_/S vssd1 vssd1 vccd1 vccd1 _13408_/D sky130_fd_sc_hd__mux2_1
XFILLER_167_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09216_ _15091_/Q _13130_/B1 _08520_/B _09215_/X vssd1 vssd1 vccd1 vccd1 _09216_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_10_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09147_ _14015_/Q _13983_/Q _09407_/S vssd1 vssd1 vccd1 vccd1 _09147_/X sky130_fd_sc_hd__mux2_1
XFILLER_148_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_230 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09078_ _13915_/Q _13119_/S _09077_/X vssd1 vssd1 vccd1 vccd1 _13915_/D sky130_fd_sc_hd__a21o_1
XFILLER_123_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08029_ _14741_/Q _08027_/X _08028_/X _12832_/C1 vssd1 vssd1 vccd1 vccd1 _13573_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_123_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11040_ _11035_/X _11039_/X _11362_/B vssd1 vssd1 vccd1 vccd1 _11136_/B sky130_fd_sc_hd__mux2_1
XFILLER_1_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_66 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12991_ _13082_/B2 _13024_/A2 _12990_/X _13024_/B2 vssd1 vssd1 vccd1 vccd1 _12991_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_3611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11942_ _12544_/A _11942_/B vssd1 vssd1 vccd1 vccd1 _11942_/X sky130_fd_sc_hd__and2_1
X_14730_ _15618_/CLK _14730_/D vssd1 vssd1 vccd1 vccd1 _14730_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_3644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14661_ _15628_/CLK _14661_/D vssd1 vssd1 vccd1 vccd1 _14661_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11873_ _15294_/Q _11873_/A1 _11883_/S vssd1 vssd1 vccd1 vccd1 _15294_/D sky130_fd_sc_hd__mux2_1
XTAP_2954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13612_ _13803_/CLK _13612_/D vssd1 vssd1 vccd1 vccd1 _13612_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10824_ _14856_/Q _07210_/A _13138_/S vssd1 vssd1 vccd1 vccd1 _14856_/D sky130_fd_sc_hd__mux2_1
XTAP_2987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14592_ _15534_/CLK _14592_/D vssd1 vssd1 vccd1 vccd1 _14592_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_2998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13543_ _14517_/CLK _13543_/D vssd1 vssd1 vccd1 vccd1 _13543_/Q sky130_fd_sc_hd__dfxtp_1
X_10755_ _15419_/Q _14787_/Q _10765_/S vssd1 vssd1 vccd1 vccd1 _14787_/D sky130_fd_sc_hd__mux2_1
XFILLER_9_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13474_ _15398_/CLK _13474_/D vssd1 vssd1 vccd1 vccd1 _13474_/Q sky130_fd_sc_hd__dfxtp_2
X_10686_ _15575_/Q _10706_/B vssd1 vssd1 vccd1 vccd1 _10686_/X sky130_fd_sc_hd__and2_1
XFILLER_173_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15213_ _15277_/CLK _15213_/D vssd1 vssd1 vccd1 vccd1 _15213_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_173_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12425_ _12563_/A _12425_/B vssd1 vssd1 vccd1 vccd1 _12425_/X sky130_fd_sc_hd__and2_1
XFILLER_126_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15144_ _15277_/CLK _15144_/D vssd1 vssd1 vccd1 vccd1 _15144_/Q sky130_fd_sc_hd__dfxtp_1
X_12356_ _12540_/A _12356_/B vssd1 vssd1 vccd1 vccd1 _12356_/X sky130_fd_sc_hd__and2_1
XFILLER_127_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11307_ _11307_/A _11307_/B vssd1 vssd1 vccd1 vccd1 _11307_/Y sky130_fd_sc_hd__nor2_1
XFILLER_5_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15075_ _15617_/CLK _15075_/D vssd1 vssd1 vccd1 vccd1 _15075_/Q sky130_fd_sc_hd__dfxtp_1
X_12287_ _12383_/A _12287_/B vssd1 vssd1 vccd1 vccd1 _12287_/X sky130_fd_sc_hd__and2_1
XFILLER_45_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14026_ _15335_/CLK _14026_/D vssd1 vssd1 vccd1 vccd1 _14026_/Q sky130_fd_sc_hd__dfxtp_1
X_11238_ _14929_/D _14927_/D _14928_/D vssd1 vssd1 vccd1 vccd1 _11240_/B sky130_fd_sc_hd__or3b_1
XFILLER_68_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11169_ _14977_/Q _11168_/Y _11202_/A vssd1 vssd1 vccd1 vccd1 _14977_/D sky130_fd_sc_hd__mux2_1
XFILLER_67_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_1098 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14928_ _15553_/CLK _14928_/D vssd1 vssd1 vccd1 vccd1 _14928_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_36_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14859_ _15434_/CLK _14859_/D vssd1 vssd1 vccd1 vccd1 _14859_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07400_ _14740_/Q _07399_/X _07500_/S vssd1 vssd1 vccd1 vccd1 _07400_/X sky130_fd_sc_hd__mux2_8
X_08380_ _13727_/Q _11346_/A2 _11351_/C1 _08379_/X vssd1 vssd1 vccd1 vccd1 _13727_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_17_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07331_ _07331_/A vssd1 vssd1 vccd1 vccd1 _07331_/Y sky130_fd_sc_hd__inv_2
XFILLER_188_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_176_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07262_ _07270_/B _07270_/C vssd1 vssd1 vccd1 vccd1 _07262_/Y sky130_fd_sc_hd__nor2_1
XFILLER_149_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09001_ _08668_/D _08997_/X _09000_/X _08996_/X vssd1 vssd1 vccd1 vccd1 _09014_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_164_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_411 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07193_ _15367_/Q _15074_/Q _07193_/S vssd1 vssd1 vccd1 vccd1 _07193_/X sky130_fd_sc_hd__mux2_8
XFILLER_160_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09903_ _11681_/A0 _14264_/Q _09925_/S vssd1 vssd1 vccd1 vccd1 _14264_/D sky130_fd_sc_hd__mux2_1
Xfanout503 _14766_/Q vssd1 vssd1 vccd1 vccd1 _08237_/A sky130_fd_sc_hd__buf_12
XFILLER_116_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout514 _09405_/A vssd1 vssd1 vccd1 vccd1 _09130_/A sky130_fd_sc_hd__buf_12
XFILLER_59_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_970 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout525 _08988_/A1 vssd1 vssd1 vccd1 vccd1 _09225_/S1 sky130_fd_sc_hd__buf_12
XFILLER_99_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout536 _08487_/A vssd1 vssd1 vccd1 vccd1 _09511_/S1 sky130_fd_sc_hd__buf_12
XFILLER_150_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09834_ _14198_/Q _13321_/A0 _09863_/S vssd1 vssd1 vccd1 vccd1 _14198_/D sky130_fd_sc_hd__mux2_1
Xfanout547 _08490_/A1 vssd1 vssd1 vccd1 vccd1 _09425_/S sky130_fd_sc_hd__buf_12
Xfanout558 _08490_/A1 vssd1 vssd1 vccd1 vccd1 _09512_/S sky130_fd_sc_hd__buf_8
XFILLER_112_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout569 _14602_/Q vssd1 vssd1 vccd1 vccd1 _12515_/C1 sky130_fd_sc_hd__buf_12
XTAP_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09765_ _14132_/Q _13320_/A0 _09795_/S vssd1 vssd1 vccd1 vccd1 _14132_/D sky130_fd_sc_hd__mux2_1
X_06977_ _06977_/A _06977_/B vssd1 vssd1 vccd1 vccd1 _06977_/Y sky130_fd_sc_hd__nor2_1
XFILLER_39_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08716_ _13801_/Q _08715_/X _12932_/S vssd1 vssd1 vccd1 vccd1 _13801_/D sky130_fd_sc_hd__mux2_1
XFILLER_132_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09696_ _11851_/A _09696_/B vssd1 vssd1 vccd1 vccd1 _09696_/X sky130_fd_sc_hd__or2_4
XTAP_2206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08647_ _13459_/Q _08684_/A2 _08683_/A2 _13523_/Q vssd1 vssd1 vccd1 vccd1 _08647_/X
+ sky130_fd_sc_hd__a22o_1
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_250 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08578_ _14511_/Q _08748_/B1 _08576_/X _08577_/X vssd1 vssd1 vccd1 vccd1 _08579_/C
+ sky130_fd_sc_hd__a211o_1
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_136 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07529_ _14759_/Q _13438_/Q _07529_/S vssd1 vssd1 vccd1 vccd1 _13438_/D sky130_fd_sc_hd__mux2_1
XFILLER_41_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_884 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_167_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10540_ _10519_/A _10524_/X _10539_/Y _10526_/B _10512_/B vssd1 vssd1 vccd1 vccd1
+ _10541_/B sky130_fd_sc_hd__o311a_1
XFILLER_22_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_826 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10471_ _10537_/A _10471_/B _10471_/C _10471_/D vssd1 vssd1 vccd1 vccd1 _10557_/B
+ sky130_fd_sc_hd__or4_2
XFILLER_10_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12210_ _15122_/Q _15090_/Q _15663_/Q _13397_/Q _12472_/S _12465_/S1 vssd1 vssd1
+ vccd1 vccd1 _12210_/X sky130_fd_sc_hd__mux4_1
X_13190_ _13229_/A _13189_/B _11476_/A _13241_/A2 vssd1 vssd1 vccd1 vccd1 _13190_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_109_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12141_ _15119_/Q _15087_/Q _15660_/Q _13394_/Q _11993_/S _11992_/A vssd1 vssd1 vccd1
+ vccd1 _12141_/X sky130_fd_sc_hd__mux4_1
XFILLER_124_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12072_ _15116_/Q _15084_/Q _15657_/Q _13391_/Q _12079_/S _12268_/A vssd1 vssd1 vccd1
+ vccd1 _12072_/X sky130_fd_sc_hd__mux4_1
XFILLER_96_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11023_ _11023_/A _13226_/B vssd1 vssd1 vccd1 vccd1 _11294_/A sky130_fd_sc_hd__nand2_1
XFILLER_173_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_943 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12974_ _15471_/Q _13105_/A2 _13025_/B1 _12973_/X vssd1 vssd1 vccd1 vccd1 _15471_/D
+ sky130_fd_sc_hd__a22o_1
XTAP_3441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_656 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14713_ _15489_/CLK _14713_/D vssd1 vssd1 vccd1 vccd1 _14713_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_3474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11925_ _12615_/A1 _11924_/X _12615_/B1 vssd1 vssd1 vccd1 vccd1 _11925_/X sky130_fd_sc_hd__a21o_1
XTAP_3485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11856_ _15277_/Q _13323_/A0 _11878_/S vssd1 vssd1 vccd1 vccd1 _15277_/D sky130_fd_sc_hd__mux2_1
X_14644_ _15429_/CLK _14644_/D vssd1 vssd1 vccd1 vccd1 _14644_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_62 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10807_ _14839_/Q _07301_/A _12481_/A vssd1 vssd1 vccd1 vccd1 _14839_/D sky130_fd_sc_hd__mux2_1
XFILLER_20_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14575_ _15286_/CLK _14575_/D vssd1 vssd1 vccd1 vccd1 _14575_/Q sky130_fd_sc_hd__dfxtp_1
X_11787_ _15210_/Q _13320_/A0 _11817_/S vssd1 vssd1 vccd1 vccd1 _15210_/D sky130_fd_sc_hd__mux2_1
XFILLER_13_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13526_ _13627_/CLK _13526_/D vssd1 vssd1 vccd1 vccd1 _13526_/Q sky130_fd_sc_hd__dfxtp_1
X_10738_ _15402_/Q _14770_/Q _10834_/S vssd1 vssd1 vccd1 vccd1 _14770_/D sky130_fd_sc_hd__mux2_1
XFILLER_186_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13457_ _15381_/CLK _13457_/D vssd1 vssd1 vccd1 vccd1 _13457_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_158_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10669_ _15061_/Q _10714_/A2 _10666_/X _10668_/X vssd1 vssd1 vccd1 vccd1 _10669_/X
+ sky130_fd_sc_hd__o22a_4
XFILLER_173_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12408_ _12592_/A1 _12407_/X _06670_/A vssd1 vssd1 vccd1 vccd1 _12408_/X sky130_fd_sc_hd__a21o_1
XFILLER_161_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13388_ _15654_/CLK _13388_/D vssd1 vssd1 vccd1 vccd1 _13388_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_154_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_892 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15127_ _15127_/CLK _15127_/D vssd1 vssd1 vccd1 vccd1 _15127_/Q sky130_fd_sc_hd__dfxtp_1
X_12339_ _12615_/A1 _12338_/X _12615_/B1 vssd1 vssd1 vccd1 vccd1 _12339_/X sky130_fd_sc_hd__a21o_1
XFILLER_99_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15058_ _15599_/CLK _15058_/D vssd1 vssd1 vccd1 vccd1 _15058_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_99_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14009_ _14572_/CLK _14009_/D vssd1 vssd1 vccd1 vccd1 _14009_/Q sky130_fd_sc_hd__dfxtp_1
X_06900_ _15374_/Q _06741_/Y _15373_/Q _06744_/Y _06899_/X vssd1 vssd1 vccd1 vccd1
+ _06900_/X sky130_fd_sc_hd__a221o_1
X_07880_ _14759_/Q _07874_/A _07879_/X _08002_/C1 vssd1 vssd1 vccd1 vccd1 _13534_/D
+ sky130_fd_sc_hd__o211a_1
X_06831_ _08756_/B _08477_/C vssd1 vssd1 vccd1 vccd1 _08390_/B sky130_fd_sc_hd__and2_2
XFILLER_68_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09550_ _09550_/A1 _09548_/X _09549_/X vssd1 vssd1 vccd1 vccd1 _09554_/B sky130_fd_sc_hd__a21o_1
XFILLER_110_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06762_ input20/X vssd1 vssd1 vccd1 vccd1 _06762_/Y sky130_fd_sc_hd__inv_2
X_08501_ _08501_/A _14609_/Q vssd1 vssd1 vccd1 vccd1 _08536_/C sky130_fd_sc_hd__nand2_1
X_09481_ _13967_/Q _13709_/Q _09481_/S vssd1 vssd1 vccd1 vccd1 _09481_/X sky130_fd_sc_hd__mux2_1
X_06693_ _15397_/Q vssd1 vssd1 vccd1 vccd1 _06693_/Y sky130_fd_sc_hd__inv_2
XFILLER_24_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08432_ _13746_/Q _12878_/S _08426_/B _08431_/X vssd1 vssd1 vccd1 vccd1 _13746_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_168_108 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08363_ _07287_/B _10523_/A2 _08362_/X vssd1 vssd1 vccd1 vccd1 _13195_/B sky130_fd_sc_hd__a21oi_4
XFILLER_23_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07314_ _07314_/A vssd1 vssd1 vccd1 vccd1 _07314_/Y sky130_fd_sc_hd__inv_2
XFILLER_176_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08294_ _08244_/A _13768_/Q _15404_/Q _08244_/B vssd1 vssd1 vccd1 vccd1 _08294_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_149_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_191 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07245_ _07265_/A _07265_/B _07242_/X _07244_/Y vssd1 vssd1 vccd1 vccd1 _07274_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_137_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_25 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07176_ _15350_/Q _15057_/Q _07188_/S vssd1 vssd1 vccd1 vccd1 _07176_/X sky130_fd_sc_hd__mux2_2
XFILLER_118_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout300 _07468_/X vssd1 vssd1 vccd1 vccd1 _13098_/B2 sky130_fd_sc_hd__buf_6
Xfanout311 _07448_/X vssd1 vssd1 vccd1 vccd1 _11870_/A1 sky130_fd_sc_hd__buf_4
XFILLER_99_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout322 _07428_/X vssd1 vssd1 vccd1 vccd1 _13078_/B2 sky130_fd_sc_hd__buf_8
XFILLER_87_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout333 _12967_/A1 vssd1 vssd1 vccd1 vccd1 _13326_/A0 sky130_fd_sc_hd__buf_6
Xfanout344 _07384_/X vssd1 vssd1 vccd1 vccd1 _11854_/A1 sky130_fd_sc_hd__buf_6
XFILLER_28_1074 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout355 _10575_/X vssd1 vssd1 vccd1 vccd1 _10733_/A2 sky130_fd_sc_hd__buf_12
XFILLER_154_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout366 _08508_/Y vssd1 vssd1 vccd1 vccd1 _08512_/B sky130_fd_sc_hd__buf_12
XFILLER_143_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09817_ _14183_/Q _13092_/B2 _09828_/S vssd1 vssd1 vccd1 vccd1 _14183_/D sky130_fd_sc_hd__mux2_1
Xfanout377 _08241_/Y vssd1 vssd1 vccd1 vccd1 _11356_/C sky130_fd_sc_hd__clkbuf_16
XFILLER_100_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout388 _08235_/Y vssd1 vssd1 vccd1 vccd1 _11047_/B sky130_fd_sc_hd__buf_12
XFILLER_47_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout399 _08227_/Y vssd1 vssd1 vccd1 vccd1 _11298_/A sky130_fd_sc_hd__buf_12
XFILLER_100_174 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09748_ _14116_/Q _13086_/B2 _09762_/S vssd1 vssd1 vccd1 vccd1 _14116_/D sky130_fd_sc_hd__mux2_1
XFILLER_185_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09679_ _14050_/Q _13082_/B2 _09690_/S vssd1 vssd1 vccd1 vccd1 _14050_/D sky130_fd_sc_hd__mux2_1
XTAP_2036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11710_ _11710_/A _11851_/B vssd1 vssd1 vccd1 vccd1 _11710_/Y sky130_fd_sc_hd__nor2_8
XTAP_2058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12690_ _15054_/Q _12689_/Y _12792_/B vssd1 vssd1 vccd1 vccd1 _12690_/X sky130_fd_sc_hd__mux2_1
XTAP_1335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11641_ _11640_/Y _15074_/Q _11641_/S vssd1 vssd1 vccd1 vccd1 _15074_/D sky130_fd_sc_hd__mux2_1
XTAP_1379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14360_ _15176_/CLK _14360_/D vssd1 vssd1 vccd1 vccd1 _14360_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11572_ _13226_/B _11572_/B vssd1 vssd1 vccd1 vccd1 _11576_/D sky130_fd_sc_hd__xnor2_4
XFILLER_128_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13311_ _15642_/Q _12799_/B _13316_/S vssd1 vssd1 vccd1 vccd1 _15642_/D sky130_fd_sc_hd__mux2_1
XFILLER_155_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput19 ext_read_data[26] vssd1 vssd1 vccd1 vccd1 input19/X sky130_fd_sc_hd__buf_8
XFILLER_122_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10523_ _07251_/A _10523_/A2 _10522_/X vssd1 vssd1 vccd1 vccd1 _13215_/B sky130_fd_sc_hd__a21oi_4
XFILLER_7_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14291_ _15203_/CLK _14291_/D vssd1 vssd1 vccd1 vccd1 _14291_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_183_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13242_ _13242_/A _13242_/B vssd1 vssd1 vccd1 vccd1 _13242_/Y sky130_fd_sc_hd__nor2_1
X_10454_ _11582_/A _11584_/A vssd1 vssd1 vccd1 vccd1 _13229_/B sky130_fd_sc_hd__nand2_1
XFILLER_171_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13173_ _13171_/Y _13172_/X _15558_/Q _13252_/B vssd1 vssd1 vccd1 vccd1 _15558_/D
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_184_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10385_ _10520_/A1 _13796_/Q _13764_/Q _10520_/B2 vssd1 vssd1 vccd1 vccd1 _10385_/X
+ sky130_fd_sc_hd__a22o_2
XFILLER_123_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12124_ _12503_/A1 _12119_/X _12122_/X _12123_/X _08449_/A vssd1 vssd1 vccd1 vccd1
+ _12136_/B sky130_fd_sc_hd__a221o_1
XFILLER_97_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12055_ _12273_/A1 _12050_/X _12053_/X _12054_/X _08449_/A vssd1 vssd1 vccd1 vccd1
+ _12067_/B sky130_fd_sc_hd__a221o_4
XFILLER_2_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11006_ _11013_/A wire360/X vssd1 vssd1 vccd1 vccd1 _11324_/A sky130_fd_sc_hd__or2_1
XFILLER_77_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_887 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12957_ _10599_/X _14866_/Q _13038_/S vssd1 vssd1 vccd1 vccd1 _12957_/X sky130_fd_sc_hd__mux2_2
XTAP_3282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11908_ _14229_/Q _14261_/Q _14293_/Q _14325_/Q _12522_/S _12521_/A vssd1 vssd1 vccd1
+ vccd1 _11908_/X sky130_fd_sc_hd__mux4_1
X_15676_ _15676_/CLK _15676_/D vssd1 vssd1 vccd1 vccd1 _15676_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12888_ _15416_/Q _15601_/Q _12928_/S vssd1 vssd1 vccd1 vccd1 _15416_/D sky130_fd_sc_hd__mux2_1
XTAP_2581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14627_ _15632_/CLK _14627_/D vssd1 vssd1 vccd1 vccd1 _14627_/Q sky130_fd_sc_hd__dfxtp_1
X_11839_ _15261_/Q _11872_/A1 _11850_/S vssd1 vssd1 vccd1 vccd1 _15261_/D sky130_fd_sc_hd__mux2_1
XTAP_1880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14558_ _15279_/CLK _14558_/D vssd1 vssd1 vccd1 vccd1 _14558_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_174_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13509_ _15615_/CLK _13509_/D vssd1 vssd1 vccd1 vccd1 _13509_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_186_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14489_ _15399_/CLK _14489_/D vssd1 vssd1 vccd1 vccd1 _14489_/Q sky130_fd_sc_hd__dfxtp_2
X_07030_ _14622_/Q _14654_/Q _07078_/S vssd1 vssd1 vccd1 vccd1 _07030_/X sky130_fd_sc_hd__mux2_1
XFILLER_173_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08981_ _08988_/A1 _08979_/X _08980_/X vssd1 vssd1 vccd1 vccd1 _08985_/B sky130_fd_sc_hd__a21o_1
XFILLER_103_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07932_ _13548_/Q _07932_/B vssd1 vssd1 vccd1 vccd1 _07932_/X sky130_fd_sc_hd__xor2_1
XFILLER_60_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07863_ _13530_/Q _07869_/D vssd1 vssd1 vccd1 vccd1 _07863_/X sky130_fd_sc_hd__or2_1
Xclkbuf_5_10_0_clk clkbuf_4_5_0_clk/X vssd1 vssd1 vccd1 vccd1 _15031_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_3_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09602_ _13976_/Q _11857_/A1 _09628_/S vssd1 vssd1 vccd1 vccd1 _13976_/D sky130_fd_sc_hd__mux2_1
XFILLER_56_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06814_ _06664_/Y _09382_/A _06810_/X _06813_/X vssd1 vssd1 vccd1 vccd1 _06814_/Y
+ sky130_fd_sc_hd__a211oi_1
XFILLER_3_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07794_ _13512_/Q _13511_/Q _07802_/C vssd1 vssd1 vccd1 vccd1 _07798_/B sky130_fd_sc_hd__and3_2
X_09533_ _08507_/A _09530_/X _09532_/X _09524_/A vssd1 vssd1 vccd1 vccd1 _09533_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_3_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06745_ _14490_/Q vssd1 vssd1 vccd1 vccd1 _06745_/Y sky130_fd_sc_hd__inv_2
XFILLER_97_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_5_25_0_clk clkbuf_5_25_0_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_5_25_0_clk/X
+ sky130_fd_sc_hd__clkbuf_8
X_09464_ _15300_/Q _15268_/Q _15236_/Q _15167_/Q _09469_/S _09546_/S1 vssd1 vssd1
+ vccd1 vccd1 _09464_/X sky130_fd_sc_hd__mux4_1
X_06676_ _06676_/A vssd1 vssd1 vccd1 vccd1 _13131_/A sky130_fd_sc_hd__inv_8
X_08415_ _14597_/Q _08390_/A _13120_/S vssd1 vssd1 vccd1 vccd1 _08415_/X sky130_fd_sc_hd__a21o_1
X_09395_ _13867_/Q _14220_/Q _09407_/S vssd1 vssd1 vccd1 vccd1 _09395_/X sky130_fd_sc_hd__mux2_1
XFILLER_52_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08346_ _11033_/B _11034_/A vssd1 vssd1 vccd1 vccd1 _08346_/X sky130_fd_sc_hd__or2_1
XFILLER_149_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08277_ _07324_/A _10481_/B _08276_/X vssd1 vssd1 vccd1 vccd1 _13168_/B sky130_fd_sc_hd__a21o_4
XFILLER_165_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07228_ _07228_/A _07228_/B vssd1 vssd1 vccd1 vccd1 _07230_/C sky130_fd_sc_hd__or2_1
XFILLER_125_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07159_ _07163_/A _07159_/B vssd1 vssd1 vccd1 vccd1 _07159_/X sky130_fd_sc_hd__and2_4
XFILLER_133_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10170_ _13323_/A0 _14554_/Q _10192_/S vssd1 vssd1 vccd1 vccd1 _14554_/D sky130_fd_sc_hd__mux2_1
XFILLER_65_1038 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout130 _13093_/A2 vssd1 vssd1 vccd1 vccd1 _10877_/S sky130_fd_sc_hd__clkbuf_16
XFILLER_87_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout141 _10871_/S vssd1 vssd1 vccd1 vccd1 _10868_/S sky130_fd_sc_hd__buf_12
Xfanout152 _12885_/S vssd1 vssd1 vccd1 vccd1 _12900_/S sky130_fd_sc_hd__buf_12
Xfanout163 _13318_/X vssd1 vssd1 vccd1 vccd1 _13345_/S sky130_fd_sc_hd__buf_12
XFILLER_93_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout174 _11743_/X vssd1 vssd1 vccd1 vccd1 _11775_/S sky130_fd_sc_hd__buf_12
XFILLER_86_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout185 _10065_/Y vssd1 vssd1 vccd1 vccd1 _10092_/S sky130_fd_sc_hd__buf_12
XFILLER_47_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout196 _09898_/Y vssd1 vssd1 vccd1 vccd1 _09930_/S sky130_fd_sc_hd__buf_12
X_13860_ _14373_/CLK _13860_/D vssd1 vssd1 vccd1 vccd1 _13860_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12811_ _15363_/Q _12810_/C _15364_/Q vssd1 vssd1 vccd1 vccd1 _12812_/B sky130_fd_sc_hd__a21oi_1
XFILLER_41_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13791_ _15628_/CLK _13791_/D vssd1 vssd1 vccd1 vccd1 _13791_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_74_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15530_ _15530_/CLK _15530_/D vssd1 vssd1 vccd1 vccd1 _15530_/Q sky130_fd_sc_hd__dfxtp_1
X_12742_ _13431_/Q _12741_/X _12764_/S vssd1 vssd1 vccd1 vccd1 _12743_/B sky130_fd_sc_hd__mux2_1
XTAP_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12673_ _15345_/Q _12679_/C vssd1 vssd1 vccd1 vccd1 _12673_/X sky130_fd_sc_hd__xor2_1
XTAP_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15461_ _15461_/CLK _15461_/D vssd1 vssd1 vccd1 vccd1 _15461_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_169_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_190_clk clkbuf_5_20_0_clk/X vssd1 vssd1 vccd1 vccd1 _15096_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14412_ _15130_/CLK _14412_/D vssd1 vssd1 vccd1 vccd1 _14412_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11624_ _11624_/A _11624_/B vssd1 vssd1 vccd1 vccd1 _11626_/B sky130_fd_sc_hd__xnor2_1
XFILLER_168_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15392_ _15393_/CLK _15392_/D vssd1 vssd1 vccd1 vccd1 _15392_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_184_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11555_ _11555_/A _11555_/B vssd1 vssd1 vccd1 vccd1 _11556_/B sky130_fd_sc_hd__nand2_1
XFILLER_11_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14343_ _15292_/CLK _14343_/D vssd1 vssd1 vccd1 vccd1 _14343_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10506_ _07265_/A _10360_/B _10505_/X vssd1 vssd1 vccd1 vccd1 _13218_/A sky130_fd_sc_hd__a21oi_4
XFILLER_183_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14274_ _14468_/CLK _14274_/D vssd1 vssd1 vccd1 vccd1 _14274_/Q sky130_fd_sc_hd__dfxtp_1
X_11486_ _15057_/Q _11614_/S _11484_/Y _11485_/X vssd1 vssd1 vccd1 vccd1 _15057_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_109_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13225_ _15575_/Q _13219_/S _13224_/X vssd1 vssd1 vccd1 vccd1 _15575_/D sky130_fd_sc_hd__o21a_1
XFILLER_155_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10437_ _07228_/A _10360_/B _10436_/X vssd1 vssd1 vccd1 vccd1 _11624_/A sky130_fd_sc_hd__a21o_4
XFILLER_6_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13156_ _14929_/D _14928_/D _14927_/D vssd1 vssd1 vccd1 vccd1 _13156_/Y sky130_fd_sc_hd__nand3_4
X_10368_ _07306_/A _10360_/B _10367_/X vssd1 vssd1 vccd1 vccd1 _11436_/A sky130_fd_sc_hd__a21oi_4
XTAP_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12107_ _12498_/A _12107_/B vssd1 vssd1 vccd1 vccd1 _12107_/X sky130_fd_sc_hd__and2_1
XFILLER_111_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13087_ _15511_/Q _13093_/A2 _13042_/A _13086_/X vssd1 vssd1 vccd1 vccd1 _15511_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_111_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10299_ _14684_/Q _14869_/Q _10615_/S vssd1 vssd1 vccd1 vccd1 _14684_/D sky130_fd_sc_hd__mux2_1
XFILLER_111_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12038_ _12590_/A _12038_/B vssd1 vssd1 vccd1 vccd1 _12038_/X sky130_fd_sc_hd__and2_1
XFILLER_66_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13989_ _15094_/CLK _13989_/D vssd1 vssd1 vccd1 vccd1 _13989_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15659_ _15659_/CLK _15659_/D vssd1 vssd1 vccd1 vccd1 _15659_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_181_clk clkbuf_5_20_0_clk/X vssd1 vssd1 vccd1 vccd1 _15094_/CLK sky130_fd_sc_hd__clkbuf_16
X_08200_ _13691_/Q _13072_/B2 _08216_/S vssd1 vssd1 vccd1 vccd1 _13691_/D sky130_fd_sc_hd__mux2_1
X_09180_ _14370_/Q _15186_/Q _13825_/Q _14564_/Q _09444_/S _09446_/A1 vssd1 vssd1
+ vccd1 vccd1 _09181_/B sky130_fd_sc_hd__mux4_1
XFILLER_105_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08131_ _08151_/S _08129_/X _08130_/Y _08121_/X vssd1 vssd1 vccd1 vccd1 _08131_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_30_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08062_ _14755_/Q _13633_/Q _08066_/S vssd1 vssd1 vccd1 vccd1 _13633_/D sky130_fd_sc_hd__mux2_1
XFILLER_134_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07013_ _07012_/X _13583_/Q _12640_/S vssd1 vssd1 vccd1 vccd1 _07013_/X sky130_fd_sc_hd__mux2_1
XFILLER_108_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_147 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08964_ _14070_/Q _09231_/A2 _09403_/B1 _14038_/Q _09221_/A vssd1 vssd1 vccd1 vccd1
+ _08964_/X sky130_fd_sc_hd__a221o_1
XFILLER_130_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07915_ _07924_/D _07914_/Y _08022_/B vssd1 vssd1 vccd1 vccd1 _07915_/Y sky130_fd_sc_hd__o21ai_1
X_08895_ _09234_/S1 _08893_/X _08894_/X vssd1 vssd1 vccd1 vccd1 _08895_/X sky130_fd_sc_hd__a21o_1
XFILLER_64_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07846_ _14750_/Q _07830_/A _07845_/Y vssd1 vssd1 vccd1 vccd1 _13525_/D sky130_fd_sc_hd__o21a_1
XFILLER_68_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07777_ _07777_/A _07777_/B _07777_/C vssd1 vssd1 vccd1 vccd1 _07777_/Y sky130_fd_sc_hd__nand3_1
XFILLER_17_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06728_ _14498_/Q vssd1 vssd1 vccd1 vccd1 _06728_/Y sky130_fd_sc_hd__clkinv_2
X_09516_ _12573_/A _09516_/B _09516_/C vssd1 vssd1 vccd1 vccd1 _09516_/X sky130_fd_sc_hd__and3_1
XFILLER_52_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09447_ _15134_/Q _15102_/Q _15675_/Q _13409_/Q _09441_/S _09448_/S1 vssd1 vssd1
+ vccd1 vccd1 _09447_/X sky130_fd_sc_hd__mux4_1
XPHY_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06659_ _14597_/Q vssd1 vssd1 vccd1 vccd1 _08754_/A sky130_fd_sc_hd__inv_2
XPHY_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_172_clk clkbuf_5_23_0_clk/X vssd1 vssd1 vccd1 vccd1 _14485_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_80_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09378_ _08494_/B _09376_/X _09377_/X vssd1 vssd1 vccd1 vccd1 _09382_/B sky130_fd_sc_hd__a21o_1
XFILLER_185_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08329_ _08305_/X _08328_/X _11088_/S vssd1 vssd1 vccd1 vccd1 _08329_/X sky130_fd_sc_hd__mux2_1
XFILLER_137_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11340_ _15040_/Q _08232_/A _08369_/X _11303_/Y _11339_/X vssd1 vssd1 vccd1 vccd1
+ _15040_/D sky130_fd_sc_hd__a221o_1
XFILLER_126_829 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11271_ _15030_/Q wire438/X _11269_/X _11270_/X vssd1 vssd1 vccd1 vccd1 _15030_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_152_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13010_ _15483_/Q _10892_/B _13116_/C _13009_/X vssd1 vssd1 vccd1 vccd1 _15483_/D
+ sky130_fd_sc_hd__a22o_1
X_10222_ input17/X _13125_/B _13309_/A vssd1 vssd1 vccd1 vccd1 _14607_/D sky130_fd_sc_hd__mux2_1
XFILLER_134_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10153_ _14538_/Q _13339_/A0 _10164_/S vssd1 vssd1 vccd1 vccd1 _14538_/D sky130_fd_sc_hd__mux2_1
XFILLER_95_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_1100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10084_ _14440_/Q _11870_/A1 _10097_/S vssd1 vssd1 vccd1 vccd1 _14440_/D sky130_fd_sc_hd__mux2_1
X_14961_ _15584_/CLK _14961_/D vssd1 vssd1 vccd1 vccd1 _14961_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_835 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold8 hold8/A vssd1 vssd1 vccd1 vccd1 hold8/X sky130_fd_sc_hd__bufbuf_16
X_13912_ _15499_/CLK _13912_/D vssd1 vssd1 vccd1 vccd1 _13912_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14892_ _14892_/CLK _14892_/D vssd1 vssd1 vccd1 vccd1 _14892_/Q sky130_fd_sc_hd__dfxtp_1
X_13843_ _15273_/CLK _13843_/D vssd1 vssd1 vccd1 vccd1 _13843_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13774_ _15462_/CLK _13774_/D vssd1 vssd1 vccd1 vccd1 _13774_/Q sky130_fd_sc_hd__dfxtp_2
X_10986_ _10986_/A _10986_/B vssd1 vssd1 vccd1 vccd1 _10987_/B sky130_fd_sc_hd__nor2_1
X_15513_ _15527_/CLK _15513_/D vssd1 vssd1 vccd1 vccd1 _15513_/Q sky130_fd_sc_hd__dfxtp_1
X_12725_ _12732_/B _12725_/B vssd1 vssd1 vccd1 vccd1 _12725_/Y sky130_fd_sc_hd__nor2_1
XFILLER_16_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_163_clk clkbuf_5_22_0_clk/X vssd1 vssd1 vccd1 vccd1 _15125_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_188_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15444_ _15630_/CLK _15444_/D vssd1 vssd1 vccd1 vccd1 _15444_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12656_ _15342_/Q _12759_/B _12655_/X _12832_/C1 vssd1 vssd1 vccd1 vccd1 _15342_/D
+ sky130_fd_sc_hd__o211a_1
X_11607_ _11614_/S _11611_/B _11606_/X vssd1 vssd1 vccd1 vccd1 _11607_/X sky130_fd_sc_hd__or3b_1
X_15375_ _15375_/CLK _15375_/D vssd1 vssd1 vccd1 vccd1 _15375_/Q sky130_fd_sc_hd__dfxtp_2
X_12587_ _13905_/Q _14420_/Q _12591_/S vssd1 vssd1 vccd1 vccd1 _12587_/X sky130_fd_sc_hd__mux2_1
XFILLER_12_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_156_464 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14326_ _15211_/CLK _14326_/D vssd1 vssd1 vccd1 vccd1 _14326_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11538_ _13236_/A _11569_/D vssd1 vssd1 vccd1 vccd1 _11539_/B sky130_fd_sc_hd__nor2_1
XFILLER_144_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_474 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11469_ _13195_/B _11470_/B vssd1 vssd1 vccd1 vccd1 _11471_/A sky130_fd_sc_hd__nor2_1
XFILLER_7_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14257_ _15335_/CLK _14257_/D vssd1 vssd1 vccd1 vccd1 _14257_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13208_ _13229_/A _13208_/B vssd1 vssd1 vccd1 vccd1 _13208_/Y sky130_fd_sc_hd__nor2_1
XFILLER_143_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14188_ _15674_/CLK _14188_/D vssd1 vssd1 vccd1 vccd1 _14188_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13139_ _14595_/Q _15536_/Q _13139_/S vssd1 vssd1 vccd1 vccd1 _15536_/D sky130_fd_sc_hd__mux2_1
XFILLER_98_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07700_ _13487_/Q _07697_/B _13488_/Q vssd1 vssd1 vccd1 vccd1 _07700_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_78_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08680_ _15378_/Q _08690_/A2 _08678_/X _08679_/X vssd1 vssd1 vccd1 vccd1 _08681_/C
+ sky130_fd_sc_hd__a211o_1
X_07631_ _13469_/Q _07655_/A _13470_/Q vssd1 vssd1 vccd1 vccd1 _07631_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_81_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07562_ _14740_/Q _07651_/A _07561_/Y _07938_/C1 vssd1 vssd1 vccd1 vccd1 _13451_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09301_ _09524_/A _09294_/X _09297_/X _08501_/A vssd1 vssd1 vccd1 vccd1 _09301_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_181_1023 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07493_ _13348_/A0 _13412_/Q _07501_/S vssd1 vssd1 vccd1 vccd1 _13412_/D sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_154_clk clkbuf_5_24_0_clk/X vssd1 vssd1 vccd1 vccd1 _15540_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_22_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09232_ _09234_/S1 _09230_/X _09231_/X vssd1 vssd1 vccd1 vccd1 _09232_/X sky130_fd_sc_hd__a21o_1
XFILLER_22_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09163_ _14467_/Q _14435_/Q _13856_/Q _14209_/Q _09444_/S _09448_/S1 vssd1 vssd1
+ vccd1 vccd1 _09163_/X sky130_fd_sc_hd__mux4_1
XFILLER_147_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08114_ input29/X input6/X input15/X input24/X _08150_/S _08151_/S vssd1 vssd1 vccd1
+ vccd1 _08114_/X sky130_fd_sc_hd__mux4_1
XFILLER_174_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09094_ _09449_/A1 _09092_/X _09093_/X _09449_/B2 vssd1 vssd1 vccd1 vccd1 _09094_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_119_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_637 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08045_ _14738_/Q _13616_/Q _08072_/S vssd1 vssd1 vccd1 vccd1 _13616_/D sky130_fd_sc_hd__mux2_1
XFILLER_102_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09996_ _13350_/A0 _14355_/Q _09996_/S vssd1 vssd1 vccd1 vccd1 _14355_/D sky130_fd_sc_hd__mux2_1
X_08947_ _15078_/Q _08540_/B _08946_/X _08501_/A vssd1 vssd1 vccd1 vccd1 _08947_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_3804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08878_ _13899_/Q _13343_/A0 _08880_/S vssd1 vssd1 vccd1 vccd1 _13899_/D sky130_fd_sc_hd__mux2_1
XFILLER_84_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07829_ _13521_/Q _07836_/D vssd1 vssd1 vccd1 vccd1 _07830_/B sky130_fd_sc_hd__xnor2_1
XTAP_3848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10840_ _14872_/Q _13796_/Q _12927_/S vssd1 vssd1 vccd1 vccd1 _14872_/D sky130_fd_sc_hd__mux2_1
XFILLER_44_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10771_ _14803_/Q _15435_/Q _12932_/S vssd1 vssd1 vccd1 vccd1 _14803_/D sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_145_clk clkbuf_5_28_0_clk/X vssd1 vssd1 vccd1 vccd1 _14493_/CLK sky130_fd_sc_hd__clkbuf_16
X_12510_ _12506_/X _12507_/X _12617_/S vssd1 vssd1 vccd1 vccd1 _12510_/X sky130_fd_sc_hd__mux2_1
X_13490_ _15383_/CLK _13490_/D vssd1 vssd1 vccd1 vccd1 _13490_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_9_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_537 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12441_ _12437_/X _12438_/X _12502_/S vssd1 vssd1 vccd1 vccd1 _12441_/X sky130_fd_sc_hd__mux2_1
XFILLER_40_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15160_ _15292_/CLK _15160_/D vssd1 vssd1 vccd1 vccd1 _15160_/Q sky130_fd_sc_hd__dfxtp_1
X_12372_ _12368_/X _12369_/X _12617_/S vssd1 vssd1 vccd1 vccd1 _12372_/X sky130_fd_sc_hd__mux2_1
XFILLER_154_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_934 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14111_ _14530_/CLK _14111_/D vssd1 vssd1 vccd1 vccd1 _14111_/Q sky130_fd_sc_hd__dfxtp_1
X_11323_ _11347_/A _11323_/B vssd1 vssd1 vccd1 vccd1 _11323_/Y sky130_fd_sc_hd__nand2_1
Xclkbuf_4_0_0_clk clkbuf_4_1_0_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_5_1_0_clk/A sky130_fd_sc_hd__clkbuf_8
X_15091_ _15664_/CLK _15091_/D vssd1 vssd1 vccd1 vccd1 _15091_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_153_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_467 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14042_ _14525_/CLK _14042_/D vssd1 vssd1 vccd1 vccd1 _14042_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_107_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11254_ _11283_/A _11311_/B vssd1 vssd1 vccd1 vccd1 _11254_/Y sky130_fd_sc_hd__nand2_1
XFILLER_4_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10205_ input30/X hold5/A _13284_/S vssd1 vssd1 vccd1 vccd1 _14590_/D sky130_fd_sc_hd__mux2_1
XFILLER_106_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11185_ _11380_/A _11185_/B vssd1 vssd1 vccd1 vccd1 _11185_/Y sky130_fd_sc_hd__nor2_1
XFILLER_133_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10136_ _14521_/Q _11680_/A0 _10159_/S vssd1 vssd1 vccd1 vccd1 _14521_/D sky130_fd_sc_hd__mux2_1
XFILLER_79_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_632 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14944_ _15020_/CLK _14944_/D vssd1 vssd1 vccd1 vccd1 _14944_/Q sky130_fd_sc_hd__dfxtp_1
X_10067_ _14423_/Q _13320_/A0 _10097_/S vssd1 vssd1 vccd1 vccd1 _14423_/D sky130_fd_sc_hd__mux2_1
XFILLER_91_911 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14875_ _15596_/CLK _14875_/D vssd1 vssd1 vccd1 vccd1 _14875_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_36_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13826_ _15306_/CLK _13826_/D vssd1 vssd1 vccd1 vccd1 _13826_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13757_ _14888_/CLK _13757_/D vssd1 vssd1 vccd1 vccd1 _13757_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_136_clk clkbuf_5_29_0_clk/X vssd1 vssd1 vccd1 vccd1 _13642_/CLK sky130_fd_sc_hd__clkbuf_16
X_10969_ _11037_/A _13208_/B vssd1 vssd1 vccd1 vccd1 _11258_/B sky130_fd_sc_hd__and2_1
XFILLER_43_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12708_ _15349_/Q _12765_/B _12707_/X _12809_/C1 vssd1 vssd1 vccd1 vccd1 _15349_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_149_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13688_ _15276_/CLK _13688_/D vssd1 vssd1 vccd1 vccd1 _13688_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_1070 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15427_ _15612_/CLK _15427_/D vssd1 vssd1 vccd1 vccd1 _15427_/Q sky130_fd_sc_hd__dfxtp_1
X_12639_ _13584_/Q _12638_/X _12785_/B vssd1 vssd1 vccd1 vccd1 _12639_/X sky130_fd_sc_hd__mux2_1
XFILLER_15_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15358_ _15638_/CLK _15358_/D vssd1 vssd1 vccd1 vccd1 _15358_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_117_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14309_ _15125_/CLK _14309_/D vssd1 vssd1 vccd1 vccd1 _14309_/Q sky130_fd_sc_hd__dfxtp_1
X_15289_ _15289_/CLK _15289_/D vssd1 vssd1 vccd1 vccd1 _15289_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_1079 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09850_ _14214_/Q _11870_/A1 _09863_/S vssd1 vssd1 vccd1 vccd1 _14214_/D sky130_fd_sc_hd__mux2_1
XTAP_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08801_ _11868_/A1 _13827_/Q _08811_/S vssd1 vssd1 vccd1 vccd1 _13827_/D sky130_fd_sc_hd__mux2_1
XTAP_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09781_ _14148_/Q _13086_/B2 _09795_/S vssd1 vssd1 vccd1 vccd1 _14148_/D sky130_fd_sc_hd__mux2_1
XFILLER_86_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06993_ _14923_/Q _10344_/S _06861_/Y _12832_/C1 _06782_/A vssd1 vssd1 vccd1 vccd1
+ _14730_/D sky130_fd_sc_hd__o2111a_1
XTAP_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08732_ _13803_/Q _12932_/S _08726_/X _08731_/X vssd1 vssd1 vccd1 vccd1 _13803_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_82_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08663_ _15380_/Q _08690_/A2 _08690_/B1 _13425_/Q vssd1 vssd1 vccd1 vccd1 _08663_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_82_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07614_ _07614_/A _07614_/B vssd1 vssd1 vccd1 vccd1 _07614_/Y sky130_fd_sc_hd__nand2_1
X_08594_ _13531_/Q _08683_/A2 _08691_/B1 _13499_/Q _08593_/X vssd1 vssd1 vccd1 vccd1
+ _08598_/B sky130_fd_sc_hd__a221o_1
XTAP_1709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07545_ _13446_/Q _13445_/Q _13447_/Q vssd1 vssd1 vccd1 vccd1 _07545_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_179_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_127_clk clkbuf_5_31_0_clk/X vssd1 vssd1 vccd1 vccd1 _13565_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_35_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07476_ _14759_/Q _07475_/X _07480_/S vssd1 vssd1 vccd1 vccd1 _07476_/X sky130_fd_sc_hd__mux2_8
X_09215_ _15664_/Q _13398_/Q _09441_/S vssd1 vssd1 vccd1 vccd1 _09215_/X sky130_fd_sc_hd__mux2_1
XFILLER_10_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09146_ _09421_/A1 _09142_/X _09145_/X _09141_/X vssd1 vssd1 vccd1 vccd1 _09146_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_108_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09077_ _12596_/A _09077_/B _09077_/C vssd1 vssd1 vccd1 vccd1 _09077_/X sky130_fd_sc_hd__and3_2
XFILLER_162_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08028_ _08028_/A _08028_/B vssd1 vssd1 vccd1 vccd1 _08028_/X sky130_fd_sc_hd__or2_1
XFILLER_162_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_1091 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09979_ _13080_/B2 _14338_/Q _09991_/S vssd1 vssd1 vccd1 vccd1 _14338_/D sky130_fd_sc_hd__mux2_1
XFILLER_58_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12990_ _10654_/X _14877_/Q _13029_/S vssd1 vssd1 vccd1 vccd1 _12990_/X sky130_fd_sc_hd__mux2_4
XFILLER_183_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11941_ _13941_/Q _13683_/Q _12543_/S vssd1 vssd1 vccd1 vccd1 _11942_/B sky130_fd_sc_hd__mux2_1
XFILLER_85_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_635 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14660_ _15446_/CLK _14660_/D vssd1 vssd1 vccd1 vccd1 _14660_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11872_ _15293_/Q _11872_/A1 _11883_/S vssd1 vssd1 vccd1 vccd1 _15293_/D sky130_fd_sc_hd__mux2_1
XFILLER_44_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13611_ _15461_/CLK _13611_/D vssd1 vssd1 vccd1 vccd1 _13611_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10823_ _14855_/Q _07206_/X _10868_/S vssd1 vssd1 vccd1 vccd1 _14855_/D sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_118_clk clkbuf_5_30_0_clk/X vssd1 vssd1 vccd1 vccd1 _15377_/CLK sky130_fd_sc_hd__clkbuf_16
X_14591_ _15530_/CLK _14591_/D vssd1 vssd1 vccd1 vccd1 _14591_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_2988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_532 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13542_ _15542_/CLK _13542_/D vssd1 vssd1 vccd1 vccd1 _13542_/Q sky130_fd_sc_hd__dfxtp_2
X_10754_ _15418_/Q _14786_/Q _10765_/S vssd1 vssd1 vccd1 vccd1 _14786_/D sky130_fd_sc_hd__mux2_1
XFILLER_158_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_536 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10685_ _14755_/Q _10684_/X _10715_/S vssd1 vssd1 vccd1 vccd1 _14755_/D sky130_fd_sc_hd__mux2_1
XFILLER_139_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13473_ _15398_/CLK _13473_/D vssd1 vssd1 vccd1 vccd1 _13473_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_139_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15212_ _15212_/CLK _15212_/D vssd1 vssd1 vccd1 vccd1 _15212_/Q sky130_fd_sc_hd__dfxtp_1
X_12424_ _13962_/Q _13704_/Q _12430_/S vssd1 vssd1 vccd1 vccd1 _12425_/B sky130_fd_sc_hd__mux2_1
X_15143_ _15212_/CLK _15143_/D vssd1 vssd1 vccd1 vccd1 _15143_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_126_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12355_ _13959_/Q _13701_/Q _12541_/S vssd1 vssd1 vccd1 vccd1 _12356_/B sky130_fd_sc_hd__mux2_1
XFILLER_4_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11306_ _11318_/S _11304_/Y _11305_/X vssd1 vssd1 vccd1 vccd1 _11307_/B sky130_fd_sc_hd__a21oi_1
X_12286_ _13956_/Q _13698_/Q _12614_/S vssd1 vssd1 vccd1 vccd1 _12287_/B sky130_fd_sc_hd__mux2_1
X_15074_ _15613_/CLK _15074_/D vssd1 vssd1 vccd1 vccd1 _15074_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_141_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14025_ _15654_/CLK _14025_/D vssd1 vssd1 vccd1 vccd1 _14025_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11237_ _11639_/A _15025_/Q _11237_/S vssd1 vssd1 vccd1 vccd1 _15025_/D sky130_fd_sc_hd__mux2_1
XFILLER_110_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11168_ _11414_/A _11165_/X _11167_/Y vssd1 vssd1 vccd1 vccd1 _11168_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_96_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10119_ _14505_/Q _14753_/Q _10131_/S vssd1 vssd1 vccd1 vccd1 _14505_/D sky130_fd_sc_hd__mux2_1
XFILLER_121_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11099_ _10988_/Y _11047_/Y _11344_/A vssd1 vssd1 vccd1 vccd1 _11099_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_49_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14927_ _15613_/CLK _14927_/D vssd1 vssd1 vccd1 vccd1 _14927_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_35_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14858_ _15500_/CLK _14858_/D vssd1 vssd1 vccd1 vccd1 _14858_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13809_ _15208_/CLK _13809_/D vssd1 vssd1 vccd1 vccd1 _13809_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_109_clk clkbuf_5_26_0_clk/X vssd1 vssd1 vccd1 vccd1 _15634_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_17_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14789_ _15641_/CLK _14789_/D vssd1 vssd1 vccd1 vccd1 _14789_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07330_ _13907_/Q _15494_/Q _07339_/S vssd1 vssd1 vccd1 vccd1 _07331_/A sky130_fd_sc_hd__mux2_4
XFILLER_177_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07261_ _07261_/A _07261_/B vssd1 vssd1 vccd1 vccd1 _07270_/C sky130_fd_sc_hd__nor2_1
XFILLER_149_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09000_ _14459_/Q _09558_/A2 _08999_/X _13049_/A1 vssd1 vssd1 vccd1 vccd1 _09000_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_118_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_3_7_0_clk clkbuf_3_7_0_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_7_0_clk/X sky130_fd_sc_hd__clkbuf_8
X_07192_ _15366_/Q _15073_/Q _07193_/S vssd1 vssd1 vccd1 vccd1 _07192_/X sky130_fd_sc_hd__mux2_8
XFILLER_117_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_968 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09902_ _13322_/A0 _14263_/Q _09925_/S vssd1 vssd1 vccd1 vccd1 _14263_/D sky130_fd_sc_hd__mux2_1
XFILLER_99_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout504 _07096_/S vssd1 vssd1 vccd1 vccd1 _07078_/S sky130_fd_sc_hd__buf_12
Xfanout515 _14606_/Q vssd1 vssd1 vccd1 vccd1 _09405_/A sky130_fd_sc_hd__buf_12
XFILLER_113_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout526 _08988_/A1 vssd1 vssd1 vccd1 vccd1 _09429_/S1 sky130_fd_sc_hd__buf_12
XFILLER_98_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout537 _09553_/A1 vssd1 vssd1 vccd1 vccd1 _08519_/A sky130_fd_sc_hd__buf_12
X_09833_ _14197_/Q _13320_/A0 _09863_/S vssd1 vssd1 vccd1 vccd1 _14197_/D sky130_fd_sc_hd__mux2_1
XFILLER_113_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout548 _09047_/S vssd1 vssd1 vccd1 vccd1 _09230_/S sky130_fd_sc_hd__buf_12
XFILLER_113_684 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout559 _09551_/S vssd1 vssd1 vccd1 vccd1 _09484_/S sky130_fd_sc_hd__buf_12
XTAP_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09764_ _14131_/Q _13319_/A0 _09790_/S vssd1 vssd1 vccd1 vccd1 _14131_/D sky130_fd_sc_hd__mux2_1
XTAP_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06976_ _06969_/D _06976_/B vssd1 vssd1 vccd1 vccd1 _06977_/B sky130_fd_sc_hd__and2b_1
X_08715_ _14491_/Q _08748_/B1 _08712_/X _08713_/X _08714_/X vssd1 vssd1 vccd1 vccd1
+ _08715_/X sky130_fd_sc_hd__a2111o_2
XFILLER_6_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09695_ _14066_/Q _11883_/A1 _09695_/S vssd1 vssd1 vccd1 vccd1 _14066_/D sky130_fd_sc_hd__mux2_1
XFILLER_66_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08646_ _13791_/Q _12917_/S _08645_/X vssd1 vssd1 vccd1 vccd1 _13791_/D sky130_fd_sc_hd__o21a_1
XFILLER_148_1024 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_262 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08577_ _13502_/Q _08747_/B1 _08693_/B1 _13637_/Q vssd1 vssd1 vccd1 vccd1 _08577_/X
+ sky130_fd_sc_hd__a22o_1
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_186_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_148 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07528_ _14758_/Q _13437_/Q _07529_/S vssd1 vssd1 vccd1 vccd1 _13437_/D sky130_fd_sc_hd__mux2_1
XFILLER_179_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_502 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07459_ _13670_/Q _07483_/A2 _07483_/B1 _14698_/Q _07458_/X vssd1 vssd1 vccd1 vccd1
+ _07459_/X sky130_fd_sc_hd__a221o_1
XFILLER_41_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10470_ _10470_/A _10470_/B _10470_/C _10470_/D vssd1 vssd1 vccd1 vccd1 _10471_/D
+ sky130_fd_sc_hd__or4_1
X_09129_ _09234_/S1 _09127_/X _09128_/X vssd1 vssd1 vccd1 vccd1 _09130_/C sky130_fd_sc_hd__a21o_1
XFILLER_108_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12140_ _14529_/Q _14142_/Q _14174_/Q _14110_/Q _11993_/S _12253_/S1 vssd1 vssd1
+ vccd1 vccd1 _12140_/X sky130_fd_sc_hd__mux4_1
XFILLER_2_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12071_ _14526_/Q _14139_/Q _14171_/Q _14107_/Q _12079_/S _12268_/A vssd1 vssd1 vccd1
+ vccd1 _12071_/X sky130_fd_sc_hd__mux4_1
XFILLER_173_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11022_ _11037_/A _11584_/A vssd1 vssd1 vccd1 vccd1 _11312_/B sky130_fd_sc_hd__nand2_1
XFILLER_131_470 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12973_ _13328_/A0 _13024_/A2 _12972_/X _13024_/B2 vssd1 vssd1 vccd1 vccd1 _12973_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_3431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14712_ _15489_/CLK _14712_/D vssd1 vssd1 vccd1 vccd1 _14712_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_3464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11924_ _14068_/Q _14036_/Q _12614_/S vssd1 vssd1 vccd1 vccd1 _11924_/X sky130_fd_sc_hd__mux2_1
XTAP_3475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14643_ _14649_/CLK _14643_/D vssd1 vssd1 vccd1 vccd1 _14643_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11855_ _15276_/Q _13322_/A0 _11878_/S vssd1 vssd1 vccd1 vccd1 _15276_/D sky130_fd_sc_hd__mux2_1
XTAP_2774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10806_ _14838_/Q _07306_/A _12481_/A vssd1 vssd1 vccd1 vccd1 _14838_/D sky130_fd_sc_hd__mux2_1
XFILLER_82_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14574_ _15652_/CLK _14574_/D vssd1 vssd1 vccd1 vccd1 _14574_/Q sky130_fd_sc_hd__dfxtp_1
X_11786_ _15209_/Q _11852_/A1 _11816_/S vssd1 vssd1 vccd1 vccd1 _15209_/D sky130_fd_sc_hd__mux2_1
XFILLER_186_632 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13525_ _13627_/CLK _13525_/D vssd1 vssd1 vccd1 vccd1 _13525_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10737_ _15401_/Q _14769_/Q _13129_/A vssd1 vssd1 vccd1 vccd1 _14769_/D sky130_fd_sc_hd__mux2_1
XFILLER_158_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_170 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13456_ _15379_/CLK _13456_/D vssd1 vssd1 vccd1 vccd1 _13456_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_158_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10668_ _14980_/Q _10718_/A2 _10722_/B1 _14948_/Q _10667_/X vssd1 vssd1 vccd1 vccd1
+ _10668_/X sky130_fd_sc_hd__a221o_1
XFILLER_9_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12407_ _14089_/Q _14057_/Q _12407_/S vssd1 vssd1 vccd1 vccd1 _12407_/X sky130_fd_sc_hd__mux2_1
XFILLER_154_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13387_ _15660_/CLK _13387_/D vssd1 vssd1 vccd1 vccd1 _13387_/Q sky130_fd_sc_hd__dfxtp_1
X_10599_ _15047_/Q _10734_/A2 _10596_/X _10598_/X vssd1 vssd1 vccd1 vccd1 _10599_/X
+ sky130_fd_sc_hd__o22a_2
XFILLER_126_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15126_ _15667_/CLK _15126_/D vssd1 vssd1 vccd1 vccd1 _15126_/Q sky130_fd_sc_hd__dfxtp_1
X_12338_ _14086_/Q _14054_/Q _12543_/S vssd1 vssd1 vccd1 vccd1 _12338_/X sky130_fd_sc_hd__mux2_1
XFILLER_5_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15057_ _15599_/CLK _15057_/D vssd1 vssd1 vccd1 vccd1 _15057_/Q sky130_fd_sc_hd__dfxtp_4
X_12269_ _14083_/Q _14051_/Q _12269_/S vssd1 vssd1 vccd1 vccd1 _12269_/X sky130_fd_sc_hd__mux2_1
XFILLER_141_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14008_ _15278_/CLK _14008_/D vssd1 vssd1 vccd1 vccd1 _14008_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06830_ _15540_/Q _13737_/Q _14896_/Q _14923_/Q _08036_/A vssd1 vssd1 vccd1 vccd1
+ _06830_/X sky130_fd_sc_hd__a221o_1
XFILLER_83_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06761_ input19/X vssd1 vssd1 vccd1 vccd1 _06761_/Y sky130_fd_sc_hd__inv_2
XFILLER_83_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08500_ _14608_/Q _14610_/Q vssd1 vssd1 vccd1 vccd1 _08536_/B sky130_fd_sc_hd__nand2b_1
X_09480_ _08510_/B _09478_/X _09479_/X _08519_/B _13049_/A1 vssd1 vssd1 vccd1 vccd1
+ _09480_/X sky130_fd_sc_hd__a221o_1
X_06692_ _14515_/Q vssd1 vssd1 vccd1 vccd1 _06692_/Y sky130_fd_sc_hd__inv_2
XFILLER_24_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08431_ _14611_/Q _08390_/C _08425_/X _10764_/S vssd1 vssd1 vccd1 vccd1 _08431_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_24_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08362_ _08244_/A _13761_/Q _15411_/Q _08244_/B vssd1 vssd1 vccd1 vccd1 _08362_/X
+ sky130_fd_sc_hd__a22o_2
XFILLER_20_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07313_ _15312_/Q _15468_/Q _07335_/S vssd1 vssd1 vccd1 vccd1 _07314_/A sky130_fd_sc_hd__mux2_8
XFILLER_149_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_833 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08293_ _11349_/B _13171_/B vssd1 vssd1 vccd1 vccd1 _10999_/B sky130_fd_sc_hd__and2_1
XFILLER_177_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07244_ _07244_/A vssd1 vssd1 vccd1 vccd1 _07244_/Y sky130_fd_sc_hd__inv_2
XFILLER_176_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07175_ _15349_/Q _15056_/Q _07193_/S vssd1 vssd1 vccd1 vccd1 _07175_/X sky130_fd_sc_hd__mux2_1
XFILLER_145_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_37 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout301 _07464_/X vssd1 vssd1 vccd1 vccd1 _11874_/A1 sky130_fd_sc_hd__buf_6
Xfanout312 _13086_/B2 vssd1 vssd1 vccd1 vccd1 _11761_/A0 sky130_fd_sc_hd__buf_6
XFILLER_132_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout323 _07424_/X vssd1 vssd1 vccd1 vccd1 _13331_/A0 sky130_fd_sc_hd__buf_6
Xfanout334 _07404_/X vssd1 vssd1 vccd1 vccd1 _12967_/A1 sky130_fd_sc_hd__clkbuf_16
XFILLER_114_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout345 _07384_/X vssd1 vssd1 vccd1 vccd1 _13321_/A0 sky130_fd_sc_hd__buf_4
XFILLER_115_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout356 _10734_/A2 vssd1 vssd1 vccd1 vccd1 _10714_/A2 sky130_fd_sc_hd__buf_12
XFILLER_28_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09816_ _14182_/Q _13338_/A0 _09828_/S vssd1 vssd1 vccd1 vccd1 _14182_/D sky130_fd_sc_hd__mux2_1
Xfanout367 _09421_/A1 vssd1 vssd1 vccd1 vccd1 _09449_/B2 sky130_fd_sc_hd__buf_12
XFILLER_86_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout378 _11356_/B vssd1 vssd1 vccd1 vccd1 _11330_/A sky130_fd_sc_hd__buf_8
Xfanout389 _08231_/X vssd1 vssd1 vccd1 vccd1 _11344_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_86_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09747_ _14115_/Q _13335_/A0 _09757_/S vssd1 vssd1 vccd1 vccd1 _14115_/D sky130_fd_sc_hd__mux2_1
XFILLER_100_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06959_ _06750_/Y _13479_/Q _06753_/Y _13478_/Q _06948_/X vssd1 vssd1 vccd1 vccd1
+ _06960_/B sky130_fd_sc_hd__o221a_1
XFILLER_39_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09678_ _14049_/Q _13333_/A0 _09690_/S vssd1 vssd1 vccd1 vccd1 _14049_/D sky130_fd_sc_hd__mux2_1
XFILLER_54_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08629_ _15385_/Q _08690_/A2 _08736_/A2 _13430_/Q vssd1 vssd1 vccd1 vccd1 _08629_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_1325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11640_ _11640_/A _11640_/B vssd1 vssd1 vccd1 vccd1 _11640_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_30_619 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11571_ _11589_/B _11571_/B vssd1 vssd1 vccd1 vccd1 _11572_/B sky130_fd_sc_hd__xnor2_4
XFILLER_22_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13310_ _15641_/Q _13309_/A _13309_/X vssd1 vssd1 vccd1 vccd1 _15641_/D sky130_fd_sc_hd__a21bo_1
XFILLER_156_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10522_ _08244_/A _13755_/Q _15417_/Q _08244_/B vssd1 vssd1 vccd1 vccd1 _10522_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_168_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14290_ _14542_/CLK _14290_/D vssd1 vssd1 vccd1 vccd1 _14290_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13241_ _15580_/Q _13241_/A2 _13239_/X _13240_/Y vssd1 vssd1 vccd1 vccd1 _15580_/D
+ sky130_fd_sc_hd__a22o_1
X_10453_ _11582_/A _11584_/A vssd1 vssd1 vccd1 vccd1 _10455_/A sky130_fd_sc_hd__or2_1
XFILLER_170_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10384_ _10384_/A vssd1 vssd1 vccd1 vccd1 _10390_/B sky130_fd_sc_hd__inv_2
X_13172_ _13251_/A _13171_/B _11414_/D _13252_/B vssd1 vssd1 vccd1 vccd1 _13172_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_108_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12123_ _08453_/A _12120_/X _08451_/A vssd1 vssd1 vccd1 vccd1 _12123_/X sky130_fd_sc_hd__o21a_1
XFILLER_124_779 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12054_ _12500_/B1 _12051_/X _12501_/C1 vssd1 vssd1 vccd1 vccd1 _12054_/X sky130_fd_sc_hd__o21a_1
XFILLER_77_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11005_ _11013_/A _13242_/B vssd1 vssd1 vccd1 vccd1 _11007_/B sky130_fd_sc_hd__nand2_1
XFILLER_81_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12956_ _15465_/Q _13081_/A2 _13025_/B1 _12955_/X vssd1 vssd1 vccd1 vccd1 _15465_/D
+ sky130_fd_sc_hd__a22o_1
XTAP_3261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11907_ _15306_/Q _13105_/A2 _11906_/X vssd1 vssd1 vccd1 vccd1 _15306_/D sky130_fd_sc_hd__a21o_1
X_15675_ _15675_/CLK _15675_/D vssd1 vssd1 vccd1 vccd1 _15675_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12887_ _15415_/Q _15600_/Q _12928_/S vssd1 vssd1 vccd1 vccd1 _15415_/D sky130_fd_sc_hd__mux2_1
XTAP_2571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14626_ _15596_/CLK _14626_/D vssd1 vssd1 vccd1 vccd1 _14626_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11838_ _15260_/Q _11838_/A1 _11850_/S vssd1 vssd1 vccd1 vccd1 _15260_/D sky130_fd_sc_hd__mux2_1
XTAP_1870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14557_ _15220_/CLK _14557_/D vssd1 vssd1 vccd1 vccd1 _14557_/Q sky130_fd_sc_hd__dfxtp_1
X_11769_ _11877_/A1 _15197_/Q _11774_/S vssd1 vssd1 vccd1 vccd1 _15197_/D sky130_fd_sc_hd__mux2_1
XFILLER_13_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_40_clk clkbuf_5_12_0_clk/X vssd1 vssd1 vccd1 vccd1 _15589_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_158_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13508_ _13642_/CLK _13508_/D vssd1 vssd1 vccd1 vccd1 _13508_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_147_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14488_ _15542_/CLK _14488_/D vssd1 vssd1 vccd1 vccd1 _14488_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_173_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13439_ _15375_/CLK _13439_/D vssd1 vssd1 vccd1 vccd1 _13439_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15109_ _15650_/CLK _15109_/D vssd1 vssd1 vccd1 vccd1 _15109_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08980_ _13879_/Q _09231_/A2 _09403_/B1 _14394_/Q _09445_/C1 vssd1 vssd1 vccd1 vccd1
+ _08980_/X sky130_fd_sc_hd__a221o_1
XFILLER_88_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07931_ _14740_/Q _08012_/A2 _07930_/X _07938_/C1 vssd1 vssd1 vccd1 vccd1 _13547_/D
+ sky130_fd_sc_hd__o211a_1
X_07862_ _13530_/Q _07869_/D vssd1 vssd1 vccd1 vccd1 _07866_/B sky130_fd_sc_hd__nand2_1
XFILLER_68_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_151 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09601_ _13975_/Q _11681_/A0 _09627_/S vssd1 vssd1 vccd1 vccd1 _13975_/D sky130_fd_sc_hd__mux2_1
X_06813_ _13732_/Q _08668_/B _09466_/A _06665_/Y _06811_/X vssd1 vssd1 vccd1 vccd1
+ _06813_/X sky130_fd_sc_hd__a221o_1
XFILLER_28_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07793_ _14736_/Q _07816_/A _07792_/Y _08084_/C1 vssd1 vssd1 vccd1 vccd1 _13511_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_3_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09532_ _09532_/A _09532_/B vssd1 vssd1 vccd1 vccd1 _09532_/X sky130_fd_sc_hd__or2_1
X_06744_ _13450_/Q vssd1 vssd1 vccd1 vccd1 _06744_/Y sky130_fd_sc_hd__inv_2
XFILLER_83_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06675_ _09532_/A vssd1 vssd1 vccd1 vccd1 _06675_/Y sky130_fd_sc_hd__clkinv_8
X_09463_ _09382_/A _09456_/X _09459_/X _09462_/X vssd1 vssd1 vccd1 vccd1 _09463_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_36_295 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08414_ _14596_/Q _14595_/Q _08777_/A _08413_/X vssd1 vssd1 vccd1 vccd1 _13739_/D
+ sky130_fd_sc_hd__a31o_1
X_09394_ _14252_/Q _14284_/Q _14316_/Q _14348_/Q _09407_/S _09406_/S1 vssd1 vssd1
+ vccd1 vccd1 _09394_/X sky130_fd_sc_hd__mux4_1
X_08345_ _11037_/A _11449_/A vssd1 vssd1 vccd1 vccd1 _11034_/A sky130_fd_sc_hd__nor2_1
XFILLER_138_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_31_clk clkbuf_5_7_0_clk/X vssd1 vssd1 vccd1 vccd1 _15519_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_137_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08276_ _10507_/A1 _13770_/Q _15402_/Q _10515_/B2 vssd1 vssd1 vccd1 vccd1 _08276_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_137_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07227_ _07227_/A _07227_/B vssd1 vssd1 vccd1 vccd1 _07227_/Y sky130_fd_sc_hd__nor2_1
XFILLER_138_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07158_ _14859_/Q _14851_/Q _14843_/Q _14835_/Q _08150_/S _08151_/S vssd1 vssd1 vccd1
+ vccd1 _07159_/B sky130_fd_sc_hd__mux4_1
XFILLER_3_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07089_ _07088_/X _14762_/Q _07098_/S vssd1 vssd1 vccd1 vccd1 _13608_/D sky130_fd_sc_hd__mux2_1
XFILLER_161_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout120 _13051_/X vssd1 vssd1 vccd1 vccd1 _13114_/B1 sky130_fd_sc_hd__buf_8
Xfanout131 fanout138/X vssd1 vssd1 vccd1 vccd1 _13093_/A2 sky130_fd_sc_hd__buf_8
Xclkbuf_leaf_98_clk clkbuf_5_25_0_clk/X vssd1 vssd1 vccd1 vccd1 _15647_/CLK sky130_fd_sc_hd__clkbuf_16
Xfanout142 _10871_/S vssd1 vssd1 vccd1 vccd1 _13138_/S sky130_fd_sc_hd__clkbuf_16
Xfanout153 _12885_/S vssd1 vssd1 vccd1 vccd1 _12917_/S sky130_fd_sc_hd__buf_12
XFILLER_75_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout164 _13318_/X vssd1 vssd1 vccd1 vccd1 _13350_/S sky130_fd_sc_hd__buf_12
Xfanout175 _11710_/Y vssd1 vssd1 vccd1 vccd1 _11741_/S sky130_fd_sc_hd__buf_12
Xfanout186 _10065_/Y vssd1 vssd1 vccd1 vccd1 _10097_/S sky130_fd_sc_hd__buf_12
Xfanout197 _09865_/Y vssd1 vssd1 vccd1 vccd1 _09892_/S sky130_fd_sc_hd__buf_12
XFILLER_75_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12810_ _15364_/Q _15363_/Q _12810_/C vssd1 vssd1 vccd1 vccd1 _12819_/B sky130_fd_sc_hd__and3_1
X_13790_ _15596_/CLK _13790_/D vssd1 vssd1 vccd1 vccd1 _13790_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_16_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12741_ _13598_/Q _12740_/X _12785_/B vssd1 vssd1 vccd1 vccd1 _12741_/X sky130_fd_sc_hd__mux2_1
XTAP_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15460_ _15622_/CLK _15460_/D vssd1 vssd1 vccd1 vccd1 _15460_/Q sky130_fd_sc_hd__dfxtp_1
X_12672_ _15344_/Q _12759_/B _12671_/X _12832_/C1 vssd1 vssd1 vccd1 vccd1 _15344_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14411_ _15680_/CLK _14411_/D vssd1 vssd1 vccd1 vccd1 _14411_/Q sky130_fd_sc_hd__dfxtp_1
X_11623_ _13236_/A _11616_/A _11616_/B vssd1 vssd1 vccd1 vccd1 _11624_/B sky130_fd_sc_hd__o21a_1
XTAP_1199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15391_ _15393_/CLK _15391_/D vssd1 vssd1 vccd1 vccd1 _15391_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_184_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_22_clk clkbuf_5_3_0_clk/X vssd1 vssd1 vccd1 vccd1 _15331_/CLK sky130_fd_sc_hd__clkbuf_16
X_14342_ _15301_/CLK _14342_/D vssd1 vssd1 vccd1 vccd1 _14342_/Q sky130_fd_sc_hd__dfxtp_1
X_11554_ _11555_/A _11555_/B vssd1 vssd1 vccd1 vccd1 _11554_/X sky130_fd_sc_hd__and2_1
XFILLER_11_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10505_ _10520_/A1 _13786_/Q _13754_/Q _10520_/B2 vssd1 vssd1 vccd1 vccd1 _10505_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_128_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14273_ _15235_/CLK _14273_/D vssd1 vssd1 vccd1 vccd1 _14273_/Q sky130_fd_sc_hd__dfxtp_1
X_11485_ _11505_/C _11484_/B _11474_/S vssd1 vssd1 vccd1 vccd1 _11485_/X sky130_fd_sc_hd__o21ba_1
XFILLER_184_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13224_ _13236_/A _10544_/X _13214_/B _13223_/Y vssd1 vssd1 vccd1 vccd1 _13224_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_155_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10436_ _10520_/A1 _13777_/Q _13745_/Q _10520_/B2 vssd1 vssd1 vccd1 vccd1 _10436_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_124_543 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13155_ _14929_/D _14928_/D _14927_/D vssd1 vssd1 vccd1 vccd1 _13219_/S sky130_fd_sc_hd__and3_4
X_10367_ _10520_/A1 _13798_/Q _13766_/Q _10520_/B2 vssd1 vssd1 vccd1 vccd1 _10367_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_88_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_576 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12106_ _14012_/Q _13980_/Q _12476_/S vssd1 vssd1 vccd1 vccd1 _12107_/B sky130_fd_sc_hd__mux2_1
XFILLER_97_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13086_ _12996_/X _13118_/A2 _13114_/B1 _13086_/B2 vssd1 vssd1 vccd1 vccd1 _13086_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_97_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10298_ _14683_/Q _14868_/Q _10610_/S vssd1 vssd1 vccd1 vccd1 _14683_/D sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_89_clk clkbuf_5_13_0_clk/X vssd1 vssd1 vccd1 vccd1 _14649_/CLK sky130_fd_sc_hd__clkbuf_16
X_12037_ _14009_/Q _13977_/Q _12591_/S vssd1 vssd1 vccd1 vccd1 _12038_/B sky130_fd_sc_hd__mux2_1
XFILLER_168_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13988_ _15651_/CLK _13988_/D vssd1 vssd1 vccd1 vccd1 _13988_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_168_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12939_ _08405_/A _09662_/B _08852_/B _12563_/A vssd1 vssd1 vccd1 vccd1 _12943_/B
+ sky130_fd_sc_hd__o22ai_1
XTAP_3091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15658_ _15658_/CLK _15658_/D vssd1 vssd1 vccd1 vccd1 _15658_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14609_ _15648_/CLK _14609_/D vssd1 vssd1 vccd1 vccd1 _14609_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_21_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15589_ _15589_/CLK _15589_/D vssd1 vssd1 vccd1 vccd1 _15589_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_13_clk clkbuf_5_2_0_clk/X vssd1 vssd1 vccd1 vccd1 _15662_/CLK sky130_fd_sc_hd__clkbuf_16
X_08130_ _08145_/S _06761_/Y _08093_/B vssd1 vssd1 vccd1 vccd1 _08130_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_179_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08061_ _14754_/Q _13632_/Q _08066_/S vssd1 vssd1 vccd1 vccd1 _13632_/D sky130_fd_sc_hd__mux2_1
XFILLER_105_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07012_ _14616_/Q _14648_/Q _07096_/S vssd1 vssd1 vccd1 vccd1 _07012_/X sky130_fd_sc_hd__mux2_1
XFILLER_175_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08963_ _14006_/Q _13974_/Q _09073_/S vssd1 vssd1 vccd1 vccd1 _08963_/X sky130_fd_sc_hd__mux2_1
XFILLER_102_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07914_ _13542_/Q _13541_/Q _07913_/D _13543_/Q vssd1 vssd1 vccd1 vccd1 _07914_/Y
+ sky130_fd_sc_hd__a31oi_1
XFILLER_130_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08894_ _14067_/Q _09231_/A2 _09403_/B1 _14035_/Q _09221_/A vssd1 vssd1 vccd1 vccd1
+ _08894_/X sky130_fd_sc_hd__a221o_1
XFILLER_69_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_994 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07845_ _07783_/X _07844_/X input35/X vssd1 vssd1 vccd1 vccd1 _07845_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_151_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_346 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07776_ _13508_/Q _13507_/Q _07776_/C vssd1 vssd1 vccd1 vccd1 _07777_/C sky130_fd_sc_hd__nand3b_1
XFILLER_140_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09515_ _08668_/D _09511_/X _09514_/X _09510_/X vssd1 vssd1 vccd1 vccd1 _09516_/C
+ sky130_fd_sc_hd__a211o_1
X_06727_ _13458_/Q vssd1 vssd1 vccd1 vccd1 _06727_/Y sky130_fd_sc_hd__inv_2
XFILLER_140_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09446_ _09446_/A1 _09444_/X _09445_/X vssd1 vssd1 vccd1 vccd1 _09446_/X sky130_fd_sc_hd__a21o_1
XPHY_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06658_ _15338_/Q vssd1 vssd1 vccd1 vccd1 _06658_/Y sky130_fd_sc_hd__inv_2
XPHY_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_287 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09377_ _13898_/Q _13123_/B _08512_/B _14413_/Q _13123_/A vssd1 vssd1 vccd1 vccd1
+ _09377_/X sky130_fd_sc_hd__a221o_1
XFILLER_33_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_782 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08328_ _11045_/B _11033_/A vssd1 vssd1 vccd1 vccd1 _08328_/X sky130_fd_sc_hd__or2_1
XFILLER_149_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08259_ _11356_/B _08259_/B vssd1 vssd1 vccd1 vccd1 _08259_/Y sky130_fd_sc_hd__nor2_4
XFILLER_126_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11270_ _11344_/A _08249_/Y _08274_/X _08232_/A vssd1 vssd1 vccd1 vccd1 _11270_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_109_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10221_ input16/X _09382_/A _13291_/S vssd1 vssd1 vccd1 vccd1 _14606_/D sky130_fd_sc_hd__mux2_1
XFILLER_3_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10152_ _14537_/Q _11838_/A1 _10164_/S vssd1 vssd1 vccd1 vccd1 _14537_/D sky130_fd_sc_hd__mux2_1
XFILLER_79_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10083_ _14439_/Q _13336_/A0 _10097_/S vssd1 vssd1 vccd1 vccd1 _14439_/D sky130_fd_sc_hd__mux2_1
X_14960_ _15581_/CLK _14960_/D vssd1 vssd1 vccd1 vccd1 _14960_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_181_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold9 hold9/A vssd1 vssd1 vccd1 vccd1 hold9/X sky130_fd_sc_hd__bufbuf_16
XFILLER_59_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13911_ _15507_/CLK _13911_/D vssd1 vssd1 vccd1 vccd1 _13911_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14891_ _15622_/CLK _14891_/D vssd1 vssd1 vccd1 vccd1 _14891_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13842_ _15326_/CLK _13842_/D vssd1 vssd1 vccd1 vccd1 _13842_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13773_ _14863_/CLK _13773_/D vssd1 vssd1 vccd1 vccd1 _13773_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10985_ _11025_/A _11440_/A _08355_/A vssd1 vssd1 vccd1 vccd1 _10985_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_167_1071 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15512_ _15525_/CLK _15512_/D vssd1 vssd1 vccd1 vccd1 _15512_/Q sky130_fd_sc_hd__dfxtp_1
X_12724_ _15351_/Q _12723_/C _15352_/Q vssd1 vssd1 vccd1 vccd1 _12725_/B sky130_fd_sc_hd__a21oi_1
XFILLER_71_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_1066 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15443_ _15632_/CLK _15443_/D vssd1 vssd1 vccd1 vccd1 _15443_/Q sky130_fd_sc_hd__dfxtp_1
X_12655_ _12743_/A _12655_/B vssd1 vssd1 vccd1 vccd1 _12655_/X sky130_fd_sc_hd__or2_1
XFILLER_90_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11606_ _11606_/A _11606_/B _11606_/C vssd1 vssd1 vccd1 vccd1 _11606_/X sky130_fd_sc_hd__or3_1
XFILLER_50_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15374_ _15374_/CLK _15374_/D vssd1 vssd1 vccd1 vccd1 _15374_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_156_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12586_ _12590_/A _12586_/B vssd1 vssd1 vccd1 vccd1 _12586_/X sky130_fd_sc_hd__and2_1
X_14325_ _14606_/CLK _14325_/D vssd1 vssd1 vccd1 vccd1 _14325_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11537_ _11537_/A _11537_/B vssd1 vssd1 vccd1 vccd1 _11569_/D sky130_fd_sc_hd__and2_1
XFILLER_172_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14256_ _14482_/CLK _14256_/D vssd1 vssd1 vccd1 vccd1 _14256_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11468_ _11475_/A _11468_/B vssd1 vssd1 vccd1 vccd1 _11470_/B sky130_fd_sc_hd__xnor2_1
XFILLER_125_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13207_ _15569_/Q _13214_/B _13205_/X _13206_/Y vssd1 vssd1 vccd1 vccd1 _15569_/D
+ sky130_fd_sc_hd__a22o_1
X_10419_ _13252_/A _13251_/B vssd1 vssd1 vccd1 vccd1 _10420_/B sky130_fd_sc_hd__nand2_1
X_14187_ _15518_/CLK _14187_/D vssd1 vssd1 vccd1 vccd1 _14187_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_5_24_0_clk clkbuf_5_25_0_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_5_24_0_clk/X
+ sky130_fd_sc_hd__clkbuf_8
X_11399_ _11399_/A _11399_/B vssd1 vssd1 vccd1 vccd1 _11400_/B sky130_fd_sc_hd__nor2_1
XTAP_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13138_ _15535_/Q _08465_/X _13138_/S vssd1 vssd1 vccd1 vccd1 _15535_/D sky130_fd_sc_hd__mux2_1
XFILLER_135_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13069_ _15502_/Q _13119_/S _13105_/B1 _13068_/X vssd1 vssd1 vccd1 vccd1 _15502_/D
+ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_2_clk clkbuf_5_0_0_clk/X vssd1 vssd1 vccd1 vccd1 _15220_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_24_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07630_ _14758_/Q _07629_/A _07629_/Y _08002_/C1 vssd1 vssd1 vccd1 vccd1 _13469_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_65_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1014 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07561_ _07576_/C _07560_/Y _07651_/A vssd1 vssd1 vccd1 vccd1 _07561_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_34_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09300_ _08519_/B _09298_/X _09299_/X _08510_/B vssd1 vssd1 vccd1 vccd1 _09300_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07492_ _14763_/Q _07491_/X _07500_/S vssd1 vssd1 vccd1 vccd1 _07492_/X sky130_fd_sc_hd__mux2_4
XFILLER_181_1035 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09231_ _13891_/Q _09231_/A2 _09403_/B1 _14406_/Q _09445_/C1 vssd1 vssd1 vccd1 vccd1
+ _09231_/X sky130_fd_sc_hd__a221o_1
XFILLER_61_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_179_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_1019 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09162_ _09437_/A1 _09159_/X _09161_/X _09405_/A vssd1 vssd1 vccd1 vccd1 _09162_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_119_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08113_ input15/X input24/X _08145_/S vssd1 vssd1 vccd1 vccd1 _08167_/B sky130_fd_sc_hd__mux2_1
X_09093_ _14527_/Q _14140_/Q _14172_/Q _14108_/Q _09425_/S _09427_/A1 vssd1 vssd1
+ vccd1 vccd1 _09093_/X sky130_fd_sc_hd__mux4_1
XFILLER_108_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08044_ _14737_/Q _13615_/Q _08072_/S vssd1 vssd1 vccd1 vccd1 _13615_/D sky130_fd_sc_hd__mux2_1
XFILLER_135_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_362 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09995_ _13349_/A0 _14354_/Q _09996_/S vssd1 vssd1 vccd1 vccd1 _14354_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08946_ _15110_/Q _09558_/A2 _08520_/B _08945_/X vssd1 vssd1 vccd1 vccd1 _08946_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_9_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08877_ _13898_/Q _13098_/B2 _08885_/S vssd1 vssd1 vccd1 vccd1 _13898_/D sky130_fd_sc_hd__mux2_1
XFILLER_85_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07828_ _14745_/Q _07830_/A _07827_/Y _12788_/C1 vssd1 vssd1 vccd1 vccd1 _13520_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_3849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07759_ _14760_/Q _07777_/A _07758_/Y _08016_/C1 vssd1 vssd1 vccd1 vccd1 _13503_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_37_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10770_ _14802_/Q _15434_/Q _12906_/S vssd1 vssd1 vccd1 vccd1 _14802_/D sky130_fd_sc_hd__mux2_1
XFILLER_25_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09429_ _14543_/Q _14156_/Q _14188_/Q _14124_/Q _09190_/S _09429_/S1 vssd1 vssd1
+ vccd1 vccd1 _09429_/X sky130_fd_sc_hd__mux4_1
XFILLER_185_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_51 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12440_ _15132_/Q _15100_/Q _15673_/Q _13407_/Q _12453_/S _12452_/A vssd1 vssd1 vccd1
+ vccd1 _12440_/X sky130_fd_sc_hd__mux4_1
XFILLER_138_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12371_ _15129_/Q _15097_/Q _15670_/Q _13404_/Q _12522_/S _12521_/A vssd1 vssd1 vccd1
+ vccd1 _12371_/X sky130_fd_sc_hd__mux4_1
XFILLER_154_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14110_ _15253_/CLK _14110_/D vssd1 vssd1 vccd1 vccd1 _14110_/Q sky130_fd_sc_hd__dfxtp_1
X_11322_ _15037_/Q _11302_/A _11321_/X vssd1 vssd1 vccd1 vccd1 _15037_/D sky130_fd_sc_hd__o21a_1
XFILLER_176_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15090_ _15658_/CLK _15090_/D vssd1 vssd1 vccd1 vccd1 _15090_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_180_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14041_ _15178_/CLK _14041_/D vssd1 vssd1 vccd1 vccd1 _14041_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11253_ _11252_/A _08367_/X _11252_/Y vssd1 vssd1 vccd1 vccd1 _11311_/B sky130_fd_sc_hd__a21oi_1
XFILLER_140_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10204_ input29/X _14589_/Q _13284_/S vssd1 vssd1 vccd1 vccd1 _14589_/D sky130_fd_sc_hd__mux2_1
X_11184_ _14984_/Q _11202_/A _11183_/X vssd1 vssd1 vccd1 vccd1 _14984_/D sky130_fd_sc_hd__o21a_1
XFILLER_122_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10135_ _14520_/Q _13321_/A0 _10164_/S vssd1 vssd1 vccd1 vccd1 _14520_/D sky130_fd_sc_hd__mux2_1
XFILLER_67_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14943_ _15580_/CLK _14943_/D vssd1 vssd1 vccd1 vccd1 _14943_/Q sky130_fd_sc_hd__dfxtp_1
X_10066_ _14422_/Q _11852_/A1 _10092_/S vssd1 vssd1 vccd1 vccd1 _14422_/D sky130_fd_sc_hd__mux2_1
XFILLER_76_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14874_ _15592_/CLK _14874_/D vssd1 vssd1 vccd1 vccd1 _14874_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13825_ _15298_/CLK _13825_/D vssd1 vssd1 vccd1 vccd1 _13825_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13756_ _14888_/CLK _13756_/D vssd1 vssd1 vccd1 vccd1 _13756_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_188_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10968_ _11272_/A _11258_/A vssd1 vssd1 vccd1 vccd1 _10972_/B sky130_fd_sc_hd__nor2_1
XFILLER_90_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12707_ _12737_/A _12707_/B vssd1 vssd1 vccd1 vccd1 _12707_/X sky130_fd_sc_hd__or2_1
XFILLER_149_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13687_ _15178_/CLK _13687_/D vssd1 vssd1 vccd1 vccd1 _13687_/Q sky130_fd_sc_hd__dfxtp_1
X_10899_ _14932_/Q _10951_/B _10898_/Y _11362_/B vssd1 vssd1 vccd1 vccd1 _14932_/D
+ sky130_fd_sc_hd__o22a_1
X_15426_ _15623_/CLK _15426_/D vssd1 vssd1 vccd1 vccd1 _15426_/Q sky130_fd_sc_hd__dfxtp_2
X_12638_ _15047_/Q _12637_/Y _12834_/B vssd1 vssd1 vccd1 vccd1 _12638_/X sky130_fd_sc_hd__mux2_1
XFILLER_157_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15357_ _15637_/CLK _15357_/D vssd1 vssd1 vccd1 vccd1 _15357_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_156_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12569_ _12592_/A1 _12568_/X _06670_/A vssd1 vssd1 vccd1 vccd1 _12569_/X sky130_fd_sc_hd__a21o_1
XFILLER_157_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14308_ _15289_/CLK _14308_/D vssd1 vssd1 vccd1 vccd1 _14308_/Q sky130_fd_sc_hd__dfxtp_1
X_15288_ _15332_/CLK _15288_/D vssd1 vssd1 vccd1 vccd1 _15288_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14239_ _15663_/CLK _14239_/D vssd1 vssd1 vccd1 vccd1 _14239_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_131_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08800_ _13334_/A0 _13826_/Q _08811_/S vssd1 vssd1 vccd1 vccd1 _13826_/D sky130_fd_sc_hd__mux2_1
XTAP_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09780_ _14147_/Q _13335_/A0 _09790_/S vssd1 vssd1 vccd1 vccd1 _14147_/D sky130_fd_sc_hd__mux2_1
XTAP_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06992_ _10507_/A1 _13120_/S _06797_/Y _08777_/A _06991_/X vssd1 vssd1 vccd1 vccd1
+ _14582_/D sky130_fd_sc_hd__a221o_1
XTAP_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08731_ _13448_/Q _08746_/A2 _08727_/X _08728_/X _08730_/X vssd1 vssd1 vccd1 vccd1
+ _08731_/X sky130_fd_sc_hd__a2111o_1
XTAP_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08662_ _13457_/Q _08684_/A2 _08691_/B1 _13489_/Q _08661_/X vssd1 vssd1 vccd1 vccd1
+ _08662_/X sky130_fd_sc_hd__a221o_1
XFILLER_38_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07613_ _13465_/Q _07617_/C vssd1 vssd1 vccd1 vccd1 _07614_/B sky130_fd_sc_hd__xnor2_1
XFILLER_53_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08593_ _13467_/Q _08684_/A2 _08750_/B1 _13634_/Q vssd1 vssd1 vccd1 vccd1 _08593_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_81_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07544_ _13447_/Q _13446_/Q _13445_/Q vssd1 vssd1 vccd1 vccd1 _07549_/B sky130_fd_sc_hd__and3_1
XFILLER_34_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07475_ _13674_/Q _07483_/A2 _07483_/B1 _14702_/Q _07474_/X vssd1 vssd1 vccd1 vccd1
+ _07475_/X sky130_fd_sc_hd__a221o_1
XFILLER_22_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09214_ _15123_/Q _09449_/A1 _09445_/A2 _09450_/B1 vssd1 vssd1 vccd1 vccd1 _09214_/X
+ sky130_fd_sc_hd__a31o_1
X_09145_ _14434_/Q _13130_/B1 _09144_/X _06676_/A vssd1 vssd1 vccd1 vccd1 _09145_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_136_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09076_ _08520_/B _09073_/X _09075_/X _09071_/X vssd1 vssd1 vccd1 vccd1 _09077_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_146_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08027_ _08027_/A _08033_/B vssd1 vssd1 vccd1 vccd1 _08027_/X sky130_fd_sc_hd__or2_1
XFILLER_1_415 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09978_ _13332_/A0 _14337_/Q _09991_/S vssd1 vssd1 vccd1 vccd1 _14337_/D sky130_fd_sc_hd__mux2_1
XFILLER_131_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08929_ _09543_/A _08929_/B vssd1 vssd1 vccd1 vccd1 _08929_/X sky130_fd_sc_hd__or2_1
XFILLER_188_1019 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11940_ _12618_/A1 _11935_/X _11938_/X _11939_/X _08405_/D vssd1 vssd1 vccd1 vccd1
+ _11952_/B sky130_fd_sc_hd__a221o_1
XFILLER_45_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_176_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11871_ _15292_/Q _13338_/A0 _11883_/S vssd1 vssd1 vccd1 vccd1 _15292_/D sky130_fd_sc_hd__mux2_1
XTAP_2934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13610_ _15461_/CLK _13610_/D vssd1 vssd1 vccd1 vccd1 _13610_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_2956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10822_ _14854_/Q _07219_/X _10868_/S vssd1 vssd1 vccd1 vccd1 _14854_/D sky130_fd_sc_hd__mux2_1
XFILLER_72_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14590_ _14612_/CLK _14590_/D vssd1 vssd1 vccd1 vccd1 hold5/A sky130_fd_sc_hd__dfxtp_2
XTAP_2978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13541_ _15542_/CLK _13541_/D vssd1 vssd1 vccd1 vccd1 _13541_/Q sky130_fd_sc_hd__dfxtp_2
X_10753_ _15417_/Q _14785_/Q _10765_/S vssd1 vssd1 vccd1 vccd1 _14785_/D sky130_fd_sc_hd__mux2_1
XFILLER_13_544 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_875 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13472_ _14513_/CLK _13472_/D vssd1 vssd1 vccd1 vccd1 _13472_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10684_ _15064_/Q _10714_/A2 _10681_/X _10683_/X vssd1 vssd1 vccd1 vccd1 _10684_/X
+ sky130_fd_sc_hd__o22a_4
XFILLER_9_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15211_ _15211_/CLK _15211_/D vssd1 vssd1 vccd1 vccd1 _15211_/Q sky130_fd_sc_hd__dfxtp_1
X_12423_ _06671_/Y _12418_/X _12421_/X _12422_/X _08405_/D vssd1 vssd1 vccd1 vccd1
+ _12435_/B sky130_fd_sc_hd__a221o_1
XFILLER_127_914 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15142_ _15142_/CLK _15142_/D vssd1 vssd1 vccd1 vccd1 _15142_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_153_210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12354_ _12595_/A1 _12349_/X _12352_/X _12353_/X _08405_/D vssd1 vssd1 vccd1 vccd1
+ _12366_/B sky130_fd_sc_hd__a221o_1
XFILLER_153_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11305_ _11330_/A _11305_/B _11305_/C vssd1 vssd1 vccd1 vccd1 _11305_/X sky130_fd_sc_hd__and3_1
X_15073_ _15613_/CLK _15073_/D vssd1 vssd1 vccd1 vccd1 _15073_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_4_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12285_ _12595_/A1 _12280_/X _12283_/X _12284_/X _08405_/D vssd1 vssd1 vccd1 vccd1
+ _12297_/B sky130_fd_sc_hd__a221o_1
XFILLER_84_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14024_ _15334_/CLK _14024_/D vssd1 vssd1 vccd1 vccd1 _14024_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11236_ _10430_/B _15024_/Q _11237_/S vssd1 vssd1 vccd1 vccd1 _15024_/D sky130_fd_sc_hd__mux2_1
XFILLER_136_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11167_ _13251_/B _11389_/B _11414_/A vssd1 vssd1 vccd1 vccd1 _11167_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_171_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10118_ _14504_/Q _14752_/Q _10124_/S vssd1 vssd1 vccd1 vccd1 _14504_/D sky130_fd_sc_hd__mux2_1
XFILLER_49_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11098_ _10973_/Y _10993_/Y _11297_/S vssd1 vssd1 vccd1 vccd1 _11098_/X sky130_fd_sc_hd__mux2_1
X_10049_ _14406_/Q _11868_/A1 _10059_/S vssd1 vssd1 vccd1 vccd1 _14406_/D sky130_fd_sc_hd__mux2_1
X_14926_ _15536_/CLK _15536_/Q vssd1 vssd1 vccd1 vccd1 _14926_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14857_ _15519_/CLK _14857_/D vssd1 vssd1 vccd1 vccd1 _14857_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_230 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13808_ _15208_/CLK _13808_/D vssd1 vssd1 vccd1 vccd1 _13808_/Q sky130_fd_sc_hd__dfxtp_1
X_14788_ _15638_/CLK _14788_/D vssd1 vssd1 vccd1 vccd1 _14788_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13739_ _14863_/CLK _13739_/D vssd1 vssd1 vccd1 vccd1 _13739_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_91_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07260_ _07260_/A _07260_/B vssd1 vssd1 vccd1 vccd1 _07270_/B sky130_fd_sc_hd__nor2_1
X_15409_ _15599_/CLK _15409_/D vssd1 vssd1 vccd1 vccd1 _15409_/Q sky130_fd_sc_hd__dfxtp_2
X_07191_ _15365_/Q _15072_/Q _07193_/S vssd1 vssd1 vccd1 vccd1 _07191_/X sky130_fd_sc_hd__mux2_4
XFILLER_118_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09901_ _13321_/A0 _14262_/Q _09930_/S vssd1 vssd1 vccd1 vccd1 _14262_/D sky130_fd_sc_hd__mux2_1
XFILLER_126_991 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout505 _14733_/Q vssd1 vssd1 vccd1 vccd1 _07096_/S sky130_fd_sc_hd__buf_12
Xfanout516 _09554_/A vssd1 vssd1 vccd1 vccd1 _09524_/A sky130_fd_sc_hd__buf_12
X_09832_ _14196_/Q _11852_/A1 _09858_/S vssd1 vssd1 vccd1 vccd1 _14196_/D sky130_fd_sc_hd__mux2_1
Xfanout527 _08988_/A1 vssd1 vssd1 vccd1 vccd1 _09427_/A1 sky130_fd_sc_hd__buf_6
Xfanout538 _09553_/A1 vssd1 vssd1 vccd1 vccd1 _09550_/A1 sky130_fd_sc_hd__buf_12
XFILLER_99_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout549 _09047_/S vssd1 vssd1 vccd1 vccd1 _09073_/S sky130_fd_sc_hd__buf_6
XFILLER_113_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09763_ _11818_/A _10132_/B vssd1 vssd1 vccd1 vccd1 _09763_/Y sky130_fd_sc_hd__nor2_8
X_06975_ _06954_/X _06958_/X _06964_/Y _06974_/X vssd1 vssd1 vccd1 vccd1 _06975_/Y
+ sky130_fd_sc_hd__a31oi_2
XTAP_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08714_ _13585_/Q _08749_/A2 _08747_/A2 _13546_/Q vssd1 vssd1 vccd1 vccd1 _08714_/X
+ sky130_fd_sc_hd__a22o_1
X_09694_ _14065_/Q _11816_/A1 _09695_/S vssd1 vssd1 vccd1 vccd1 _14065_/D sky130_fd_sc_hd__mux2_1
XFILLER_27_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08645_ _08722_/A _08645_/B _08645_/C vssd1 vssd1 vccd1 vccd1 _08645_/X sky130_fd_sc_hd__or3_4
XFILLER_187_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_14 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08576_ _15393_/Q _08748_/A2 _08736_/A2 _13438_/Q vssd1 vssd1 vccd1 vccd1 _08576_/X
+ sky130_fd_sc_hd__a22o_1
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07527_ _14757_/Q _13436_/Q _07529_/S vssd1 vssd1 vccd1 vccd1 _13436_/D sky130_fd_sc_hd__mux2_1
XFILLER_167_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07458_ _14666_/Q _07490_/B _14710_/Q vssd1 vssd1 vccd1 vccd1 _07458_/X sky130_fd_sc_hd__and3_1
XFILLER_23_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07389_ _11680_/A0 _13386_/Q _07481_/S vssd1 vssd1 vccd1 vccd1 _13386_/D sky130_fd_sc_hd__mux2_1
XFILLER_41_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09128_ _14078_/Q _09231_/A2 _09403_/B1 _14046_/Q _09221_/A vssd1 vssd1 vccd1 vccd1
+ _09128_/X sky130_fd_sc_hd__a221o_1
XFILLER_109_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09059_ _14011_/Q _13979_/Q _09230_/S vssd1 vssd1 vccd1 vccd1 _09059_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12070_ _14462_/Q _14430_/Q _13851_/Q _14204_/Q _12470_/S _12080_/A vssd1 vssd1 vccd1
+ vccd1 _12070_/X sky130_fd_sc_hd__mux4_1
XFILLER_123_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11021_ _11017_/X _11020_/Y _11318_/S vssd1 vssd1 vccd1 vccd1 _11021_/X sky130_fd_sc_hd__mux2_1
XFILLER_77_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12972_ _10624_/X _14871_/Q _13029_/S vssd1 vssd1 vccd1 vccd1 _12972_/X sky130_fd_sc_hd__mux2_8
XFILLER_46_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11923_ _12383_/A _11923_/B vssd1 vssd1 vccd1 vccd1 _11923_/X sky130_fd_sc_hd__and2_1
XFILLER_73_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14711_ _15530_/CLK _14711_/D vssd1 vssd1 vccd1 vccd1 _14711_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14642_ _15645_/CLK _14642_/D vssd1 vssd1 vccd1 vccd1 _14642_/Q sky130_fd_sc_hd__dfxtp_1
X_11854_ _15275_/Q _11854_/A1 _11883_/S vssd1 vssd1 vccd1 vccd1 _15275_/D sky130_fd_sc_hd__mux2_1
XTAP_2764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10805_ _14837_/Q _07352_/A _13138_/S vssd1 vssd1 vccd1 vccd1 _14837_/D sky130_fd_sc_hd__mux2_1
XTAP_2797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14573_ _15336_/CLK _14573_/D vssd1 vssd1 vccd1 vccd1 _14573_/Q sky130_fd_sc_hd__dfxtp_1
X_11785_ _13318_/D _11851_/B vssd1 vssd1 vccd1 vccd1 _11785_/Y sky130_fd_sc_hd__nor2_8
X_13524_ _13627_/CLK _13524_/D vssd1 vssd1 vccd1 vccd1 _13524_/Q sky130_fd_sc_hd__dfxtp_1
X_10736_ _15400_/Q _14768_/Q _13129_/A vssd1 vssd1 vccd1 vccd1 _14768_/D sky130_fd_sc_hd__mux2_1
XFILLER_9_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13455_ _15377_/CLK _13455_/D vssd1 vssd1 vccd1 vccd1 _13455_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10667_ _15012_/Q _10717_/A2 _10602_/B _15029_/Q _10717_/C1 vssd1 vssd1 vccd1 vccd1
+ _10667_/X sky130_fd_sc_hd__a221o_1
X_12406_ _12406_/A _12406_/B vssd1 vssd1 vccd1 vccd1 _12406_/X sky130_fd_sc_hd__and2_1
XFILLER_12_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13386_ _15652_/CLK _13386_/D vssd1 vssd1 vccd1 vccd1 _13386_/Q sky130_fd_sc_hd__dfxtp_1
X_10598_ _13717_/Q _10602_/B _10597_/X vssd1 vssd1 vccd1 vccd1 _10598_/X sky130_fd_sc_hd__a21o_1
XFILLER_182_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15125_ _15125_/CLK _15125_/D vssd1 vssd1 vccd1 vccd1 _15125_/Q sky130_fd_sc_hd__dfxtp_1
X_12337_ _12544_/A _12337_/B vssd1 vssd1 vccd1 vccd1 _12337_/X sky130_fd_sc_hd__and2_1
XFILLER_115_939 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15056_ _15599_/CLK _15056_/D vssd1 vssd1 vccd1 vccd1 _15056_/Q sky130_fd_sc_hd__dfxtp_4
X_12268_ _12268_/A _12268_/B vssd1 vssd1 vccd1 vccd1 _12268_/X sky130_fd_sc_hd__and2_1
X_14007_ _15253_/CLK _14007_/D vssd1 vssd1 vccd1 vccd1 _14007_/Q sky130_fd_sc_hd__dfxtp_1
X_11219_ _10366_/B _10390_/B _11232_/S _11218_/Y vssd1 vssd1 vccd1 vccd1 _15007_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_122_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12199_ _12498_/A _12199_/B vssd1 vssd1 vccd1 vccd1 _12199_/X sky130_fd_sc_hd__and2_1
Xoutput90 _07161_/X vssd1 vssd1 vccd1 vccd1 ext_write_data[30] sky130_fd_sc_hd__clkbuf_2
XFILLER_96_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_772 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06760_ input18/X vssd1 vssd1 vccd1 vccd1 _06760_/Y sky130_fd_sc_hd__inv_2
X_14909_ _15499_/CLK _14909_/D vssd1 vssd1 vccd1 vccd1 _14909_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_37_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06691_ _13475_/Q vssd1 vssd1 vccd1 vccd1 _06691_/Y sky130_fd_sc_hd__inv_2
XFILLER_64_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08430_ _13745_/Q _12878_/S _08426_/B _08429_/X vssd1 vssd1 vccd1 vccd1 _13745_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_63_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08361_ _11023_/A _08361_/B vssd1 vssd1 vccd1 vccd1 _11034_/B sky130_fd_sc_hd__nor2_1
XFILLER_177_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_1091 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07312_ _13913_/Q _15500_/Q _07334_/S vssd1 vssd1 vccd1 vccd1 _07312_/X sky130_fd_sc_hd__mux2_8
XFILLER_108_1042 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08292_ _11297_/S _08292_/B vssd1 vssd1 vccd1 vccd1 _08299_/B sky130_fd_sc_hd__or2_1
XFILLER_165_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07243_ _15327_/Q _15483_/Q _07335_/S vssd1 vssd1 vccd1 vccd1 _07244_/A sky130_fd_sc_hd__mux2_8
XFILLER_176_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07174_ _15348_/Q _15055_/Q _07188_/S vssd1 vssd1 vccd1 vccd1 _07174_/X sky130_fd_sc_hd__mux2_8
XFILLER_11_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_883 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout302 _07464_/X vssd1 vssd1 vccd1 vccd1 _13341_/A0 sky130_fd_sc_hd__buf_4
Xfanout313 _13086_/B2 vssd1 vssd1 vccd1 vccd1 _13336_/A0 sky130_fd_sc_hd__buf_2
XFILLER_120_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout324 _07424_/X vssd1 vssd1 vccd1 vccd1 _11689_/A0 sky130_fd_sc_hd__buf_4
XFILLER_59_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout335 _13325_/A0 vssd1 vssd1 vccd1 vccd1 _11858_/A1 sky130_fd_sc_hd__buf_6
XFILLER_115_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout346 _13320_/A0 vssd1 vssd1 vccd1 vccd1 _11853_/A1 sky130_fd_sc_hd__buf_6
X_09815_ _14181_/Q _13337_/A0 _09828_/S vssd1 vssd1 vccd1 vccd1 _14181_/D sky130_fd_sc_hd__mux2_1
Xfanout357 _10569_/Y vssd1 vssd1 vccd1 vccd1 _10734_/A2 sky130_fd_sc_hd__buf_12
Xfanout368 _08507_/Y vssd1 vssd1 vccd1 vccd1 _09421_/A1 sky130_fd_sc_hd__buf_12
XFILLER_87_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout379 _11053_/S vssd1 vssd1 vccd1 vccd1 _11356_/B sky130_fd_sc_hd__buf_12
XFILLER_115_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09746_ _14114_/Q _13334_/A0 _09757_/S vssd1 vssd1 vccd1 vccd1 _14114_/D sky130_fd_sc_hd__mux2_1
X_06958_ _06941_/A _06957_/X _06936_/Y vssd1 vssd1 vccd1 vccd1 _06958_/X sky130_fd_sc_hd__a21bo_1
XFILLER_27_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09677_ _14048_/Q _13078_/B2 _09690_/S vssd1 vssd1 vccd1 vccd1 _14048_/D sky130_fd_sc_hd__mux2_1
XTAP_2016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06889_ _15395_/Q _06699_/Y _15394_/Q _06701_/Y _06888_/Y vssd1 vssd1 vccd1 vccd1
+ _06889_/X sky130_fd_sc_hd__o221a_1
XTAP_2027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08628_ _13597_/Q _08691_/A2 _08685_/A2 _13558_/Q _08627_/X vssd1 vssd1 vccd1 vccd1
+ _08632_/B sky130_fd_sc_hd__a221o_1
XFILLER_42_403 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08559_ _08722_/A _08559_/B _08559_/C vssd1 vssd1 vccd1 vccd1 _08559_/X sky130_fd_sc_hd__or3_1
XFILLER_30_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11570_ _13236_/A _11589_/C vssd1 vssd1 vccd1 vccd1 _11571_/B sky130_fd_sc_hd__or2_4
XFILLER_74_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_1044 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10521_ _07264_/A _10360_/B _10520_/X vssd1 vssd1 vccd1 vccd1 _13214_/A sky130_fd_sc_hd__a21oi_4
XFILLER_22_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13240_ _13217_/A wire360/X _13241_/A2 vssd1 vssd1 vccd1 vccd1 _13240_/Y sky130_fd_sc_hd__a21oi_1
X_10452_ _07221_/A _10481_/B _10451_/X vssd1 vssd1 vccd1 vccd1 _11584_/A sky130_fd_sc_hd__a21o_4
XFILLER_109_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13171_ _13251_/A _13171_/B vssd1 vssd1 vccd1 vccd1 _13171_/Y sky130_fd_sc_hd__nor2_1
X_10383_ _13195_/B _11475_/A vssd1 vssd1 vccd1 vccd1 _10384_/A sky130_fd_sc_hd__nand2_1
XFILLER_164_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12122_ _12490_/A _12122_/B vssd1 vssd1 vccd1 vccd1 _12122_/X sky130_fd_sc_hd__or2_1
XFILLER_184_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_972 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12053_ _12260_/A _12053_/B vssd1 vssd1 vccd1 vccd1 _12053_/X sky130_fd_sc_hd__or2_1
XFILLER_89_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11004_ _14962_/Q _11003_/X _11202_/A vssd1 vssd1 vccd1 vccd1 _14962_/D sky130_fd_sc_hd__mux2_1
XFILLER_120_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_3_6_0_clk clkbuf_3_7_0_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_6_0_clk/X sky130_fd_sc_hd__clkbuf_8
XFILLER_58_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12955_ _07388_/X _13024_/A2 _12954_/X _13024_/B2 vssd1 vssd1 vccd1 vccd1 _12955_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_3251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11906_ _12596_/A _11906_/B _11906_/C vssd1 vssd1 vccd1 vccd1 _11906_/X sky130_fd_sc_hd__and3_4
XTAP_3284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12886_ _15414_/Q _15599_/Q _12917_/S vssd1 vssd1 vccd1 vccd1 _15414_/D sky130_fd_sc_hd__mux2_1
XTAP_3295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15674_ _15674_/CLK _15674_/D vssd1 vssd1 vccd1 vccd1 _15674_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14625_ _15596_/CLK _14625_/D vssd1 vssd1 vccd1 vccd1 _14625_/Q sky130_fd_sc_hd__dfxtp_1
X_11837_ _15259_/Q _11870_/A1 _11850_/S vssd1 vssd1 vccd1 vccd1 _15259_/D sky130_fd_sc_hd__mux2_1
XFILLER_61_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1103 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_110 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14556_ _15279_/CLK _14556_/D vssd1 vssd1 vccd1 vccd1 _14556_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11768_ _13343_/A0 _15196_/Q _11774_/S vssd1 vssd1 vccd1 vccd1 _15196_/D sky130_fd_sc_hd__mux2_1
XFILLER_147_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13507_ _13642_/CLK _13507_/D vssd1 vssd1 vccd1 vccd1 _13507_/Q sky130_fd_sc_hd__dfxtp_2
X_10719_ _15071_/Q _10734_/A2 _10716_/X _10718_/X vssd1 vssd1 vccd1 vccd1 _10719_/X
+ sky130_fd_sc_hd__o22a_4
XFILLER_9_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14487_ _15542_/CLK _14487_/D vssd1 vssd1 vccd1 vccd1 _14487_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_173_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11699_ _13341_/A0 _15130_/Q _11703_/S vssd1 vssd1 vccd1 vccd1 _15130_/D sky130_fd_sc_hd__mux2_1
XFILLER_173_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13438_ _15393_/CLK _13438_/D vssd1 vssd1 vccd1 vccd1 _13438_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_174_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_248_clk clkbuf_5_4_0_clk/X vssd1 vssd1 vccd1 vccd1 _15184_/CLK sky130_fd_sc_hd__clkbuf_16
X_13369_ _14472_/Q vssd1 vssd1 vccd1 vccd1 _14472_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_54_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15108_ _15108_/CLK _15108_/D vssd1 vssd1 vccd1 vccd1 _15108_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_142_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15039_ _15041_/CLK _15039_/D vssd1 vssd1 vccd1 vccd1 _15039_/Q sky130_fd_sc_hd__dfxtp_1
X_07930_ _07932_/B _07929_/X _08012_/A2 vssd1 vssd1 vccd1 vccd1 _07930_/X sky130_fd_sc_hd__a21bo_1
XFILLER_69_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07861_ _14754_/Q _07874_/A _07860_/Y _08002_/C1 vssd1 vssd1 vccd1 vccd1 _13529_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_111_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09600_ _13974_/Q _11680_/A0 _09627_/S vssd1 vssd1 vccd1 vccd1 _13974_/D sky130_fd_sc_hd__mux2_1
X_06812_ _13732_/Q _08668_/B _09382_/A _06664_/Y vssd1 vssd1 vccd1 vccd1 _06812_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_95_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07792_ _07816_/A _07792_/B vssd1 vssd1 vccd1 vccd1 _07792_/Y sky130_fd_sc_hd__nand2_1
X_09531_ _14386_/Q _15202_/Q _13841_/Q _14580_/Q _09521_/S _08494_/B vssd1 vssd1 vccd1
+ vccd1 _09532_/B sky130_fd_sc_hd__mux4_1
XFILLER_3_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06743_ _13482_/Q vssd1 vssd1 vccd1 vccd1 _06743_/Y sky130_fd_sc_hd__inv_2
XFILLER_52_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09462_ _08510_/B _09460_/X _09461_/X _08519_/B _13131_/A vssd1 vssd1 vccd1 vccd1
+ _09462_/X sky130_fd_sc_hd__a221o_1
XFILLER_92_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06674_ _08508_/B vssd1 vssd1 vccd1 vccd1 _08668_/B sky130_fd_sc_hd__inv_6
XFILLER_19_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08413_ _13242_/A _13138_/S _08412_/X vssd1 vssd1 vccd1 vccd1 _08413_/X sky130_fd_sc_hd__o21a_1
XFILLER_52_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09393_ _09437_/A1 _09392_/X _09391_/X _09130_/A vssd1 vssd1 vccd1 vccd1 _09393_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_51_255 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08344_ _11449_/A vssd1 vssd1 vccd1 vccd1 _13189_/B sky130_fd_sc_hd__inv_2
XFILLER_149_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_631 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08275_ _11351_/C1 _08249_/Y _08274_/X _08232_/A _13716_/Q vssd1 vssd1 vccd1 vccd1
+ _13716_/D sky130_fd_sc_hd__a32o_1
XFILLER_138_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07226_ _07227_/A _07227_/B _07197_/X vssd1 vssd1 vccd1 vccd1 _07231_/C sky130_fd_sc_hd__a21o_1
XFILLER_118_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_239_clk clkbuf_5_5_0_clk/X vssd1 vssd1 vccd1 vccd1 _14462_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_164_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_179 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07157_ _07157_/A _07157_/B vssd1 vssd1 vccd1 vccd1 _07157_/X sky130_fd_sc_hd__and2_2
XFILLER_121_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07088_ _07087_/X _13608_/Q _12662_/S vssd1 vssd1 vccd1 vccd1 _07088_/X sky130_fd_sc_hd__mux2_1
XFILLER_160_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout110 _13288_/S vssd1 vssd1 vccd1 vccd1 _13300_/S sky130_fd_sc_hd__buf_12
Xfanout121 _10834_/S vssd1 vssd1 vccd1 vccd1 _13081_/A2 sky130_fd_sc_hd__buf_8
Xfanout132 fanout138/X vssd1 vssd1 vccd1 vccd1 _13129_/A sky130_fd_sc_hd__buf_12
Xfanout143 _12320_/A vssd1 vssd1 vccd1 vccd1 _10871_/S sky130_fd_sc_hd__buf_8
Xfanout154 _12927_/S vssd1 vssd1 vccd1 vccd1 _12918_/S sky130_fd_sc_hd__buf_6
Xfanout165 _12871_/S vssd1 vssd1 vccd1 vccd1 _12866_/S sky130_fd_sc_hd__buf_12
XFILLER_59_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout176 _11710_/Y vssd1 vssd1 vccd1 vccd1 _11742_/S sky130_fd_sc_hd__buf_12
XFILLER_47_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout187 _10032_/Y vssd1 vssd1 vccd1 vccd1 _10059_/S sky130_fd_sc_hd__buf_12
Xfanout198 _09865_/Y vssd1 vssd1 vccd1 vccd1 _09897_/S sky130_fd_sc_hd__buf_12
XFILLER_86_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09729_ _14715_/Q _13318_/C _14714_/Q vssd1 vssd1 vccd1 vccd1 _10132_/B sky130_fd_sc_hd__or3b_4
XFILLER_55_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12740_ _15061_/Q _12739_/X _12792_/B vssd1 vssd1 vccd1 vccd1 _12740_/X sky130_fd_sc_hd__mux2_1
XFILLER_16_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12671_ _12743_/A _12671_/B vssd1 vssd1 vccd1 vccd1 _12671_/X sky130_fd_sc_hd__or2_1
XTAP_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14410_ _15096_/CLK _14410_/D vssd1 vssd1 vccd1 vccd1 _14410_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11622_ _11621_/X _15071_/Q _11641_/S vssd1 vssd1 vccd1 vccd1 _15071_/D sky130_fd_sc_hd__mux2_1
XFILLER_24_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_187_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15390_ _15393_/CLK _15390_/D vssd1 vssd1 vccd1 vccd1 _15390_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14341_ _15125_/CLK _14341_/D vssd1 vssd1 vccd1 vccd1 _14341_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_168_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11553_ _11555_/A _11555_/B vssd1 vssd1 vccd1 vccd1 _11556_/A sky130_fd_sc_hd__or2_1
XFILLER_7_602 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10504_ _10543_/B _10542_/A vssd1 vssd1 vccd1 vccd1 _10527_/C sky130_fd_sc_hd__nand2_1
XFILLER_7_635 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14272_ _14530_/CLK _14272_/D vssd1 vssd1 vccd1 vccd1 _14272_/Q sky130_fd_sc_hd__dfxtp_1
X_11484_ _11505_/C _11484_/B vssd1 vssd1 vccd1 vccd1 _11484_/Y sky130_fd_sc_hd__nand2_1
XFILLER_144_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_171_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13223_ _13236_/A _13223_/B vssd1 vssd1 vccd1 vccd1 _13223_/Y sky130_fd_sc_hd__nor2_1
X_10435_ _11616_/A _13242_/B vssd1 vssd1 vccd1 vccd1 _10471_/B sky130_fd_sc_hd__xnor2_2
XFILLER_170_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13154_ _14614_/Q _15552_/Q _13154_/S vssd1 vssd1 vccd1 vccd1 _15552_/D sky130_fd_sc_hd__mux2_1
XFILLER_128_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10366_ _10366_/A _10366_/B _10366_/C vssd1 vssd1 vccd1 vccd1 _10557_/A sky130_fd_sc_hd__or3_2
XFILLER_3_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12105_ _12477_/A1 _12104_/X _12260_/A vssd1 vssd1 vccd1 vccd1 _12105_/X sky130_fd_sc_hd__a21o_1
XFILLER_69_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13085_ _15510_/Q _13119_/S _13105_/B1 _13084_/X vssd1 vssd1 vccd1 vccd1 _15510_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_88_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10297_ _14682_/Q _14867_/Q _10730_/S vssd1 vssd1 vccd1 vccd1 _14682_/D sky130_fd_sc_hd__mux2_1
XFILLER_78_631 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12036_ _12592_/A1 _12035_/X _12594_/S vssd1 vssd1 vccd1 vccd1 _12036_/X sky130_fd_sc_hd__a21o_1
XFILLER_78_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13987_ _14083_/CLK _13987_/D vssd1 vssd1 vccd1 vccd1 _13987_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12938_ _06671_/A _11743_/C _08817_/Y _06670_/A vssd1 vssd1 vccd1 vccd1 _12943_/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15657_ _15657_/CLK _15657_/D vssd1 vssd1 vccd1 vccd1 _15657_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12869_ _14763_/Q _15397_/Q _12871_/S vssd1 vssd1 vccd1 vccd1 _15397_/D sky130_fd_sc_hd__mux2_1
XFILLER_178_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14608_ _15461_/CLK _14608_/D vssd1 vssd1 vccd1 vccd1 _14608_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_1690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15588_ _15588_/CLK _15588_/D vssd1 vssd1 vccd1 vccd1 _15588_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_187_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14539_ _15161_/CLK _14539_/D vssd1 vssd1 vccd1 vccd1 _14539_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_179_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08060_ _14753_/Q _13631_/Q _08072_/S vssd1 vssd1 vccd1 vccd1 _13631_/D sky130_fd_sc_hd__mux2_1
XFILLER_119_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07011_ _07010_/X _14736_/Q _07098_/S vssd1 vssd1 vccd1 vccd1 _13582_/D sky130_fd_sc_hd__mux2_1
XFILLER_108_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08962_ _09530_/S1 _08960_/X _08961_/X vssd1 vssd1 vccd1 vccd1 _08962_/X sky130_fd_sc_hd__a21o_1
XFILLER_88_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07913_ _13543_/Q _13542_/Q _13541_/Q _07913_/D vssd1 vssd1 vccd1 vccd1 _07924_/D
+ sky130_fd_sc_hd__and4_2
X_08893_ _14003_/Q _13971_/Q _09230_/S vssd1 vssd1 vccd1 vccd1 _08893_/X sky130_fd_sc_hd__mux2_1
XFILLER_111_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07844_ _13525_/Q _07844_/B vssd1 vssd1 vccd1 vccd1 _07844_/X sky130_fd_sc_hd__xor2_1
XFILLER_151_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_859 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07775_ _13507_/Q _07776_/C _13508_/Q vssd1 vssd1 vccd1 vccd1 _07777_/B sky130_fd_sc_hd__a21bo_1
XFILLER_37_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09514_ _15137_/Q _09558_/A2 _09513_/X _08501_/A vssd1 vssd1 vccd1 vccd1 _09514_/X
+ sky130_fd_sc_hd__a211o_1
X_06726_ _13490_/Q vssd1 vssd1 vccd1 vccd1 _06726_/Y sky130_fd_sc_hd__inv_2
XFILLER_65_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09445_ _13901_/Q _09445_/A2 _09522_/B1 _14416_/Q _09445_/C1 vssd1 vssd1 vccd1 vccd1
+ _09445_/X sky130_fd_sc_hd__a221o_1
XFILLER_13_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09376_ _13962_/Q _13704_/Q _09512_/S vssd1 vssd1 vccd1 vccd1 _09376_/X sky130_fd_sc_hd__mux2_1
XFILLER_24_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08327_ _11037_/A _11431_/A vssd1 vssd1 vccd1 vccd1 _11033_/A sky130_fd_sc_hd__nor2_1
XFILLER_165_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_1088 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08258_ _08259_/B vssd1 vssd1 vccd1 vccd1 _08258_/Y sky130_fd_sc_hd__inv_2
XFILLER_166_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07209_ _13933_/Q _15520_/Q _07339_/S vssd1 vssd1 vccd1 vccd1 _07210_/A sky130_fd_sc_hd__mux2_8
X_08189_ _11710_/A _10032_/A vssd1 vssd1 vccd1 vccd1 _08189_/Y sky130_fd_sc_hd__nor2_8
XFILLER_165_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10220_ input15/X _09435_/A _13282_/S vssd1 vssd1 vccd1 vccd1 _14605_/D sky130_fd_sc_hd__mux2_1
XFILLER_165_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10151_ _14536_/Q _13337_/A0 _10164_/S vssd1 vssd1 vccd1 vccd1 _14536_/D sky130_fd_sc_hd__mux2_1
XFILLER_79_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_855 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10082_ _14438_/Q _11868_/A1 _10092_/S vssd1 vssd1 vccd1 vccd1 _14438_/D sky130_fd_sc_hd__mux2_1
X_13910_ _15497_/CLK _13910_/D vssd1 vssd1 vccd1 vccd1 _13910_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14890_ _15623_/CLK _14890_/D vssd1 vssd1 vccd1 vccd1 _14890_/Q sky130_fd_sc_hd__dfxtp_1
X_13841_ _15303_/CLK _13841_/D vssd1 vssd1 vccd1 vccd1 _13841_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13772_ _14861_/CLK _13772_/D vssd1 vssd1 vccd1 vccd1 _13772_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10984_ _14928_/D _14927_/D _14929_/D vssd1 vssd1 vccd1 vccd1 _10984_/Y sky130_fd_sc_hd__nand3b_4
XFILLER_55_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15511_ _15525_/CLK _15511_/D vssd1 vssd1 vccd1 vccd1 _15511_/Q sky130_fd_sc_hd__dfxtp_1
X_12723_ _15352_/Q _15351_/Q _12723_/C vssd1 vssd1 vccd1 vccd1 _12732_/B sky130_fd_sc_hd__and3_2
XFILLER_167_1083 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15442_ _15628_/CLK _15442_/D vssd1 vssd1 vccd1 vccd1 _15442_/Q sky130_fd_sc_hd__dfxtp_1
X_12654_ _13419_/Q _12653_/X _12662_/S vssd1 vssd1 vccd1 vccd1 _12655_/B sky130_fd_sc_hd__mux2_1
XFILLER_130_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11605_ _11606_/A _11606_/C _11606_/B vssd1 vssd1 vccd1 vccd1 _11611_/B sky130_fd_sc_hd__o21a_1
X_12585_ _13969_/Q _13711_/Q _12591_/S vssd1 vssd1 vccd1 vccd1 _12586_/B sky130_fd_sc_hd__mux2_1
X_15373_ _15374_/CLK _15373_/D vssd1 vssd1 vccd1 vccd1 _15373_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11536_ _11536_/A _11536_/B _11536_/C _13214_/A vssd1 vssd1 vccd1 vccd1 _11537_/B
+ sky130_fd_sc_hd__and4_1
X_14324_ _15172_/CLK _14324_/D vssd1 vssd1 vccd1 vccd1 _14324_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_172_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_488 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14255_ _15199_/CLK _14255_/D vssd1 vssd1 vccd1 vccd1 _14255_/Q sky130_fd_sc_hd__dfxtp_1
X_11467_ _06769_/Y _11475_/B _11455_/B vssd1 vssd1 vccd1 vccd1 _11468_/B sky130_fd_sc_hd__a21boi_1
XFILLER_125_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13206_ _13233_/A _11500_/A _13214_/B vssd1 vssd1 vccd1 vccd1 _13206_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_143_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10418_ _11496_/A _10418_/B _13199_/B vssd1 vssd1 vccd1 vccd1 _10418_/Y sky130_fd_sc_hd__nand3b_1
XFILLER_87_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14186_ _15672_/CLK _14186_/D vssd1 vssd1 vccd1 vccd1 _14186_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_125_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11398_ _11399_/A _11399_/B vssd1 vssd1 vccd1 vccd1 _11421_/A sky130_fd_sc_hd__and2_1
XFILLER_180_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13137_ _15534_/Q _08400_/C _13138_/S vssd1 vssd1 vccd1 vccd1 _15534_/D sky130_fd_sc_hd__mux2_1
XFILLER_125_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10349_ _07197_/B _10481_/B _10348_/X vssd1 vssd1 vccd1 vccd1 _13251_/B sky130_fd_sc_hd__a21o_4
XFILLER_97_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_856 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13068_ _12969_/X _13104_/A2 _13104_/B1 _07408_/X vssd1 vssd1 vccd1 vccd1 _13068_/X
+ sky130_fd_sc_hd__a22o_1
X_12019_ _12002_/X _12003_/X _12594_/S vssd1 vssd1 vccd1 vccd1 _12019_/X sky130_fd_sc_hd__mux2_1
XFILLER_17_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_954 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07560_ _13451_/Q _07560_/B vssd1 vssd1 vccd1 vccd1 _07560_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07491_ _13678_/Q _07499_/A2 _07499_/B1 _14706_/Q _07490_/X vssd1 vssd1 vccd1 vccd1
+ _07491_/X sky130_fd_sc_hd__a221o_1
XFILLER_179_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09230_ _13955_/Q _13697_/Q _09230_/S vssd1 vssd1 vccd1 vccd1 _09230_/X sky130_fd_sc_hd__mux2_1
XFILLER_181_1047 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09161_ _09221_/A _09161_/B vssd1 vssd1 vccd1 vccd1 _09161_/X sky130_fd_sc_hd__or2_1
XFILLER_119_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08112_ _13654_/Q _10344_/S _08096_/X _08111_/X vssd1 vssd1 vccd1 vccd1 _13654_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_30_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09092_ _15117_/Q _15085_/Q _15658_/Q _13392_/Q _09190_/S _09429_/S1 vssd1 vssd1
+ vccd1 vccd1 _09092_/X sky130_fd_sc_hd__mux4_1
XFILLER_119_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08043_ _14736_/Q _13614_/Q _08072_/S vssd1 vssd1 vccd1 vccd1 _13614_/D sky130_fd_sc_hd__mux2_1
XFILLER_135_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09994_ _13110_/B2 _14353_/Q _09996_/S vssd1 vssd1 vccd1 vccd1 _14353_/D sky130_fd_sc_hd__mux2_1
XFILLER_135_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08945_ _15651_/Q _13385_/Q _09005_/S vssd1 vssd1 vccd1 vccd1 _08945_/X sky130_fd_sc_hd__mux2_1
XFILLER_85_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08876_ _13897_/Q _13341_/A0 _08880_/S vssd1 vssd1 vccd1 vccd1 _13897_/D sky130_fd_sc_hd__mux2_1
XTAP_3806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07827_ _07836_/D _07826_/Y _07830_/A vssd1 vssd1 vccd1 vccd1 _07827_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_28_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07758_ _07756_/Y _07765_/C _07777_/A vssd1 vssd1 vccd1 vccd1 _07758_/Y sky130_fd_sc_hd__o21ai_1
X_06709_ _13467_/Q vssd1 vssd1 vccd1 vccd1 _07621_/A sky130_fd_sc_hd__inv_2
XFILLER_13_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07689_ _14741_/Q _07676_/A _07688_/Y _07938_/C1 vssd1 vssd1 vccd1 vccd1 _13484_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_44_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09428_ _15133_/Q _15101_/Q _15674_/Q _13408_/Q _09190_/S _09429_/S1 vssd1 vssd1
+ vccd1 vccd1 _09428_/X sky130_fd_sc_hd__mux4_1
XFILLER_25_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09359_ _09511_/S1 _09357_/X _09358_/X vssd1 vssd1 vccd1 vccd1 _09359_/X sky130_fd_sc_hd__a21o_1
XFILLER_100_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12370_ _14539_/Q _14152_/Q _14184_/Q _14120_/Q _12518_/S _12521_/A vssd1 vssd1 vccd1
+ vccd1 _12370_/X sky130_fd_sc_hd__mux4_1
XFILLER_121_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11321_ _11344_/A _08339_/X _11320_/Y _11346_/A2 vssd1 vssd1 vccd1 vccd1 _11321_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_107_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14040_ _15295_/CLK _14040_/D vssd1 vssd1 vccd1 vccd1 _14040_/Q sky130_fd_sc_hd__dfxtp_1
X_11252_ _11252_/A _11252_/B vssd1 vssd1 vccd1 vccd1 _11252_/Y sky130_fd_sc_hd__nor2_1
XFILLER_109_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10203_ input28/X _14588_/Q _13284_/S vssd1 vssd1 vccd1 vccd1 _14588_/D sky130_fd_sc_hd__mux2_1
XFILLER_106_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11183_ _08233_/B _11114_/X _11170_/X vssd1 vssd1 vccd1 vccd1 _11183_/X sky130_fd_sc_hd__a21o_1
XFILLER_79_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10134_ _14519_/Q _13320_/A0 _10164_/S vssd1 vssd1 vccd1 vccd1 _14519_/D sky130_fd_sc_hd__mux2_1
XFILLER_79_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14942_ _15006_/CLK _14942_/D vssd1 vssd1 vccd1 vccd1 _14942_/Q sky130_fd_sc_hd__dfxtp_1
X_10065_ _10065_/A _11818_/A vssd1 vssd1 vccd1 vccd1 _10065_/Y sky130_fd_sc_hd__nor2_8
XFILLER_48_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_954 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14873_ _15591_/CLK _14873_/D vssd1 vssd1 vccd1 vccd1 _14873_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13824_ _15218_/CLK _13824_/D vssd1 vssd1 vccd1 vccd1 _13824_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_165_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10967_ _11025_/A _11521_/A vssd1 vssd1 vccd1 vccd1 _11258_/A sky130_fd_sc_hd__and2_1
XFILLER_50_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13755_ _14888_/CLK _13755_/D vssd1 vssd1 vccd1 vccd1 _13755_/Q sky130_fd_sc_hd__dfxtp_1
X_12706_ _13426_/Q _12705_/X _12728_/S vssd1 vssd1 vccd1 vccd1 _12707_/B sky130_fd_sc_hd__mux2_1
X_13686_ _15278_/CLK _13686_/D vssd1 vssd1 vccd1 vccd1 _13686_/Q sky130_fd_sc_hd__dfxtp_1
X_10898_ _13162_/B _10951_/B vssd1 vssd1 vccd1 vccd1 _10898_/Y sky130_fd_sc_hd__nand2_1
X_15425_ _15623_/CLK _15425_/D vssd1 vssd1 vccd1 vccd1 _15425_/Q sky130_fd_sc_hd__dfxtp_2
X_12637_ _12644_/B _12637_/B vssd1 vssd1 vccd1 vccd1 _12637_/Y sky130_fd_sc_hd__nor2_1
XFILLER_12_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15356_ _15636_/CLK _15356_/D vssd1 vssd1 vccd1 vccd1 _15356_/Q sky130_fd_sc_hd__dfxtp_2
X_12568_ _14096_/Q _14064_/Q _12568_/S vssd1 vssd1 vccd1 vccd1 _12568_/X sky130_fd_sc_hd__mux2_1
XFILLER_172_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11519_ _11536_/C _11519_/B vssd1 vssd1 vccd1 vccd1 _11521_/B sky130_fd_sc_hd__xnor2_1
XFILLER_7_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14307_ _15306_/CLK _14307_/D vssd1 vssd1 vccd1 vccd1 _14307_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12499_ _14093_/Q _14061_/Q _12499_/S vssd1 vssd1 vccd1 vccd1 _12499_/X sky130_fd_sc_hd__mux2_1
X_15287_ _15287_/CLK _15287_/D vssd1 vssd1 vccd1 vccd1 _15287_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_171_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14238_ _15235_/CLK _14238_/D vssd1 vssd1 vccd1 vccd1 _14238_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14169_ _14462_/CLK _14169_/D vssd1 vssd1 vccd1 vccd1 _14169_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06991_ _13138_/S _06991_/B vssd1 vssd1 vccd1 vccd1 _06991_/X sky130_fd_sc_hd__and2_1
XFILLER_98_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08730_ _13577_/Q _08668_/X _08729_/X _13154_/S vssd1 vssd1 vccd1 vccd1 _08730_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08661_ _13521_/Q _08683_/A2 _08685_/A2 _13553_/Q vssd1 vssd1 vccd1 vccd1 _08661_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_27_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07612_ _14753_/Q _07607_/A _07611_/Y _07987_/C1 vssd1 vssd1 vccd1 vccd1 _13464_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_54_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08592_ _13783_/Q _08591_/X _08626_/S vssd1 vssd1 vccd1 vccd1 _13783_/D sky130_fd_sc_hd__mux2_1
XFILLER_82_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07543_ _14735_/Q _07644_/A _07542_/Y _08084_/C1 vssd1 vssd1 vccd1 vccd1 _13446_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_53_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07474_ _14670_/Q _07474_/B _07482_/C vssd1 vssd1 vccd1 vccd1 _07474_/X sky130_fd_sc_hd__and3_1
X_09213_ _14533_/Q _14146_/Q _14178_/Q _14114_/Q _09441_/S _09446_/A1 vssd1 vssd1
+ vccd1 vccd1 _09213_/X sky130_fd_sc_hd__mux4_1
XFILLER_33_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09144_ _14466_/Q _09536_/A2 _08520_/B _09143_/X vssd1 vssd1 vccd1 vccd1 _09144_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_182_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09075_ _09421_/A1 _09072_/X _09074_/X vssd1 vssd1 vccd1 vccd1 _09075_/X sky130_fd_sc_hd__a21o_1
X_08026_ _08027_/A _08033_/B vssd1 vssd1 vccd1 vccd1 _08028_/B sky130_fd_sc_hd__nor2_1
XFILLER_123_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_523 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09977_ _13331_/A0 _14336_/Q _09991_/S vssd1 vssd1 vccd1 vccd1 _14336_/D sky130_fd_sc_hd__mux2_1
XFILLER_77_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08928_ _14358_/Q _15174_/Q _13813_/Q _14552_/Q _09484_/S _08519_/A vssd1 vssd1 vccd1
+ vccd1 _08929_/B sky130_fd_sc_hd__mux4_1
XFILLER_40_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08859_ _13880_/Q _11649_/A0 _08885_/S vssd1 vssd1 vccd1 vccd1 _13880_/D sky130_fd_sc_hd__mux2_1
XFILLER_84_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11870_ _15291_/Q _11870_/A1 _11883_/S vssd1 vssd1 vccd1 vccd1 _15291_/D sky130_fd_sc_hd__mux2_1
XTAP_3669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10821_ _14853_/Q _07233_/A _12906_/S vssd1 vssd1 vccd1 vccd1 _14853_/D sky130_fd_sc_hd__mux2_1
XTAP_2957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_1023 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_1083 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_5_23_0_clk clkbuf_5_23_0_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_5_23_0_clk/X
+ sky130_fd_sc_hd__clkbuf_8
X_10752_ _15416_/Q _14784_/Q _10765_/S vssd1 vssd1 vccd1 vccd1 _14784_/D sky130_fd_sc_hd__mux2_1
X_13540_ _14517_/CLK _13540_/D vssd1 vssd1 vccd1 vccd1 _13540_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_1078 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13471_ _14513_/CLK _13471_/D vssd1 vssd1 vccd1 vccd1 _13471_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_9_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10683_ _15032_/Q _10652_/B _10682_/X vssd1 vssd1 vccd1 vccd1 _10683_/X sky130_fd_sc_hd__a21o_1
XFILLER_41_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12422_ _06670_/A _12419_/X _06671_/A vssd1 vssd1 vccd1 vccd1 _12422_/X sky130_fd_sc_hd__o21a_1
XFILLER_71_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15210_ _15676_/CLK _15210_/D vssd1 vssd1 vccd1 vccd1 _15210_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_185_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12353_ _12615_/B1 _12350_/X _12616_/C1 vssd1 vssd1 vccd1 vccd1 _12353_/X sky130_fd_sc_hd__o21a_1
X_15141_ _15676_/CLK _15141_/D vssd1 vssd1 vccd1 vccd1 _15141_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_153_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11304_ _11037_/A _13226_/B _10958_/B vssd1 vssd1 vccd1 vccd1 _11304_/Y sky130_fd_sc_hd__a21oi_2
X_15072_ _15581_/CLK _15072_/D vssd1 vssd1 vccd1 vccd1 _15072_/Q sky130_fd_sc_hd__dfxtp_4
X_12284_ _06670_/A _12281_/X _06671_/A vssd1 vssd1 vccd1 vccd1 _12284_/X sky130_fd_sc_hd__o21a_1
XFILLER_141_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14023_ _15292_/CLK _14023_/D vssd1 vssd1 vccd1 vccd1 _14023_/Q sky130_fd_sc_hd__dfxtp_1
X_11235_ _10471_/C _15023_/Q _11237_/S vssd1 vssd1 vccd1 vccd1 _15023_/D sky130_fd_sc_hd__mux2_1
XFILLER_171_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11166_ _11298_/A _11047_/B _11088_/S _11356_/C _13251_/A vssd1 vssd1 vccd1 vccd1
+ _11389_/B sky130_fd_sc_hd__a41o_4
X_10117_ _14503_/Q _14751_/Q _10124_/S vssd1 vssd1 vccd1 vccd1 _14503_/D sky130_fd_sc_hd__mux2_1
XFILLER_95_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11097_ _11371_/A _11093_/X _11096_/X vssd1 vssd1 vccd1 vccd1 _11179_/B sky130_fd_sc_hd__o21ai_4
XFILLER_67_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10048_ _14405_/Q _13082_/B2 _10059_/S vssd1 vssd1 vccd1 vccd1 _14405_/D sky130_fd_sc_hd__mux2_1
X_14925_ _15529_/CLK _14925_/D vssd1 vssd1 vccd1 vccd1 _14925_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14856_ _15519_/CLK _14856_/D vssd1 vssd1 vccd1 vccd1 _14856_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_136 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1071 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13807_ _15489_/CLK _13807_/D vssd1 vssd1 vccd1 vccd1 _13807_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14787_ _15638_/CLK _14787_/D vssd1 vssd1 vccd1 vccd1 _14787_/Q sky130_fd_sc_hd__dfxtp_1
X_11999_ _15310_/Q _10834_/S _11998_/X vssd1 vssd1 vccd1 vccd1 _15310_/D sky130_fd_sc_hd__a21o_1
XFILLER_90_275 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13738_ _15540_/CLK _13738_/D vssd1 vssd1 vccd1 vccd1 _13738_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_528 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13669_ _15645_/CLK _13669_/D vssd1 vssd1 vccd1 vccd1 _13669_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15408_ _15626_/CLK _15408_/D vssd1 vssd1 vccd1 vccd1 _15408_/Q sky130_fd_sc_hd__dfxtp_2
X_07190_ _15364_/Q _15071_/Q _07193_/S vssd1 vssd1 vccd1 vccd1 _07190_/X sky130_fd_sc_hd__mux2_8
XFILLER_157_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15339_ _15619_/CLK _15339_/D vssd1 vssd1 vccd1 vccd1 _15339_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_145_756 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09900_ _11853_/A1 _14261_/Q _09930_/S vssd1 vssd1 vccd1 vccd1 _14261_/D sky130_fd_sc_hd__mux2_1
XFILLER_116_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout506 _07490_/B vssd1 vssd1 vccd1 vccd1 _07474_/B sky130_fd_sc_hd__buf_6
XFILLER_63_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09831_ _11710_/A _10065_/A vssd1 vssd1 vccd1 vccd1 _09831_/Y sky130_fd_sc_hd__nor2_8
Xfanout517 _09554_/A vssd1 vssd1 vccd1 vccd1 _09382_/A sky130_fd_sc_hd__buf_12
XFILLER_99_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout528 _08487_/A vssd1 vssd1 vccd1 vccd1 _08988_/A1 sky130_fd_sc_hd__clkbuf_16
XFILLER_112_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout539 _08487_/A vssd1 vssd1 vccd1 vccd1 _09553_/A1 sky130_fd_sc_hd__clkbuf_16
XFILLER_59_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06974_ _06974_/A _06974_/B _06973_/X vssd1 vssd1 vccd1 vccd1 _06974_/X sky130_fd_sc_hd__or3b_2
XFILLER_140_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09762_ _14130_/Q _11883_/A1 _09762_/S vssd1 vssd1 vccd1 vccd1 _14130_/D sky130_fd_sc_hd__mux2_1
XTAP_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08713_ _15373_/Q _08748_/A2 _08736_/A2 _13418_/Q vssd1 vssd1 vccd1 vccd1 _08713_/X
+ sky130_fd_sc_hd__a22o_1
X_09693_ _14064_/Q _11881_/A1 _09695_/S vssd1 vssd1 vccd1 vccd1 _14064_/D sky130_fd_sc_hd__mux2_1
XFILLER_66_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08644_ _15383_/Q _08690_/A2 _08642_/X _08643_/X vssd1 vssd1 vccd1 vccd1 _08645_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_26_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08575_ _13605_/Q _08749_/A2 _08685_/A2 _13566_/Q _08574_/X vssd1 vssd1 vccd1 vccd1
+ _08579_/B sky130_fd_sc_hd__a221o_1
XFILLER_25_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_155_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07526_ _14756_/Q _13435_/Q _07529_/S vssd1 vssd1 vccd1 vccd1 _13435_/D sky130_fd_sc_hd__mux2_1
XFILLER_23_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07457_ _13339_/A0 _13403_/Q _07501_/S vssd1 vssd1 vccd1 vccd1 _13403_/D sky130_fd_sc_hd__mux2_1
XFILLER_183_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07388_ _14737_/Q _07387_/X _07500_/S vssd1 vssd1 vccd1 vccd1 _07388_/X sky130_fd_sc_hd__mux2_8
XFILLER_6_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09127_ _14014_/Q _13982_/Q _09230_/S vssd1 vssd1 vccd1 vccd1 _09127_/X sky130_fd_sc_hd__mux2_1
XFILLER_41_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09058_ _09530_/S1 _09056_/X _09057_/X vssd1 vssd1 vccd1 vccd1 _09062_/B sky130_fd_sc_hd__a21o_1
XFILLER_151_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08009_ _14761_/Q _08012_/A2 _08008_/Y _08016_/C1 vssd1 vssd1 vccd1 vccd1 _13568_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_104_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11020_ _11020_/A _11249_/A vssd1 vssd1 vccd1 vccd1 _11020_/Y sky130_fd_sc_hd__nor2_1
XFILLER_173_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12971_ _15470_/Q _13119_/S _13025_/B1 _12970_/X vssd1 vssd1 vccd1 vccd1 _15470_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_57_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14710_ _15646_/CLK _14710_/D vssd1 vssd1 vccd1 vccd1 _14710_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_3444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11922_ _14004_/Q _13972_/Q _12614_/S vssd1 vssd1 vccd1 vccd1 _11923_/B sky130_fd_sc_hd__mux2_1
XTAP_3455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1096 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_916 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14641_ _15647_/CLK _14641_/D vssd1 vssd1 vccd1 vccd1 _14641_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11853_ _15274_/Q _11853_/A1 _11883_/S vssd1 vssd1 vccd1 vccd1 _15274_/D sky130_fd_sc_hd__mux2_1
XTAP_2754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10804_ _14836_/Q _07312_/X _10871_/S vssd1 vssd1 vccd1 vccd1 _14836_/D sky130_fd_sc_hd__mux2_1
X_14572_ _14572_/CLK _14572_/D vssd1 vssd1 vccd1 vccd1 _14572_/Q sky130_fd_sc_hd__dfxtp_1
X_11784_ _15208_/Q _10892_/B _11781_/A _13808_/Q vssd1 vssd1 vccd1 vccd1 _15208_/D
+ sky130_fd_sc_hd__a22o_1
XTAP_2798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13523_ _15381_/CLK _13523_/D vssd1 vssd1 vccd1 vccd1 _13523_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_185_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10735_ _14765_/Q _10734_/X _10735_/S vssd1 vssd1 vccd1 vccd1 _14765_/D sky130_fd_sc_hd__mux2_1
XFILLER_186_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_695 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10666_ _15571_/Q _10706_/B vssd1 vssd1 vccd1 vccd1 _10666_/X sky130_fd_sc_hd__and2_1
X_13454_ _15377_/CLK _13454_/D vssd1 vssd1 vccd1 vccd1 _13454_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_139_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12405_ _14025_/Q _13993_/Q _12407_/S vssd1 vssd1 vccd1 vccd1 _12406_/B sky130_fd_sc_hd__mux2_1
XFILLER_139_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13385_ _15651_/CLK _13385_/D vssd1 vssd1 vccd1 vccd1 _13385_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_126_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10597_ _15557_/Q _10731_/B _10733_/B1 _14934_/Q vssd1 vssd1 vccd1 vccd1 _10597_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_12_1059 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15124_ _15665_/CLK _15124_/D vssd1 vssd1 vccd1 vccd1 _15124_/Q sky130_fd_sc_hd__dfxtp_1
X_12336_ _14022_/Q _13990_/Q _12543_/S vssd1 vssd1 vccd1 vccd1 _12337_/B sky130_fd_sc_hd__mux2_1
XFILLER_5_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15055_ _15569_/CLK _15055_/D vssd1 vssd1 vccd1 vccd1 _15055_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_141_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12267_ _14019_/Q _13987_/Q _12269_/S vssd1 vssd1 vccd1 vccd1 _12268_/B sky130_fd_sc_hd__mux2_1
X_11218_ _15007_/Q _11232_/S vssd1 vssd1 vccd1 vccd1 _11218_/Y sky130_fd_sc_hd__nand2b_1
X_14006_ _14462_/CLK _14006_/D vssd1 vssd1 vccd1 vccd1 _14006_/Q sky130_fd_sc_hd__dfxtp_1
X_12198_ _14016_/Q _13984_/Q _12476_/S vssd1 vssd1 vccd1 vccd1 _12199_/B sky130_fd_sc_hd__mux2_1
XFILLER_96_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput80 _07143_/X vssd1 vssd1 vccd1 vccd1 ext_write_data[21] sky130_fd_sc_hd__clkbuf_2
Xoutput91 _07163_/X vssd1 vssd1 vccd1 vccd1 ext_write_data[31] sky130_fd_sc_hd__clkbuf_2
X_11149_ _14973_/Q _10984_/Y _11146_/Y _11148_/Y vssd1 vssd1 vccd1 vccd1 _14973_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_23_1100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14908_ _15499_/CLK _14908_/D vssd1 vssd1 vccd1 vccd1 _14908_/Q sky130_fd_sc_hd__dfxtp_2
X_06690_ _15398_/Q vssd1 vssd1 vccd1 vccd1 _06690_/Y sky130_fd_sc_hd__inv_2
XFILLER_64_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14839_ _15508_/CLK _14839_/D vssd1 vssd1 vccd1 vccd1 _14839_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_45_990 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08360_ _13725_/Q _11346_/A2 _11351_/C1 _08359_/X vssd1 vssd1 vccd1 vccd1 _13725_/D
+ sky130_fd_sc_hd__a22o_1
X_07311_ _07348_/B _07310_/X _07350_/A vssd1 vssd1 vccd1 vccd1 _07311_/X sky130_fd_sc_hd__o21a_1
XFILLER_32_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08291_ _11298_/A _11351_/C1 _08290_/X _08232_/A _13718_/Q vssd1 vssd1 vccd1 vccd1
+ _13718_/D sky130_fd_sc_hd__a32o_1
XFILLER_108_1054 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07242_ _13928_/Q _15515_/Q _07334_/S vssd1 vssd1 vccd1 vccd1 _07242_/X sky130_fd_sc_hd__mux2_8
XFILLER_118_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07173_ _15347_/Q _15054_/Q _07188_/S vssd1 vssd1 vccd1 vccd1 _07173_/X sky130_fd_sc_hd__mux2_8
XFILLER_157_380 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1022 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout303 _13340_/A0 vssd1 vssd1 vccd1 vccd1 _11873_/A1 sky130_fd_sc_hd__buf_6
XFILLER_132_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout314 _07444_/X vssd1 vssd1 vccd1 vccd1 _13086_/B2 sky130_fd_sc_hd__clkbuf_8
XFILLER_99_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout325 _07420_/X vssd1 vssd1 vccd1 vccd1 _13330_/A0 sky130_fd_sc_hd__buf_6
XFILLER_98_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout336 _07400_/X vssd1 vssd1 vccd1 vccd1 _13325_/A0 sky130_fd_sc_hd__buf_6
X_09814_ _14180_/Q _13086_/B2 _09828_/S vssd1 vssd1 vccd1 vccd1 _14180_/D sky130_fd_sc_hd__mux2_1
Xfanout347 _07380_/X vssd1 vssd1 vccd1 vccd1 _13320_/A0 sky130_fd_sc_hd__buf_6
Xfanout358 _10732_/C1 vssd1 vssd1 vccd1 vccd1 _10717_/C1 sky130_fd_sc_hd__clkbuf_16
XFILLER_98_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout369 _08668_/D vssd1 vssd1 vccd1 vccd1 _08510_/B sky130_fd_sc_hd__buf_12
X_09745_ _14113_/Q _13333_/A0 _09757_/S vssd1 vssd1 vccd1 vccd1 _14113_/D sky130_fd_sc_hd__mux2_1
X_06957_ _06941_/C _06956_/Y _06944_/B vssd1 vssd1 vccd1 vccd1 _06957_/X sky130_fd_sc_hd__a21o_1
XFILLER_39_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06888_ _06888_/A _06929_/B vssd1 vssd1 vccd1 vccd1 _06888_/Y sky130_fd_sc_hd__nand2_1
XFILLER_28_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09676_ _14047_/Q _11689_/A0 _09690_/S vssd1 vssd1 vccd1 vccd1 _14047_/D sky130_fd_sc_hd__mux2_1
XTAP_2017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08627_ _13462_/Q _08684_/A2 _08683_/A2 _13526_/Q vssd1 vssd1 vccd1 vccd1 _08627_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_1305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08558_ _14514_/Q _08748_/B1 _08556_/X _08557_/X vssd1 vssd1 vccd1 vccd1 _08559_/C
+ sky130_fd_sc_hd__a211o_1
X_07509_ _14739_/Q _13418_/Q _07535_/S vssd1 vssd1 vccd1 vccd1 _13418_/D sky130_fd_sc_hd__mux2_1
XFILLER_23_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08489_ _13773_/Q _08488_/X _12481_/A vssd1 vssd1 vccd1 vccd1 _13773_/D sky130_fd_sc_hd__mux2_1
XFILLER_168_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10520_ _10520_/A1 _13787_/Q _13755_/Q _10520_/B2 vssd1 vssd1 vccd1 vccd1 _10520_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_167_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10451_ _08244_/A _13750_/Q _15422_/Q _08244_/B vssd1 vssd1 vccd1 vccd1 _10451_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_6_327 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13170_ _15557_/Q _13252_/B _13168_/Y _13169_/X vssd1 vssd1 vccd1 vccd1 _15557_/D
+ sky130_fd_sc_hd__a22o_1
X_10382_ _10382_/A _10382_/B _10382_/C _10382_/D vssd1 vssd1 vccd1 vccd1 _10390_/A
+ sky130_fd_sc_hd__or4_1
XFILLER_136_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12121_ _15283_/Q _15251_/Q _15219_/Q _15150_/Q _12489_/S0 _12489_/S1 vssd1 vssd1
+ vccd1 vccd1 _12122_/B sky130_fd_sc_hd__mux4_1
XFILLER_123_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12052_ _15280_/Q _15248_/Q _15216_/Q _15147_/Q _12154_/S _12253_/S1 vssd1 vssd1
+ vccd1 vccd1 _12053_/B sky130_fd_sc_hd__mux4_1
XFILLER_151_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_910 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11003_ _10982_/X _11002_/X _11414_/A vssd1 vssd1 vccd1 vccd1 _11003_/X sky130_fd_sc_hd__mux2_1
XFILLER_77_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12954_ _10594_/X _14865_/Q _13038_/S vssd1 vssd1 vccd1 vccd1 _12954_/X sky130_fd_sc_hd__mux2_2
XFILLER_46_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11905_ _12273_/A1 _11904_/X _11903_/X _12503_/C1 vssd1 vssd1 vccd1 vccd1 _11906_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_93_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15673_ _15673_/CLK _15673_/D vssd1 vssd1 vccd1 vccd1 _15673_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12885_ _15413_/Q _15598_/Q _12885_/S vssd1 vssd1 vccd1 vccd1 _15413_/D sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_193_clk clkbuf_5_20_0_clk/X vssd1 vssd1 vccd1 vccd1 _14537_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_18_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14624_ _15596_/CLK _14624_/D vssd1 vssd1 vccd1 vccd1 _14624_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11836_ _15258_/Q _13336_/A0 _11850_/S vssd1 vssd1 vccd1 vccd1 _15258_/D sky130_fd_sc_hd__mux2_1
XTAP_2584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14555_ _15278_/CLK _14555_/D vssd1 vssd1 vccd1 vccd1 _14555_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_122 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11767_ _13098_/B2 _15195_/Q _11775_/S vssd1 vssd1 vccd1 vccd1 _15195_/D sky130_fd_sc_hd__mux2_1
XTAP_1894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13506_ _13569_/CLK _13506_/D vssd1 vssd1 vccd1 vccd1 _13506_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_186_464 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10718_ _14990_/Q _10718_/A2 _10722_/B1 _14958_/Q _10717_/X vssd1 vssd1 vccd1 vccd1
+ _10718_/X sky130_fd_sc_hd__a221o_2
X_14486_ _15543_/CLK _14486_/D vssd1 vssd1 vccd1 vccd1 _14486_/Q sky130_fd_sc_hd__dfxtp_1
X_11698_ _11873_/A1 _15129_/Q _11708_/S vssd1 vssd1 vccd1 vccd1 _15129_/D sky130_fd_sc_hd__mux2_1
X_13437_ _15393_/CLK _13437_/D vssd1 vssd1 vccd1 vccd1 _13437_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_339 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10649_ _15057_/Q _10734_/A2 _10646_/X _10648_/X vssd1 vssd1 vccd1 vccd1 _10649_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_155_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13368_ _14471_/Q vssd1 vssd1 vccd1 vccd1 _14471_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_155_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15107_ _15680_/CLK _15107_/D vssd1 vssd1 vccd1 vccd1 _15107_/Q sky130_fd_sc_hd__dfxtp_1
X_12319_ _12595_/A1 _12318_/X _12317_/X _12618_/C1 vssd1 vssd1 vccd1 vccd1 _12320_/C
+ sky130_fd_sc_hd__a211o_1
X_13299_ _12717_/X _15631_/Q _13300_/S vssd1 vssd1 vccd1 vccd1 _15631_/D sky130_fd_sc_hd__mux2_1
XFILLER_5_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15038_ _15041_/CLK _15038_/D vssd1 vssd1 vccd1 vccd1 _15038_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_142_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07860_ _07869_/D _07859_/Y _07874_/A vssd1 vssd1 vccd1 vccd1 _07860_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_3_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06811_ _06663_/Y _08910_/S _13123_/A _13731_/Q vssd1 vssd1 vccd1 vccd1 _06811_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_68_378 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07791_ _13511_/Q _07802_/C vssd1 vssd1 vccd1 vccd1 _07792_/B sky130_fd_sc_hd__xnor2_1
XFILLER_77_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09530_ _15303_/Q _15271_/Q _15239_/Q _15170_/Q _09047_/S _09530_/S1 vssd1 vssd1
+ vccd1 vccd1 _09530_/X sky130_fd_sc_hd__mux4_1
XFILLER_97_1020 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06742_ _14491_/Q vssd1 vssd1 vccd1 vccd1 _06742_/Y sky130_fd_sc_hd__inv_2
XFILLER_36_220 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09461_ _15135_/Q _15103_/Q _15676_/Q _13410_/Q _09469_/S _09546_/S1 vssd1 vssd1
+ vccd1 vccd1 _09461_/X sky130_fd_sc_hd__mux4_1
X_06673_ _08910_/S vssd1 vssd1 vccd1 vccd1 _08668_/C sky130_fd_sc_hd__inv_6
Xclkbuf_leaf_184_clk clkbuf_5_21_0_clk/X vssd1 vssd1 vccd1 vccd1 _15200_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_92_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_1048 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08412_ _14613_/Q _08390_/A _08411_/X _13120_/S vssd1 vssd1 vccd1 vccd1 _08412_/X
+ sky130_fd_sc_hd__a31o_1
X_09392_ _15297_/Q _15265_/Q _15233_/Q _15164_/Q _09047_/S _09406_/S1 vssd1 vssd1
+ vccd1 vccd1 _09392_/X sky130_fd_sc_hd__mux4_1
XFILLER_52_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08343_ _07298_/X _10523_/A2 _08342_/X vssd1 vssd1 vccd1 vccd1 _11449_/A sky130_fd_sc_hd__a21oi_4
XFILLER_33_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08274_ _08258_/Y _08273_/X _11088_/S vssd1 vssd1 vccd1 vccd1 _08274_/X sky130_fd_sc_hd__mux2_4
XFILLER_165_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07225_ _07225_/A vssd1 vssd1 vccd1 vccd1 _07227_/B sky130_fd_sc_hd__inv_2
XFILLER_20_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_542 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07156_ _14858_/Q _14850_/Q _14842_/Q _14834_/Q _08094_/S _07104_/C vssd1 vssd1 vccd1
+ vccd1 _07157_/B sky130_fd_sc_hd__mux4_1
XFILLER_161_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07087_ _14641_/Q _14673_/Q _07096_/S vssd1 vssd1 vccd1 vccd1 _07087_/X sky130_fd_sc_hd__mux2_1
XFILLER_154_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout111 _13288_/S vssd1 vssd1 vccd1 vccd1 _13309_/A sky130_fd_sc_hd__buf_12
Xfanout122 _10834_/S vssd1 vssd1 vccd1 vccd1 _13105_/A2 sky130_fd_sc_hd__buf_8
Xfanout133 fanout138/X vssd1 vssd1 vccd1 vccd1 _10892_/B sky130_fd_sc_hd__buf_6
Xfanout144 _12320_/A vssd1 vssd1 vccd1 vccd1 _12596_/A sky130_fd_sc_hd__buf_12
XFILLER_59_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout155 _12885_/S vssd1 vssd1 vccd1 vccd1 _12927_/S sky130_fd_sc_hd__buf_12
XFILLER_87_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout166 _12839_/X vssd1 vssd1 vccd1 vccd1 _12871_/S sky130_fd_sc_hd__buf_12
Xfanout177 _11676_/X vssd1 vssd1 vccd1 vccd1 _11703_/S sky130_fd_sc_hd__buf_12
Xfanout188 _10032_/Y vssd1 vssd1 vccd1 vccd1 _10064_/S sky130_fd_sc_hd__buf_12
XFILLER_86_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_14 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout199 _09796_/Y vssd1 vssd1 vccd1 vccd1 _09823_/S sky130_fd_sc_hd__buf_12
X_07989_ _13563_/Q _07995_/D vssd1 vssd1 vccd1 vccd1 _07989_/X sky130_fd_sc_hd__or2_1
XFILLER_47_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_68 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09728_ _11883_/A1 _14098_/Q _09728_/S vssd1 vssd1 vccd1 vccd1 _14098_/D sky130_fd_sc_hd__mux2_1
XFILLER_83_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09659_ _14032_/Q _11881_/A1 _09661_/S vssd1 vssd1 vccd1 vccd1 _14032_/D sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_175_clk clkbuf_5_23_0_clk/X vssd1 vssd1 vccd1 vccd1 _15301_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12670_ _13421_/Q _12669_/X _12764_/S vssd1 vssd1 vccd1 vccd1 _12671_/B sky130_fd_sc_hd__mux2_1
XTAP_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11621_ _11621_/A _11621_/B vssd1 vssd1 vccd1 vccd1 _11621_/X sky130_fd_sc_hd__xor2_1
XFILLER_30_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14340_ _15289_/CLK _14340_/D vssd1 vssd1 vccd1 vccd1 _14340_/Q sky130_fd_sc_hd__dfxtp_1
X_11552_ _11569_/B _11552_/B vssd1 vssd1 vccd1 vccd1 _11555_/B sky130_fd_sc_hd__xor2_2
XFILLER_184_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10503_ _11569_/B _13220_/B vssd1 vssd1 vccd1 vccd1 _10542_/A sky130_fd_sc_hd__or2_1
XFILLER_128_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11483_ _11472_/B _11505_/B _11482_/X vssd1 vssd1 vccd1 vccd1 _11484_/B sky130_fd_sc_hd__a21o_1
X_14271_ _15181_/CLK _14271_/D vssd1 vssd1 vccd1 vccd1 _14271_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_155_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13222_ _13220_/Y _13221_/X _15574_/Q _13214_/B vssd1 vssd1 vccd1 vccd1 _15574_/D
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_10_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10434_ _07204_/A _10523_/A2 _10433_/X vssd1 vssd1 vccd1 vccd1 _13242_/B sky130_fd_sc_hd__a21o_4
XFILLER_12_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10365_ _10418_/B _10365_/B vssd1 vssd1 vccd1 vccd1 _10366_/C sky130_fd_sc_hd__nand2_1
XFILLER_152_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13153_ _14613_/Q _15551_/Q _13154_/S vssd1 vssd1 vccd1 vccd1 _15551_/D sky130_fd_sc_hd__mux2_1
XFILLER_151_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12104_ _13884_/Q _14399_/Q _12476_/S vssd1 vssd1 vccd1 vccd1 _12104_/X sky130_fd_sc_hd__mux2_1
X_13084_ _12993_/X _13104_/A2 _13104_/B1 _07440_/X vssd1 vssd1 vccd1 vccd1 _13084_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10296_ _14681_/Q _14866_/Q _10615_/S vssd1 vssd1 vccd1 vccd1 _14681_/D sky130_fd_sc_hd__mux2_1
XFILLER_124_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12035_ _13881_/Q _14396_/Q _12591_/S vssd1 vssd1 vccd1 vccd1 _12035_/X sky130_fd_sc_hd__mux2_1
XFILLER_105_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13986_ _15088_/CLK _13986_/D vssd1 vssd1 vccd1 vccd1 _13986_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12937_ _10578_/X _14862_/Q _13038_/S vssd1 vssd1 vccd1 vccd1 _12937_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_166_clk clkbuf_5_22_0_clk/X vssd1 vssd1 vccd1 vccd1 _15676_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_3071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15656_ _15656_/CLK _15656_/D vssd1 vssd1 vccd1 vccd1 _15656_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12868_ _14762_/Q _15396_/Q _12871_/S vssd1 vssd1 vccd1 vccd1 _15396_/D sky130_fd_sc_hd__mux2_1
XFILLER_178_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14607_ _15375_/CLK _14607_/D vssd1 vssd1 vccd1 vccd1 _14607_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_33_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11819_ _15241_/Q _11852_/A1 _11849_/S vssd1 vssd1 vccd1 vccd1 _15241_/D sky130_fd_sc_hd__mux2_1
XTAP_1680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15587_ _15587_/CLK _15587_/D vssd1 vssd1 vccd1 vccd1 _15587_/Q sky130_fd_sc_hd__dfxtp_1
X_12799_ _12828_/A _12799_/B vssd1 vssd1 vccd1 vccd1 _12799_/X sky130_fd_sc_hd__or2_1
XTAP_1691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14538_ _15669_/CLK _14538_/D vssd1 vssd1 vccd1 vccd1 _14538_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_175_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_1046 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14469_ _15664_/CLK _14469_/D vssd1 vssd1 vccd1 vccd1 _14469_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_162_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07010_ _07009_/X _13582_/Q _12662_/S vssd1 vssd1 vccd1 vccd1 _07010_/X sky130_fd_sc_hd__mux2_1
XFILLER_134_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08961_ _13878_/Q _09231_/A2 _09403_/B1 _14393_/Q _09445_/C1 vssd1 vssd1 vccd1 vccd1
+ _08961_/X sky130_fd_sc_hd__a221o_1
XFILLER_103_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07912_ _14735_/Q _08022_/B _07911_/Y _08016_/C1 vssd1 vssd1 vccd1 vccd1 _13542_/D
+ sky130_fd_sc_hd__o211a_1
X_08892_ _09449_/A1 _08890_/X _08891_/X _09449_/B2 _08889_/X vssd1 vssd1 vccd1 vccd1
+ _08892_/X sky130_fd_sc_hd__a221o_1
XFILLER_124_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07843_ _14749_/Q _07830_/A _07842_/X _07949_/C1 vssd1 vssd1 vccd1 vccd1 _13524_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_68_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07774_ _14764_/Q _07777_/A _07773_/Y _08016_/C1 vssd1 vssd1 vccd1 vccd1 _13507_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_84_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09513_ _15105_/Q _08540_/B _13130_/C1 _09512_/X vssd1 vssd1 vccd1 vccd1 _09513_/X
+ sky130_fd_sc_hd__a22o_1
X_06725_ _13459_/Q vssd1 vssd1 vccd1 vccd1 _07595_/B sky130_fd_sc_hd__inv_2
XFILLER_140_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_157_clk clkbuf_5_25_0_clk/X vssd1 vssd1 vccd1 vccd1 _15208_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_52_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09444_ _13965_/Q _13707_/Q _09444_/S vssd1 vssd1 vccd1 vccd1 _09444_/X sky130_fd_sc_hd__mux2_1
XPHY_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09375_ _08668_/D _09373_/X _09374_/X _08519_/B _13049_/A1 vssd1 vssd1 vccd1 vccd1
+ _09375_/X sky130_fd_sc_hd__a221o_1
XFILLER_178_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08326_ _11431_/A vssd1 vssd1 vccd1 vccd1 _13183_/B sky130_fd_sc_hd__inv_2
XFILLER_166_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08257_ _11349_/B _13159_/B _10551_/B vssd1 vssd1 vccd1 vccd1 _08259_/B sky130_fd_sc_hd__o21ai_4
XFILLER_20_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_3_5_0_clk clkbuf_3_5_0_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_5_0_clk/X sky130_fd_sc_hd__clkbuf_8
X_07208_ _07208_/A vssd1 vssd1 vccd1 vccd1 _07208_/Y sky130_fd_sc_hd__inv_2
XFILLER_137_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08188_ _14714_/Q _14715_/Q _14716_/Q _08817_/B vssd1 vssd1 vccd1 vccd1 _10032_/A
+ sky130_fd_sc_hd__nand4_4
XFILLER_119_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07139_ _14833_/Q _07104_/X _07138_/X _07131_/A vssd1 vssd1 vccd1 vccd1 _07139_/X
+ sky130_fd_sc_hd__a22o_4
XFILLER_3_138 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10150_ _14535_/Q _13086_/B2 _10164_/S vssd1 vssd1 vccd1 vccd1 _14535_/D sky130_fd_sc_hd__mux2_1
XFILLER_161_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10081_ _14437_/Q _13334_/A0 _10092_/S vssd1 vssd1 vccd1 vccd1 _14437_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13840_ _15335_/CLK _13840_/D vssd1 vssd1 vccd1 vccd1 _13840_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_74_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13771_ _15588_/CLK _13771_/D vssd1 vssd1 vccd1 vccd1 _13771_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_148_clk clkbuf_5_25_0_clk/X vssd1 vssd1 vccd1 vccd1 _13803_/CLK sky130_fd_sc_hd__clkbuf_16
X_10983_ _14928_/D _14927_/D _14929_/D vssd1 vssd1 vccd1 vccd1 _10983_/X sky130_fd_sc_hd__and3b_4
XFILLER_43_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15510_ _15510_/CLK _15510_/D vssd1 vssd1 vccd1 vccd1 _15510_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12722_ _15351_/Q _12765_/B _12721_/X _12809_/C1 vssd1 vssd1 vccd1 vccd1 _15351_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_167_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_1095 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15441_ _15632_/CLK _15441_/D vssd1 vssd1 vccd1 vccd1 _15441_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12653_ _13586_/Q _12652_/X _12785_/B vssd1 vssd1 vccd1 vccd1 _12653_/X sky130_fd_sc_hd__mux2_1
XFILLER_157_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11604_ _11604_/A _11604_/B vssd1 vssd1 vccd1 vccd1 _11606_/C sky130_fd_sc_hd__nor2_1
XFILLER_90_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15372_ _15372_/CLK _15372_/D vssd1 vssd1 vccd1 vccd1 _15372_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_168_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12584_ _12595_/A1 _12579_/X _12582_/X _12583_/X _08405_/D vssd1 vssd1 vccd1 vccd1
+ _12596_/B sky130_fd_sc_hd__a221o_1
XFILLER_7_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14323_ _15203_/CLK _14323_/D vssd1 vssd1 vccd1 vccd1 _14323_/Q sky130_fd_sc_hd__dfxtp_1
X_11535_ _11534_/Y _15062_/Q _11614_/S vssd1 vssd1 vccd1 vccd1 _15062_/D sky130_fd_sc_hd__mux2_1
XFILLER_11_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_967 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14254_ _15332_/CLK _14254_/D vssd1 vssd1 vccd1 vccd1 _14254_/Q sky130_fd_sc_hd__dfxtp_1
X_11466_ _15055_/Q _11474_/S _11465_/X vssd1 vssd1 vccd1 vccd1 _15055_/D sky130_fd_sc_hd__a21bo_1
XFILLER_172_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13205_ _13233_/A _11500_/A _11536_/B vssd1 vssd1 vccd1 vccd1 _13205_/X sky130_fd_sc_hd__o21ba_1
X_10417_ _10381_/A _10384_/A _10413_/X _10416_/X _10557_/A vssd1 vssd1 vccd1 vccd1
+ _10417_/X sky130_fd_sc_hd__a41o_1
X_14185_ _15679_/CLK _14185_/D vssd1 vssd1 vccd1 vccd1 _14185_/Q sky130_fd_sc_hd__dfxtp_1
X_11397_ _11414_/C _11397_/B vssd1 vssd1 vccd1 vccd1 _11399_/B sky130_fd_sc_hd__xnor2_1
XFILLER_125_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13136_ _15533_/Q _10892_/B _13129_/Y vssd1 vssd1 vccd1 vccd1 _15533_/D sky130_fd_sc_hd__a21o_1
XTAP_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10348_ _10507_/A1 _13743_/Q _15429_/Q _10515_/B2 vssd1 vssd1 vccd1 vccd1 _10348_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10279_ _14664_/Q _14817_/Q _10665_/S vssd1 vssd1 vccd1 vccd1 _14664_/D sky130_fd_sc_hd__mux2_1
XTAP_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13067_ _15501_/Q _13120_/S _13105_/B1 _13066_/X vssd1 vssd1 vccd1 vccd1 _15501_/D
+ sky130_fd_sc_hd__a22o_1
X_12018_ _12011_/X _12013_/X _12015_/X _12017_/X _06671_/A vssd1 vssd1 vccd1 vccd1
+ _12018_/X sky130_fd_sc_hd__o221a_1
XFILLER_94_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13969_ _15679_/CLK _13969_/D vssd1 vssd1 vccd1 vccd1 _13969_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_139_clk clkbuf_5_29_0_clk/X vssd1 vssd1 vccd1 vccd1 _15542_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_19_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07490_ _14674_/Q _07490_/B _07498_/C vssd1 vssd1 vccd1 vccd1 _07490_/X sky130_fd_sc_hd__and3_1
X_15639_ _15641_/CLK _15639_/D vssd1 vssd1 vccd1 vccd1 _15639_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_179_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09160_ _14369_/Q _15185_/Q _13824_/Q _14563_/Q _09190_/S _09429_/S1 vssd1 vssd1
+ vccd1 vccd1 _09161_/B sky130_fd_sc_hd__mux4_1
X_08111_ input28/X input5/X input14/X input22/X _08150_/S _08151_/S vssd1 vssd1 vccd1
+ vccd1 _08111_/X sky130_fd_sc_hd__mux4_1
X_09091_ _09429_/S1 _09089_/X _09090_/X vssd1 vssd1 vccd1 vccd1 _09091_/X sky130_fd_sc_hd__a21o_1
XFILLER_175_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08042_ _14735_/Q _13613_/Q _08072_/S vssd1 vssd1 vccd1 vccd1 _13613_/D sky130_fd_sc_hd__mux2_1
XFILLER_162_404 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09993_ _11847_/A1 _14352_/Q _09996_/S vssd1 vssd1 vccd1 vccd1 _14352_/D sky130_fd_sc_hd__mux2_1
XFILLER_142_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_548 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08944_ _14520_/Q _14133_/Q _14165_/Q _14101_/Q _09005_/S _09511_/S1 vssd1 vssd1
+ vccd1 vccd1 _08944_/X sky130_fd_sc_hd__mux4_1
XFILLER_130_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08875_ _13896_/Q _11873_/A1 _08885_/S vssd1 vssd1 vccd1 vccd1 _13896_/D sky130_fd_sc_hd__mux2_1
XFILLER_57_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07826_ _13519_/Q _13518_/Q _07825_/D _13520_/Q vssd1 vssd1 vccd1 vccd1 _07826_/Y
+ sky130_fd_sc_hd__a31oi_1
XTAP_3829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07757_ _13503_/Q _13502_/Q _13501_/Q _07757_/D vssd1 vssd1 vccd1 vccd1 _07765_/C
+ sky130_fd_sc_hd__and4_1
XFILLER_25_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06708_ _14508_/Q vssd1 vssd1 vccd1 vccd1 _06708_/Y sky130_fd_sc_hd__inv_2
XFILLER_53_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07688_ _07686_/Y _07717_/A _07676_/A vssd1 vssd1 vccd1 vccd1 _07688_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_52_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09427_ _09427_/A1 _09425_/X _09426_/X vssd1 vssd1 vccd1 vccd1 _09427_/X sky130_fd_sc_hd__a21o_1
XFILLER_12_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09358_ _14089_/Q _09522_/A2 _09519_/B1 _14057_/Q _09532_/A vssd1 vssd1 vccd1 vccd1
+ _09358_/X sky130_fd_sc_hd__a221o_1
XFILLER_8_208 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08309_ _11371_/A _08309_/B vssd1 vssd1 vccd1 vccd1 _08309_/Y sky130_fd_sc_hd__nor2_1
XFILLER_154_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09289_ _14441_/Q _08540_/B _08520_/B _09288_/X vssd1 vssd1 vccd1 vccd1 _09289_/X
+ sky130_fd_sc_hd__a22o_1
X_11320_ _11347_/A _11260_/X _11319_/X vssd1 vssd1 vccd1 vccd1 _11320_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_158_1006 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_990 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11251_ _11252_/B vssd1 vssd1 vccd1 vccd1 _11251_/Y sky130_fd_sc_hd__inv_2
XFILLER_181_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10202_ input27/X _14587_/Q _13284_/S vssd1 vssd1 vccd1 vccd1 _14587_/D sky130_fd_sc_hd__mux2_1
XFILLER_122_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11182_ _14983_/Q _11164_/S _11170_/X _11181_/Y vssd1 vssd1 vccd1 vccd1 _14983_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_69_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10133_ _14518_/Q _11852_/A1 _10159_/S vssd1 vssd1 vccd1 vccd1 _14518_/D sky130_fd_sc_hd__mux2_1
XFILLER_79_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14941_ _15580_/CLK _14941_/D vssd1 vssd1 vccd1 vccd1 _14941_/Q sky130_fd_sc_hd__dfxtp_1
X_10064_ _14421_/Q _13350_/A0 _10064_/S vssd1 vssd1 vccd1 vccd1 _14421_/D sky130_fd_sc_hd__mux2_1
XFILLER_88_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14872_ _15422_/CLK _14872_/D vssd1 vssd1 vccd1 vccd1 _14872_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_668 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13823_ _15184_/CLK _13823_/D vssd1 vssd1 vccd1 vccd1 _13823_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13754_ _14868_/CLK _13754_/D vssd1 vssd1 vccd1 vccd1 _13754_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_188_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10966_ _11025_/A _13215_/B vssd1 vssd1 vccd1 vccd1 _11272_/A sky130_fd_sc_hd__nor2_1
XFILLER_31_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_576 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12705_ _13593_/Q _12704_/X _12763_/S vssd1 vssd1 vccd1 vccd1 _12705_/X sky130_fd_sc_hd__mux2_1
XFILLER_71_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13685_ _15665_/CLK _13685_/D vssd1 vssd1 vccd1 vccd1 _13685_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10897_ _14931_/Q _10554_/A _10951_/B vssd1 vssd1 vccd1 vccd1 _14931_/D sky130_fd_sc_hd__mux2_1
XFILLER_176_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15424_ _15624_/CLK _15424_/D vssd1 vssd1 vccd1 vccd1 _15424_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_148_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12636_ _15339_/Q _15338_/Q _15340_/Q vssd1 vssd1 vccd1 vccd1 _12637_/B sky130_fd_sc_hd__a21oi_1
XFILLER_157_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_579 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15355_ _15635_/CLK _15355_/D vssd1 vssd1 vccd1 vccd1 _15355_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_156_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12567_ _12567_/A _12567_/B vssd1 vssd1 vccd1 vccd1 _12567_/X sky130_fd_sc_hd__and2_1
XFILLER_156_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14306_ _14468_/CLK _14306_/D vssd1 vssd1 vccd1 vccd1 _14306_/Q sky130_fd_sc_hd__dfxtp_1
X_11518_ _11536_/A _11536_/B _11537_/A _13236_/A vssd1 vssd1 vccd1 vccd1 _11519_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_117_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15286_ _15286_/CLK _15286_/D vssd1 vssd1 vccd1 vccd1 _15286_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12498_ _12498_/A _12498_/B vssd1 vssd1 vccd1 vccd1 _12498_/X sky130_fd_sc_hd__and2_1
XFILLER_172_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14237_ _15181_/CLK _14237_/D vssd1 vssd1 vccd1 vccd1 _14237_/Q sky130_fd_sc_hd__dfxtp_1
X_11449_ _11449_/A _11449_/B vssd1 vssd1 vccd1 vccd1 _11450_/B sky130_fd_sc_hd__or2_1
XFILLER_153_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14168_ _15081_/CLK _14168_/D vssd1 vssd1 vccd1 vccd1 _14168_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13119_ _14596_/Q _15528_/Q _13119_/S vssd1 vssd1 vccd1 vccd1 _15528_/D sky130_fd_sc_hd__mux2_1
XFILLER_98_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14099_ _15172_/CLK _14099_/D vssd1 vssd1 vccd1 vccd1 _14099_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06990_ _08773_/A _09829_/C vssd1 vssd1 vccd1 vccd1 _06991_/B sky130_fd_sc_hd__nor2_1
XTAP_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08660_ _13793_/Q _12917_/S _08659_/X vssd1 vssd1 vccd1 vccd1 _13793_/D sky130_fd_sc_hd__o21a_1
XFILLER_66_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07611_ _07609_/Y _07617_/C _07614_/A vssd1 vssd1 vccd1 vccd1 _07611_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_82_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08591_ _14509_/Q _08693_/A2 _08588_/X _08589_/X _08590_/X vssd1 vssd1 vccd1 vccd1
+ _08591_/X sky130_fd_sc_hd__a2111o_1
XFILLER_35_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07542_ _07644_/A _07542_/B vssd1 vssd1 vccd1 vccd1 _07542_/Y sky130_fd_sc_hd__nand2_1
XFILLER_50_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07473_ _13343_/A0 _13407_/Q _07481_/S vssd1 vssd1 vccd1 vccd1 _13407_/D sky130_fd_sc_hd__mux2_1
XFILLER_50_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09212_ _09405_/A _09212_/B _09212_/C vssd1 vssd1 vccd1 vccd1 _09212_/X sky130_fd_sc_hd__and3_1
XFILLER_33_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09143_ _13855_/Q _14208_/Q _09407_/S vssd1 vssd1 vccd1 vccd1 _09143_/X sky130_fd_sc_hd__mux2_1
XFILLER_147_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09074_ _14462_/Q _09536_/A2 _13130_/B1 _14430_/Q _06676_/A vssd1 vssd1 vccd1 vccd1
+ _09074_/X sky130_fd_sc_hd__a221o_1
XFILLER_135_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08025_ _14717_/Q _14718_/Q _08025_/C vssd1 vssd1 vccd1 vccd1 _08033_/B sky130_fd_sc_hd__or3_4
XFILLER_89_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_1050 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_25 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09976_ _13330_/A0 _14335_/Q _09991_/S vssd1 vssd1 vccd1 vccd1 _14335_/D sky130_fd_sc_hd__mux2_1
XFILLER_39_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08927_ _13908_/Q _13139_/S _08926_/X vssd1 vssd1 vccd1 vccd1 _13908_/D sky130_fd_sc_hd__a21o_1
XFILLER_103_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08858_ _13879_/Q _11681_/A0 _08880_/S vssd1 vssd1 vccd1 vccd1 _13879_/D sky130_fd_sc_hd__mux2_1
XFILLER_58_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07809_ _14740_/Q _07816_/A _07808_/X _07938_/C1 vssd1 vssd1 vccd1 vccd1 _13515_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_3659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08789_ _13323_/A0 _13815_/Q _08811_/S vssd1 vssd1 vccd1 vccd1 _13815_/D sky130_fd_sc_hd__mux2_1
XFILLER_55_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10820_ _14852_/Q _07237_/A _10868_/S vssd1 vssd1 vccd1 vccd1 _14852_/D sky130_fd_sc_hd__mux2_1
XTAP_2947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_351 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10751_ _15415_/Q _14783_/Q _10765_/S vssd1 vssd1 vccd1 vccd1 _14783_/D sky130_fd_sc_hd__mux2_1
XFILLER_77_1095 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13470_ _15393_/CLK _13470_/D vssd1 vssd1 vccd1 vccd1 _13470_/Q sky130_fd_sc_hd__dfxtp_2
X_10682_ _15574_/Q _10731_/B _10733_/B1 _14951_/Q vssd1 vssd1 vccd1 vccd1 _10682_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_40_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12421_ _12559_/A _12421_/B vssd1 vssd1 vccd1 vccd1 _12421_/X sky130_fd_sc_hd__or2_1
XFILLER_138_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15140_ _15209_/CLK _15140_/D vssd1 vssd1 vccd1 vccd1 _15140_/Q sky130_fd_sc_hd__dfxtp_1
X_12352_ _12536_/A _12352_/B vssd1 vssd1 vccd1 vccd1 _12352_/X sky130_fd_sc_hd__or2_1
XFILLER_126_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11303_ _11303_/A vssd1 vssd1 vccd1 vccd1 _11303_/Y sky130_fd_sc_hd__inv_2
XFILLER_154_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15071_ _15591_/CLK _15071_/D vssd1 vssd1 vccd1 vccd1 _15071_/Q sky130_fd_sc_hd__dfxtp_4
X_12283_ _12594_/S _12283_/B vssd1 vssd1 vccd1 vccd1 _12283_/X sky130_fd_sc_hd__or2_1
XFILLER_153_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14022_ _14537_/CLK _14022_/D vssd1 vssd1 vccd1 vccd1 _14022_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_107_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11234_ _10471_/B _15022_/Q _11237_/S vssd1 vssd1 vccd1 vccd1 _15022_/D sky130_fd_sc_hd__mux2_1
XFILLER_20_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_131 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11165_ _11122_/X _11124_/X _11298_/A vssd1 vssd1 vccd1 vccd1 _11165_/X sky130_fd_sc_hd__mux2_1
XFILLER_171_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10116_ _14502_/Q _14750_/Q _10124_/S vssd1 vssd1 vccd1 vccd1 _14502_/D sky130_fd_sc_hd__mux2_1
X_11096_ _11129_/A _11096_/B vssd1 vssd1 vccd1 vccd1 _11096_/X sky130_fd_sc_hd__or2_2
XFILLER_48_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10047_ _14404_/Q _13333_/A0 _10059_/S vssd1 vssd1 vccd1 vccd1 _14404_/D sky130_fd_sc_hd__mux2_1
X_14924_ _15648_/CLK _14924_/D vssd1 vssd1 vccd1 vccd1 _14924_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_64_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14855_ _15519_/CLK _14855_/D vssd1 vssd1 vccd1 vccd1 _14855_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13806_ _15462_/CLK _13806_/D vssd1 vssd1 vccd1 vccd1 _13806_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_1083 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14786_ _15637_/CLK _14786_/D vssd1 vssd1 vccd1 vccd1 _14786_/Q sky130_fd_sc_hd__dfxtp_1
X_11998_ _12596_/A _11998_/B _11998_/C vssd1 vssd1 vccd1 vccd1 _11998_/X sky130_fd_sc_hd__and3_2
XFILLER_90_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13737_ _15540_/CLK _13737_/D vssd1 vssd1 vccd1 vccd1 _13737_/Q sky130_fd_sc_hd__dfxtp_2
X_10949_ _14959_/Q _10948_/B _10948_/Y _11624_/A vssd1 vssd1 vccd1 vccd1 _14959_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_31_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_70_clk clkbuf_5_14_0_clk/X vssd1 vssd1 vccd1 vccd1 _15569_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_177_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13668_ _15606_/CLK _13668_/D vssd1 vssd1 vccd1 vccd1 _13668_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_188_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15407_ _15592_/CLK _15407_/D vssd1 vssd1 vccd1 vccd1 _15407_/Q sky130_fd_sc_hd__dfxtp_2
X_12619_ _13134_/A _12619_/B _12619_/C vssd1 vssd1 vccd1 vccd1 _12619_/X sky130_fd_sc_hd__and3_1
X_13599_ _15635_/CLK _13599_/D vssd1 vssd1 vccd1 vccd1 _13599_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_77_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15338_ _15429_/CLK _15338_/D vssd1 vssd1 vccd1 vccd1 _15338_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_129_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_768 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15269_ _15301_/CLK _15269_/D vssd1 vssd1 vccd1 vccd1 _15269_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_160_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout507 _07498_/B vssd1 vssd1 vccd1 vccd1 _07490_/B sky130_fd_sc_hd__buf_4
X_09830_ _10515_/B2 _13138_/S _09829_/X vssd1 vssd1 vccd1 vccd1 _14195_/D sky130_fd_sc_hd__o21a_1
XFILLER_112_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout518 _14606_/Q vssd1 vssd1 vccd1 vccd1 _09554_/A sky130_fd_sc_hd__buf_12
Xfanout529 _09530_/S1 vssd1 vssd1 vccd1 vccd1 _09234_/S1 sky130_fd_sc_hd__buf_12
XFILLER_98_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09761_ _14129_/Q _13349_/A0 _09762_/S vssd1 vssd1 vccd1 vccd1 _14129_/D sky130_fd_sc_hd__mux2_1
X_06973_ _06720_/Y _13493_/Q _06971_/X _06972_/X vssd1 vssd1 vccd1 vccd1 _06973_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08712_ _13450_/Q _08746_/A2 _08747_/B1 _13482_/Q _08711_/X vssd1 vssd1 vccd1 vccd1
+ _08712_/X sky130_fd_sc_hd__a221o_1
X_09692_ _14063_/Q _13347_/A0 _09695_/S vssd1 vssd1 vccd1 vccd1 _14063_/D sky130_fd_sc_hd__mux2_1
XFILLER_132_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08643_ _13556_/Q _08685_/A2 _08693_/B1 _13627_/Q vssd1 vssd1 vccd1 vccd1 _08643_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_54_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08574_ _13470_/Q _08746_/A2 _08750_/A2 _13534_/Q vssd1 vssd1 vccd1 vccd1 _08574_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_26_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07525_ _14755_/Q _13434_/Q _07529_/S vssd1 vssd1 vccd1 vccd1 _13434_/D sky130_fd_sc_hd__mux2_1
XFILLER_23_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_61_clk _15031_/CLK vssd1 vssd1 vccd1 vccd1 _15006_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_62_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07456_ _14754_/Q _07455_/X _07480_/S vssd1 vssd1 vccd1 vccd1 _07456_/X sky130_fd_sc_hd__mux2_4
XFILLER_22_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07387_ _13652_/Q _07499_/A2 _07499_/B1 _14680_/Q _07386_/X vssd1 vssd1 vccd1 vccd1
+ _07387_/X sky130_fd_sc_hd__a221o_1
XFILLER_182_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_551 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09126_ _09234_/S1 _09124_/X _09125_/X vssd1 vssd1 vccd1 vccd1 _09130_/B sky130_fd_sc_hd__a21o_1
XFILLER_124_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09057_ _13883_/Q _09231_/A2 _09522_/B1 _14398_/Q _09445_/C1 vssd1 vssd1 vccd1 vccd1
+ _09057_/X sky130_fd_sc_hd__a221o_1
XFILLER_136_768 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08008_ _08017_/D _08007_/Y _08012_/A2 vssd1 vssd1 vccd1 vccd1 _08008_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_1_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09959_ _11879_/A1 _14319_/Q _09963_/S vssd1 vssd1 vccd1 vccd1 _14319_/D sky130_fd_sc_hd__mux2_1
XFILLER_103_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12970_ _07408_/X _13024_/A2 _12969_/X _13024_/B2 vssd1 vssd1 vccd1 vccd1 _12970_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_181_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11921_ _12615_/A1 _11920_/X _12617_/S vssd1 vssd1 vccd1 vccd1 _11921_/X sky130_fd_sc_hd__a21o_1
XTAP_2700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14640_ _15644_/CLK _14640_/D vssd1 vssd1 vccd1 vccd1 _14640_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11852_ _15273_/Q _11852_/A1 _11878_/S vssd1 vssd1 vccd1 vccd1 _15273_/D sky130_fd_sc_hd__mux2_1
XTAP_2744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10803_ _14835_/Q _07319_/X _10868_/S vssd1 vssd1 vccd1 vccd1 _14835_/D sky130_fd_sc_hd__mux2_1
XTAP_2777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14571_ _15304_/CLK _14571_/D vssd1 vssd1 vccd1 vccd1 _14571_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11783_ _15207_/Q _12904_/S _11781_/Y _13809_/Q vssd1 vssd1 vccd1 vccd1 _15207_/D
+ sky130_fd_sc_hd__o22a_1
XTAP_2799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_52_clk clkbuf_5_8_0_clk/X vssd1 vssd1 vccd1 vccd1 _15042_/CLK sky130_fd_sc_hd__clkbuf_16
X_13522_ _15381_/CLK _13522_/D vssd1 vssd1 vccd1 vccd1 _13522_/Q sky130_fd_sc_hd__dfxtp_1
X_10734_ _15074_/Q _10734_/A2 _10731_/X _10733_/X vssd1 vssd1 vccd1 vccd1 _10734_/X
+ sky130_fd_sc_hd__o22a_4
XFILLER_9_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13453_ _15377_/CLK _13453_/D vssd1 vssd1 vccd1 vccd1 _13453_/Q sky130_fd_sc_hd__dfxtp_1
X_10665_ _14751_/Q _10664_/X _10665_/S vssd1 vssd1 vccd1 vccd1 _14751_/D sky130_fd_sc_hd__mux2_1
XFILLER_185_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12404_ _12592_/A1 _12403_/X _12548_/S vssd1 vssd1 vccd1 vccd1 _12404_/X sky130_fd_sc_hd__a21o_1
XFILLER_51_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13384_ _15650_/CLK _13384_/D vssd1 vssd1 vccd1 vccd1 _13384_/Q sky130_fd_sc_hd__dfxtp_1
X_10596_ _14998_/Q _10569_/B _10733_/A2 _14966_/Q _10732_/C1 vssd1 vssd1 vccd1 vccd1
+ _10596_/X sky130_fd_sc_hd__a221o_1
XFILLER_182_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15123_ _15507_/CLK _15123_/D vssd1 vssd1 vccd1 vccd1 _15123_/Q sky130_fd_sc_hd__dfxtp_1
X_12335_ _12615_/A1 _12334_/X _12536_/A vssd1 vssd1 vccd1 vccd1 _12335_/X sky130_fd_sc_hd__a21o_1
XFILLER_181_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15054_ _15054_/CLK _15054_/D vssd1 vssd1 vccd1 vccd1 _15054_/Q sky130_fd_sc_hd__dfxtp_4
X_12266_ _12500_/A1 _12265_/X _12582_/A vssd1 vssd1 vccd1 vccd1 _12266_/X sky130_fd_sc_hd__a21o_1
X_14005_ _15142_/CLK _14005_/D vssd1 vssd1 vccd1 vccd1 _14005_/Q sky130_fd_sc_hd__dfxtp_1
X_11217_ _10382_/D _15006_/Q _11232_/S vssd1 vssd1 vccd1 vccd1 _15006_/D sky130_fd_sc_hd__mux2_1
X_12197_ _12477_/A1 _12196_/X _12490_/A vssd1 vssd1 vccd1 vccd1 _12197_/X sky130_fd_sc_hd__a21o_1
XFILLER_68_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput70 _07125_/X vssd1 vssd1 vccd1 vccd1 ext_write_data[12] sky130_fd_sc_hd__clkbuf_2
Xoutput81 _07145_/X vssd1 vssd1 vccd1 vccd1 ext_write_data[22] sky130_fd_sc_hd__clkbuf_2
Xoutput92 _07111_/X vssd1 vssd1 vccd1 vccd1 ext_write_data[3] sky130_fd_sc_hd__clkbuf_2
X_11148_ _08233_/B _11147_/X _10984_/Y vssd1 vssd1 vccd1 vccd1 _11148_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_1_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11079_ _11259_/S _11079_/B vssd1 vssd1 vccd1 vccd1 _11079_/Y sky130_fd_sc_hd__nor2_1
XFILLER_48_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14907_ _15499_/CLK _14907_/D vssd1 vssd1 vccd1 vccd1 _14907_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_63_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14838_ _15497_/CLK _14838_/D vssd1 vssd1 vccd1 vccd1 _14838_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_1000 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14769_ _15620_/CLK _14769_/D vssd1 vssd1 vccd1 vccd1 _14769_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_43_clk clkbuf_5_9_0_clk/X vssd1 vssd1 vccd1 vccd1 _15584_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_16_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07310_ _07292_/A _07292_/B _07351_/B _07309_/X _07287_/X vssd1 vssd1 vccd1 vccd1
+ _07310_/X sky130_fd_sc_hd__o221a_1
XFILLER_108_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08290_ _08259_/Y _08289_/X _11047_/B vssd1 vssd1 vccd1 vccd1 _08290_/X sky130_fd_sc_hd__mux2_2
XFILLER_149_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_1066 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07241_ _07241_/A vssd1 vssd1 vccd1 vccd1 _07265_/B sky130_fd_sc_hd__inv_2
XFILLER_20_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07172_ _15346_/Q _15053_/Q _07188_/S vssd1 vssd1 vccd1 vccd1 _07172_/X sky130_fd_sc_hd__mux2_8
XFILLER_164_329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_395 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_5_22_0_clk clkbuf_5_23_0_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_5_22_0_clk/X
+ sky130_fd_sc_hd__clkbuf_8
Xfanout304 _07460_/X vssd1 vssd1 vccd1 vccd1 _13340_/A0 sky130_fd_sc_hd__buf_6
XFILLER_28_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout315 _07440_/X vssd1 vssd1 vccd1 vccd1 _11868_/A1 sky130_fd_sc_hd__buf_6
XFILLER_59_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout326 _07420_/X vssd1 vssd1 vccd1 vccd1 _13074_/B2 sky130_fd_sc_hd__buf_6
XFILLER_99_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09813_ _14179_/Q _13335_/A0 _09823_/S vssd1 vssd1 vccd1 vccd1 _14179_/D sky130_fd_sc_hd__mux2_1
Xfanout337 _13324_/A0 vssd1 vssd1 vccd1 vccd1 _11857_/A1 sky130_fd_sc_hd__buf_6
Xfanout348 _13319_/A0 vssd1 vssd1 vccd1 vccd1 _11852_/A1 sky130_fd_sc_hd__buf_6
XFILLER_101_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout359 _10568_/X vssd1 vssd1 vccd1 vccd1 _10732_/C1 sky130_fd_sc_hd__buf_12
XFILLER_101_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09744_ _14112_/Q _13332_/A0 _09757_/S vssd1 vssd1 vccd1 vccd1 _14112_/D sky130_fd_sc_hd__mux2_1
XFILLER_100_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06956_ _06728_/Y _13489_/Q _06730_/Y _13488_/Q _06955_/X vssd1 vssd1 vccd1 vccd1
+ _06956_/Y sky130_fd_sc_hd__o221ai_4
XFILLER_86_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09675_ _14046_/Q _13074_/B2 _09690_/S vssd1 vssd1 vccd1 vccd1 _14046_/D sky130_fd_sc_hd__mux2_1
X_06887_ _06702_/Y _13470_/Q _06704_/Y _13469_/Q vssd1 vssd1 vccd1 vccd1 _06929_/B
+ sky130_fd_sc_hd__a22o_1
XTAP_2007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08626_ _13788_/Q _08625_/X _08626_/S vssd1 vssd1 vccd1 vccd1 _13788_/D sky130_fd_sc_hd__mux2_1
XTAP_1306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08557_ _13608_/Q _08749_/A2 _08747_/A2 _13569_/Q vssd1 vssd1 vccd1 vccd1 _08557_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_168_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_34_clk clkbuf_5_13_0_clk/X vssd1 vssd1 vccd1 vccd1 _15537_/CLK sky130_fd_sc_hd__clkbuf_16
X_07508_ _14738_/Q _13417_/Q _07535_/S vssd1 vssd1 vccd1 vccd1 _13417_/D sky130_fd_sc_hd__mux2_1
X_08488_ _14591_/Q _08465_/B _08477_/X _14599_/Q _08487_/X vssd1 vssd1 vccd1 vccd1
+ _08488_/X sky130_fd_sc_hd__a221o_1
XFILLER_35_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_167_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07439_ _13665_/Q _07483_/A2 _07483_/B1 _14693_/Q _07438_/X vssd1 vssd1 vccd1 vccd1
+ _07439_/X sky130_fd_sc_hd__a221o_1
XFILLER_10_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10450_ _07219_/X _10360_/B _10449_/X vssd1 vssd1 vccd1 vccd1 _11582_/A sky130_fd_sc_hd__a21o_4
XFILLER_109_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09109_ _14077_/Q _09445_/A2 _09522_/B1 _14045_/Q _09221_/A vssd1 vssd1 vccd1 vccd1
+ _09109_/X sky130_fd_sc_hd__a221o_1
X_10381_ _10381_/A _10381_/B vssd1 vssd1 vccd1 vccd1 _10382_/D sky130_fd_sc_hd__nand2_1
XFILLER_124_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12120_ _14366_/Q _15182_/Q _13821_/Q _14560_/Q _12489_/S0 _12489_/S1 vssd1 vssd1
+ vccd1 vccd1 _12120_/X sky130_fd_sc_hd__mux4_1
XFILLER_163_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12051_ _14363_/Q _15179_/Q _13818_/Q _14557_/Q _12154_/S _12253_/S1 vssd1 vssd1
+ vccd1 vccd1 _12051_/X sky130_fd_sc_hd__mux4_1
XFILLER_77_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11002_ _10994_/X _11001_/X _11298_/A vssd1 vssd1 vccd1 vccd1 _11002_/X sky130_fd_sc_hd__mux2_1
XFILLER_120_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12953_ _15464_/Q _10877_/S _13116_/C _12952_/X vssd1 vssd1 vccd1 vccd1 _15464_/D
+ sky130_fd_sc_hd__a22o_1
XTAP_3231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11904_ _11887_/X _11888_/X _12260_/A vssd1 vssd1 vccd1 vccd1 _11904_/X sky130_fd_sc_hd__mux2_1
XTAP_3264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15672_ _15672_/CLK _15672_/D vssd1 vssd1 vccd1 vccd1 _15672_/Q sky130_fd_sc_hd__dfxtp_1
X_12884_ _15412_/Q _15597_/Q _12918_/S vssd1 vssd1 vccd1 vccd1 _15412_/D sky130_fd_sc_hd__mux2_1
XTAP_3275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14623_ _15626_/CLK _14623_/D vssd1 vssd1 vccd1 vccd1 _14623_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_2_3_1_clk clkbuf_2_3_1_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_7_0_clk/A sky130_fd_sc_hd__clkbuf_8
X_11835_ _15257_/Q _11868_/A1 _11849_/S vssd1 vssd1 vccd1 vccd1 _15257_/D sky130_fd_sc_hd__mux2_1
XFILLER_61_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_25_clk clkbuf_5_6_0_clk/X vssd1 vssd1 vccd1 vccd1 _15088_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_2585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_922 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_624 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14554_ _15176_/CLK _14554_/D vssd1 vssd1 vccd1 vccd1 _14554_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11766_ _11874_/A1 _15194_/Q _11775_/S vssd1 vssd1 vccd1 vccd1 _15194_/D sky130_fd_sc_hd__mux2_1
XTAP_1884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13505_ _14513_/CLK _13505_/D vssd1 vssd1 vccd1 vccd1 _13505_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_187_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10717_ _15022_/Q _10717_/A2 _10652_/B _15039_/Q _10717_/C1 vssd1 vssd1 vccd1 vccd1
+ _10717_/X sky130_fd_sc_hd__a221o_1
X_14485_ _14485_/CLK _14485_/D vssd1 vssd1 vccd1 vccd1 _14485_/Q sky130_fd_sc_hd__dfxtp_1
X_11697_ _11872_/A1 _15128_/Q _11708_/S vssd1 vssd1 vccd1 vccd1 _15128_/D sky130_fd_sc_hd__mux2_1
XFILLER_9_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13436_ _15393_/CLK _13436_/D vssd1 vssd1 vccd1 vccd1 _13436_/Q sky130_fd_sc_hd__dfxtp_1
X_10648_ _14976_/Q _10718_/A2 _10722_/B1 _14944_/Q _10647_/X vssd1 vssd1 vccd1 vccd1
+ _10648_/X sky130_fd_sc_hd__a221o_2
XFILLER_9_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13367_ _14470_/Q vssd1 vssd1 vccd1 vccd1 _14470_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_6_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10579_ _14734_/Q _10578_/X _10615_/S vssd1 vssd1 vccd1 vccd1 _14734_/D sky130_fd_sc_hd__mux2_1
XFILLER_127_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15106_ _15678_/CLK _15106_/D vssd1 vssd1 vccd1 vccd1 _15106_/Q sky130_fd_sc_hd__dfxtp_1
X_12318_ _12301_/X _12302_/X _12536_/A vssd1 vssd1 vccd1 vccd1 _12318_/X sky130_fd_sc_hd__mux2_1
XFILLER_138_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13298_ _12711_/X _15630_/Q _13309_/A vssd1 vssd1 vccd1 vccd1 _15630_/D sky130_fd_sc_hd__mux2_1
XFILLER_181_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15037_ _15041_/CLK _15037_/D vssd1 vssd1 vccd1 vccd1 _15037_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12249_ _12232_/X _12233_/X _12502_/S vssd1 vssd1 vccd1 vccd1 _12249_/X sky130_fd_sc_hd__mux2_1
XFILLER_96_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06810_ _13733_/Q _08668_/C _13049_/A1 _06666_/Y vssd1 vssd1 vccd1 vccd1 _06810_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_56_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07790_ _14735_/Q _07816_/A _07789_/Y _08084_/C1 vssd1 vssd1 vccd1 vccd1 _13510_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_110_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06741_ _13451_/Q vssd1 vssd1 vccd1 vccd1 _06741_/Y sky130_fd_sc_hd__inv_2
XFILLER_64_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_232 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09460_ _14545_/Q _14158_/Q _14190_/Q _14126_/Q _09469_/S _09546_/S1 vssd1 vssd1
+ vccd1 vccd1 _09460_/X sky130_fd_sc_hd__mux4_1
X_06672_ _08449_/A vssd1 vssd1 vccd1 vccd1 _06672_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_97_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08411_ _14597_/Q _08765_/A _14595_/Q _14588_/Q vssd1 vssd1 vccd1 vccd1 _08411_/X
+ sky130_fd_sc_hd__a31o_1
X_09391_ _09391_/A _09391_/B vssd1 vssd1 vccd1 vccd1 _09391_/X sky130_fd_sc_hd__or2_1
XFILLER_91_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_16_clk clkbuf_5_2_0_clk/X vssd1 vssd1 vccd1 vccd1 _15235_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_178_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08342_ _08244_/A _13763_/Q _15409_/Q _08244_/B vssd1 vssd1 vccd1 vccd1 _08342_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_178_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08273_ _08273_/A _11041_/A vssd1 vssd1 vccd1 vccd1 _08273_/X sky130_fd_sc_hd__or2_1
XFILLER_137_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07224_ _13937_/Q _15524_/Q _15527_/Q vssd1 vssd1 vccd1 vccd1 _07225_/A sky130_fd_sc_hd__mux2_8
XFILLER_146_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07155_ _07157_/A _07155_/B vssd1 vssd1 vccd1 vccd1 _07155_/X sky130_fd_sc_hd__and2_4
XFILLER_118_554 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07086_ _07085_/X _14761_/Q _07098_/S vssd1 vssd1 vccd1 vccd1 _13607_/D sky130_fd_sc_hd__mux2_1
XFILLER_65_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout112 _06852_/Y vssd1 vssd1 vccd1 vccd1 _13288_/S sky130_fd_sc_hd__buf_12
XFILLER_102_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout123 fanout138/X vssd1 vssd1 vccd1 vccd1 _10834_/S sky130_fd_sc_hd__buf_6
Xfanout134 _13149_/S vssd1 vssd1 vccd1 vccd1 _13154_/S sky130_fd_sc_hd__buf_12
Xfanout145 _12320_/A vssd1 vssd1 vccd1 vccd1 _12573_/A sky130_fd_sc_hd__buf_12
XFILLER_113_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout156 _06781_/X vssd1 vssd1 vccd1 vccd1 _12885_/S sky130_fd_sc_hd__buf_12
Xfanout167 _11851_/Y vssd1 vssd1 vccd1 vccd1 _11878_/S sky130_fd_sc_hd__buf_12
XFILLER_59_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout178 _11676_/X vssd1 vssd1 vccd1 vccd1 _11708_/S sky130_fd_sc_hd__buf_12
XFILLER_86_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07988_ _13563_/Q _07995_/D vssd1 vssd1 vccd1 vccd1 _07992_/B sky130_fd_sc_hd__nand2_1
Xfanout189 _09997_/X vssd1 vssd1 vccd1 vccd1 _10028_/S sky130_fd_sc_hd__buf_12
XFILLER_170_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09727_ _11816_/A1 _14097_/Q _09728_/S vssd1 vssd1 vccd1 vccd1 _14097_/D sky130_fd_sc_hd__mux2_1
XFILLER_74_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06939_ _13489_/Q _06728_/Y _06726_/Y _14499_/Q vssd1 vssd1 vccd1 vccd1 _06941_/C
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_28_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_243 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09658_ _14031_/Q _13347_/A0 _09661_/S vssd1 vssd1 vccd1 vccd1 _14031_/D sky130_fd_sc_hd__mux2_1
XTAP_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08609_ _15388_/Q _08748_/A2 _08736_/A2 _13433_/Q vssd1 vssd1 vccd1 vccd1 _08609_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_82_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09589_ _13965_/Q _13104_/B2 _09589_/S vssd1 vssd1 vccd1 vccd1 _13965_/D sky130_fd_sc_hd__mux2_1
XTAP_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_555 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11620_ wire360/X _11612_/B _11619_/X vssd1 vssd1 vccd1 vccd1 _11621_/B sky130_fd_sc_hd__o21a_1
XTAP_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11551_ _13218_/A _11537_/A _11537_/B _13236_/A vssd1 vssd1 vccd1 vccd1 _11552_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_168_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10502_ _11569_/B _13220_/B vssd1 vssd1 vccd1 vccd1 _10543_/B sky130_fd_sc_hd__nand2_1
XFILLER_184_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14270_ _15287_/CLK _14270_/D vssd1 vssd1 vccd1 vccd1 _14270_/Q sky130_fd_sc_hd__dfxtp_1
X_11482_ _11472_/A _11471_/A _11471_/B vssd1 vssd1 vccd1 vccd1 _11482_/X sky130_fd_sc_hd__o21ba_1
XFILLER_137_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13221_ _13236_/A _13220_/B _13214_/B _11569_/B vssd1 vssd1 vccd1 vccd1 _13221_/X
+ sky130_fd_sc_hd__a211o_1
X_10433_ _08244_/A _13746_/Q _15426_/Q _08244_/B vssd1 vssd1 vccd1 vccd1 _10433_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_137_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13152_ _14612_/Q _15550_/Q _13154_/S vssd1 vssd1 vccd1 vccd1 _15550_/D sky130_fd_sc_hd__mux2_1
X_10364_ _13202_/B _11496_/B vssd1 vssd1 vccd1 vccd1 _10365_/B sky130_fd_sc_hd__or2_1
XFILLER_128_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12103_ _12498_/A _12103_/B vssd1 vssd1 vccd1 vccd1 _12103_/X sky130_fd_sc_hd__and2_1
XTAP_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13083_ _15509_/Q _10834_/S _13105_/B1 _13082_/X vssd1 vssd1 vccd1 vccd1 _15509_/D
+ sky130_fd_sc_hd__a22o_1
X_10295_ _14680_/Q _14865_/Q _10615_/S vssd1 vssd1 vccd1 vccd1 _14680_/D sky130_fd_sc_hd__mux2_1
XFILLER_105_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12034_ _12590_/A _12034_/B vssd1 vssd1 vccd1 vccd1 _12034_/X sky130_fd_sc_hd__and2_1
XFILLER_77_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13985_ _15658_/CLK _13985_/D vssd1 vssd1 vccd1 vccd1 _13985_/Q sky130_fd_sc_hd__dfxtp_1
X_12936_ _06844_/X _12934_/Y _12935_/Y _06846_/X vssd1 vssd1 vccd1 vccd1 _12936_/X
+ sky130_fd_sc_hd__o211a_2
XFILLER_92_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12867_ _14761_/Q _15395_/Q _12871_/S vssd1 vssd1 vccd1 vccd1 _15395_/D sky130_fd_sc_hd__mux2_1
X_15655_ _15655_/CLK _15655_/D vssd1 vssd1 vccd1 vccd1 _15655_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_2_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11818_ _11818_/A _11851_/B vssd1 vssd1 vccd1 vccd1 _11818_/Y sky130_fd_sc_hd__nor2_8
X_14606_ _14606_/CLK _14606_/D vssd1 vssd1 vccd1 vccd1 _14606_/Q sky130_fd_sc_hd__dfxtp_4
X_15586_ _15620_/CLK _15586_/D vssd1 vssd1 vccd1 vccd1 _15586_/Q sky130_fd_sc_hd__dfxtp_1
X_12798_ _12810_/C _12798_/B vssd1 vssd1 vccd1 vccd1 _12799_/B sky130_fd_sc_hd__and2b_1
XTAP_1670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_942 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14537_ _14537_/CLK _14537_/D vssd1 vssd1 vccd1 vccd1 _14537_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11749_ _11857_/A1 _15177_/Q _11775_/S vssd1 vssd1 vccd1 vccd1 _15177_/D sky130_fd_sc_hd__mux2_1
XFILLER_186_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14468_ _14468_/CLK _14468_/D vssd1 vssd1 vccd1 vccd1 _14468_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_159 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13419_ _15374_/CLK _13419_/D vssd1 vssd1 vccd1 vccd1 _13419_/Q sky130_fd_sc_hd__dfxtp_2
X_14399_ _14530_/CLK _14399_/D vssd1 vssd1 vccd1 vccd1 _14399_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_155_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08960_ _13942_/Q _13684_/Q _09073_/S vssd1 vssd1 vccd1 vccd1 _08960_/X sky130_fd_sc_hd__mux2_1
XFILLER_142_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_5_clk clkbuf_5_1_0_clk/X vssd1 vssd1 vccd1 vccd1 _15660_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_102_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07911_ _08022_/B _07911_/B vssd1 vssd1 vccd1 vccd1 _07911_/Y sky130_fd_sc_hd__nand2_1
X_08891_ _14228_/Q _14260_/Q _14292_/Q _14324_/Q _09132_/S _08988_/A1 vssd1 vssd1
+ vccd1 vccd1 _08891_/X sky130_fd_sc_hd__mux4_1
XFILLER_97_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07842_ _07844_/B _07841_/X _07830_/A vssd1 vssd1 vccd1 vccd1 _07842_/X sky130_fd_sc_hd__a21bo_1
XFILLER_69_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07773_ _07777_/A _07773_/B vssd1 vssd1 vccd1 vccd1 _07773_/Y sky130_fd_sc_hd__nand2_1
XFILLER_17_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09512_ _15678_/Q _13412_/Q _09512_/S vssd1 vssd1 vccd1 vccd1 _09512_/X sky130_fd_sc_hd__mux2_1
X_06724_ _13491_/Q vssd1 vssd1 vccd1 vccd1 _06724_/Y sky130_fd_sc_hd__inv_2
XFILLER_71_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09443_ _09446_/A1 _09441_/X _09442_/X vssd1 vssd1 vccd1 vccd1 _09443_/X sky130_fd_sc_hd__a21o_1
XFILLER_52_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09374_ _14477_/Q _14445_/Q _13866_/Q _14219_/Q _09535_/S _08508_/B vssd1 vssd1 vccd1
+ vccd1 _09374_/X sky130_fd_sc_hd__mux4_1
XFILLER_33_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08325_ _07302_/X _10523_/A2 _08324_/X vssd1 vssd1 vccd1 vccd1 _11431_/A sky130_fd_sc_hd__a21oi_4
XFILLER_21_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08256_ _11356_/C _10895_/B vssd1 vssd1 vccd1 vccd1 _10551_/B sky130_fd_sc_hd__or2_2
XFILLER_165_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07207_ _15331_/Q _15487_/Q _07340_/S vssd1 vssd1 vccd1 vccd1 _07208_/A sky130_fd_sc_hd__mux2_4
XFILLER_4_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08187_ _14715_/Q _08817_/B vssd1 vssd1 vccd1 vccd1 _11743_/C sky130_fd_sc_hd__nand2_4
XFILLER_118_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_822 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07138_ _14849_/Q _14841_/Q _07146_/S vssd1 vssd1 vccd1 vccd1 _07138_/X sky130_fd_sc_hd__mux2_1
XFILLER_134_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07069_ _14635_/Q _14667_/Q _07078_/S vssd1 vssd1 vccd1 vccd1 _07069_/X sky130_fd_sc_hd__mux2_1
XFILLER_121_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10080_ _14436_/Q _13080_/B2 _10092_/S vssd1 vssd1 vccd1 vccd1 _14436_/D sky130_fd_sc_hd__mux2_1
XFILLER_58_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13770_ _15587_/CLK _13770_/D vssd1 vssd1 vccd1 vccd1 _13770_/Q sky130_fd_sc_hd__dfxtp_1
X_10982_ _10965_/X _10981_/X _11129_/A vssd1 vssd1 vccd1 vccd1 _10982_/X sky130_fd_sc_hd__mux2_2
XFILLER_74_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_179 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12721_ _12737_/A _12721_/B vssd1 vssd1 vccd1 vccd1 _12721_/X sky130_fd_sc_hd__or2_1
XFILLER_55_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_516 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15440_ _15626_/CLK _15440_/D vssd1 vssd1 vccd1 vccd1 _15440_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12652_ _15049_/Q _12651_/X _12834_/B vssd1 vssd1 vccd1 vccd1 _12652_/X sky130_fd_sc_hd__mux2_1
XFILLER_71_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11603_ _11611_/A _11603_/B vssd1 vssd1 vccd1 vccd1 _11606_/B sky130_fd_sc_hd__nor2_1
X_15371_ _15372_/CLK _15371_/D vssd1 vssd1 vccd1 vccd1 _15371_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12583_ _06670_/A _12580_/X _06671_/A vssd1 vssd1 vccd1 vccd1 _12583_/X sky130_fd_sc_hd__o21a_1
XFILLER_129_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14322_ _15303_/CLK _14322_/D vssd1 vssd1 vccd1 vccd1 _14322_/Q sky130_fd_sc_hd__dfxtp_1
X_11534_ _11534_/A _11544_/B vssd1 vssd1 vccd1 vccd1 _11534_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_129_638 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14253_ _15662_/CLK _14253_/D vssd1 vssd1 vccd1 vccd1 _14253_/Q sky130_fd_sc_hd__dfxtp_1
X_11465_ _11474_/S _11472_/B _11465_/C vssd1 vssd1 vccd1 vccd1 _11465_/X sky130_fd_sc_hd__or3_1
XFILLER_125_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13204_ _10362_/X _13202_/X _13203_/Y _13214_/B _15568_/Q vssd1 vssd1 vccd1 vccd1
+ _15568_/D sky130_fd_sc_hd__a32o_1
XFILLER_104_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10416_ _13189_/B _11476_/A _10379_/Y _10415_/X vssd1 vssd1 vccd1 vccd1 _10416_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_171_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14184_ _15161_/CLK _14184_/D vssd1 vssd1 vccd1 vccd1 _14184_/Q sky130_fd_sc_hd__dfxtp_1
X_11396_ _11414_/A _11437_/A _11414_/D _13242_/A vssd1 vssd1 vccd1 vccd1 _11397_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_174_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13135_ _15532_/Q _10892_/B _13129_/Y _13134_/X vssd1 vssd1 vccd1 vccd1 _15532_/D
+ sky130_fd_sc_hd__a211o_1
X_10347_ _07197_/A _10457_/A2 _10346_/X vssd1 vssd1 vccd1 vccd1 _13252_/A sky130_fd_sc_hd__a21oi_4
XFILLER_124_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13066_ _12966_/X _13104_/A2 _13104_/B1 _13326_/A0 vssd1 vssd1 vccd1 vccd1 _13066_/X
+ sky130_fd_sc_hd__a22o_1
X_10278_ _14663_/Q _14816_/Q _10665_/S vssd1 vssd1 vccd1 vccd1 _14663_/D sky130_fd_sc_hd__mux2_1
XFILLER_140_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12017_ _12592_/A1 _12016_/X _06670_/A vssd1 vssd1 vccd1 vccd1 _12017_/X sky130_fd_sc_hd__a21o_1
XFILLER_38_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_1070 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13968_ _15651_/CLK _13968_/D vssd1 vssd1 vccd1 vccd1 _13968_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12919_ hold2/A _15633_/Q _12928_/S vssd1 vssd1 vccd1 vccd1 _15447_/D sky130_fd_sc_hd__mux2_1
XFILLER_179_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13899_ _15673_/CLK _13899_/D vssd1 vssd1 vccd1 vccd1 _13899_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15638_ _15638_/CLK _15638_/D vssd1 vssd1 vccd1 vccd1 _15638_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15569_ _15569_/CLK _15569_/D vssd1 vssd1 vccd1 vccd1 _15569_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_148_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08110_ input14/X input22/X _08133_/S vssd1 vssd1 vccd1 vccd1 _08165_/B sky130_fd_sc_hd__mux2_1
X_09090_ _13884_/Q _09231_/A2 _09403_/B1 _14399_/Q _09437_/A1 vssd1 vssd1 vccd1 vccd1
+ _09090_/X sky130_fd_sc_hd__a221o_1
X_08041_ _14734_/Q _13612_/Q _08072_/S vssd1 vssd1 vccd1 vccd1 _13612_/D sky130_fd_sc_hd__mux2_1
XFILLER_162_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09992_ _11879_/A1 _14351_/Q _09996_/S vssd1 vssd1 vccd1 vccd1 _14351_/D sky130_fd_sc_hd__mux2_1
XFILLER_103_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_227 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08943_ _09524_/A _08943_/B _08943_/C vssd1 vssd1 vccd1 vccd1 _08943_/X sky130_fd_sc_hd__and3_1
XFILLER_130_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_4_15_0_clk clkbuf_3_7_0_clk/X vssd1 vssd1 vccd1 vccd1 clkbuf_5_31_0_clk/A
+ sky130_fd_sc_hd__clkbuf_8
X_08874_ _13895_/Q _11872_/A1 _08885_/S vssd1 vssd1 vccd1 vccd1 _13895_/D sky130_fd_sc_hd__mux2_1
XFILLER_57_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07825_ _13520_/Q _13519_/Q _13518_/Q _07825_/D vssd1 vssd1 vccd1 vccd1 _07836_/D
+ sky130_fd_sc_hd__and4_4
XTAP_3819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07756_ _13503_/Q _07756_/B vssd1 vssd1 vccd1 vccd1 _07756_/Y sky130_fd_sc_hd__nor2_1
XFILLER_25_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06707_ _13500_/Q vssd1 vssd1 vccd1 vccd1 _06707_/Y sky130_fd_sc_hd__inv_2
XFILLER_37_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07687_ _13484_/Q _13483_/Q _07687_/C vssd1 vssd1 vccd1 vccd1 _07717_/A sky130_fd_sc_hd__and3_4
XFILLER_13_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09426_ _13900_/Q _09445_/A2 _09522_/B1 _14415_/Q _09437_/A1 vssd1 vssd1 vccd1 vccd1
+ _09426_/X sky130_fd_sc_hd__a221o_1
XFILLER_80_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09357_ _14025_/Q _13993_/Q _09521_/S vssd1 vssd1 vccd1 vccd1 _09357_/X sky130_fd_sc_hd__mux2_1
X_08308_ _11047_/B _08274_/X _08307_/X vssd1 vssd1 vccd1 vccd1 _08309_/B sky130_fd_sc_hd__o21ai_1
XFILLER_166_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09288_ _13862_/Q _14215_/Q _09484_/S vssd1 vssd1 vccd1 vccd1 _09288_/X sky130_fd_sc_hd__mux2_1
X_08239_ _08240_/A _13805_/Q _07327_/A _10457_/A2 _08237_/X vssd1 vssd1 vccd1 vccd1
+ _11053_/S sky130_fd_sc_hd__a221o_4
XFILLER_107_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11250_ _08385_/Y _11249_/Y _11318_/S vssd1 vssd1 vccd1 vccd1 _11252_/B sky130_fd_sc_hd__mux2_1
XFILLER_153_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10201_ input26/X _14586_/Q _13284_/S vssd1 vssd1 vccd1 vccd1 _14586_/D sky130_fd_sc_hd__mux2_1
XFILLER_106_343 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11181_ _11199_/A _11181_/B vssd1 vssd1 vccd1 vccd1 _11181_/Y sky130_fd_sc_hd__nor2_1
XFILLER_106_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10132_ _11851_/A _10132_/B vssd1 vssd1 vccd1 vccd1 _10132_/Y sky130_fd_sc_hd__nor2_8
XFILLER_122_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14940_ _15006_/CLK _14940_/D vssd1 vssd1 vccd1 vccd1 _14940_/Q sky130_fd_sc_hd__dfxtp_1
X_10063_ _14420_/Q _11816_/A1 _10064_/S vssd1 vssd1 vccd1 vccd1 _14420_/D sky130_fd_sc_hd__mux2_1
XFILLER_76_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14871_ _15422_/CLK _14871_/D vssd1 vssd1 vccd1 vccd1 _14871_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13822_ _15220_/CLK _13822_/D vssd1 vssd1 vccd1 vccd1 _13822_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_141_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13753_ _14649_/CLK _13753_/D vssd1 vssd1 vccd1 vccd1 _13753_/Q sky130_fd_sc_hd__dfxtp_1
X_10965_ _10959_/Y _10964_/X _11252_/A vssd1 vssd1 vccd1 vccd1 _10965_/X sky130_fd_sc_hd__mux2_1
XFILLER_43_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12704_ _15056_/Q _12703_/X _12792_/B vssd1 vssd1 vccd1 vccd1 _12704_/X sky130_fd_sc_hd__mux2_1
XFILLER_188_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13684_ _15202_/CLK _13684_/D vssd1 vssd1 vccd1 vccd1 _13684_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10896_ _14930_/Q _10895_/X _10951_/B vssd1 vssd1 vccd1 vccd1 _14930_/D sky130_fd_sc_hd__mux2_1
X_15423_ _15608_/CLK _15423_/D vssd1 vssd1 vccd1 vccd1 _15423_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12635_ _15340_/Q _15339_/Q _15338_/Q vssd1 vssd1 vccd1 vccd1 _12644_/B sky130_fd_sc_hd__and3_1
XFILLER_34_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15354_ _15354_/CLK _15354_/D vssd1 vssd1 vccd1 vccd1 _15354_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_157_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12566_ _14032_/Q _14000_/Q _12568_/S vssd1 vssd1 vccd1 vccd1 _12567_/B sky130_fd_sc_hd__mux2_1
XFILLER_180_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11517_ _11516_/X _15060_/Q _11614_/S vssd1 vssd1 vccd1 vccd1 _15060_/D sky130_fd_sc_hd__mux2_1
X_14305_ _15287_/CLK _14305_/D vssd1 vssd1 vccd1 vccd1 _14305_/Q sky130_fd_sc_hd__dfxtp_1
X_15285_ _15285_/CLK _15285_/D vssd1 vssd1 vccd1 vccd1 _15285_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_172_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12497_ _14029_/Q _13997_/Q _12499_/S vssd1 vssd1 vccd1 vccd1 _12498_/B sky130_fd_sc_hd__mux2_1
XFILLER_138_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_438 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14236_ _14462_/CLK _14236_/D vssd1 vssd1 vccd1 vccd1 _14236_/Q sky130_fd_sc_hd__dfxtp_1
X_11448_ _11449_/A _11449_/B vssd1 vssd1 vccd1 vccd1 _11450_/A sky130_fd_sc_hd__nand2_1
XFILLER_153_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14167_ _15273_/CLK _14167_/D vssd1 vssd1 vccd1 vccd1 _14167_/Q sky130_fd_sc_hd__dfxtp_1
X_11379_ _11378_/Y _15046_/Q _11641_/S vssd1 vssd1 vccd1 vccd1 _15046_/D sky130_fd_sc_hd__mux2_1
XFILLER_4_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13118_ _13042_/Y _13118_/A2 _13051_/B _12904_/S _07334_/S vssd1 vssd1 vccd1 vccd1
+ _15527_/D sky130_fd_sc_hd__o32a_1
XTAP_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_492 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14098_ _14439_/CLK _14098_/D vssd1 vssd1 vccd1 vccd1 _14098_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13049_ _13049_/A1 _13318_/C _08817_/Y _09466_/A _13048_/X vssd1 vssd1 vccd1 vccd1
+ _13050_/C sky130_fd_sc_hd__o221a_1
XFILLER_22_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07610_ _13464_/Q _13463_/Q _07610_/C vssd1 vssd1 vccd1 vccd1 _07617_/C sky130_fd_sc_hd__and3_2
XFILLER_66_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08590_ _13564_/Q _08747_/A2 _08691_/B1 _13500_/Q vssd1 vssd1 vccd1 vccd1 _08590_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_38_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_3_4_0_clk clkbuf_3_5_0_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_9_0_clk/A sky130_fd_sc_hd__clkbuf_8
XFILLER_19_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07541_ _13446_/Q _13445_/Q vssd1 vssd1 vccd1 vccd1 _07542_/B sky130_fd_sc_hd__xnor2_1
XFILLER_46_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07472_ _14758_/Q _07471_/X _07480_/S vssd1 vssd1 vccd1 vccd1 _07472_/X sky130_fd_sc_hd__mux2_8
XFILLER_35_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09211_ _09406_/S1 _09209_/X _09210_/X vssd1 vssd1 vccd1 vccd1 _09212_/C sky130_fd_sc_hd__a21o_1
XFILLER_14_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09142_ _14240_/Q _14272_/Q _14304_/Q _14336_/Q _09407_/S _09406_/S1 vssd1 vssd1
+ vccd1 vccd1 _09142_/X sky130_fd_sc_hd__mux4_1
XFILLER_175_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09073_ _13851_/Q _14204_/Q _09073_/S vssd1 vssd1 vccd1 vccd1 _09073_/X sky130_fd_sc_hd__mux2_1
XFILLER_129_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_747 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08024_ _13574_/Q _12640_/S _06863_/B _13573_/Q vssd1 vssd1 vccd1 vccd1 _08028_/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_135_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09975_ _13329_/A0 _14334_/Q _09991_/S vssd1 vssd1 vccd1 vccd1 _14334_/D sky130_fd_sc_hd__mux2_1
XFILLER_103_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_208 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08926_ _13134_/A _08926_/B _08926_/C vssd1 vssd1 vccd1 vccd1 _08926_/X sky130_fd_sc_hd__and3_2
XFILLER_162_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08857_ _13878_/Q _11680_/A0 _08880_/S vssd1 vssd1 vccd1 vccd1 _13878_/D sky130_fd_sc_hd__mux2_1
XFILLER_111_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_220_clk clkbuf_5_18_0_clk/X vssd1 vssd1 vccd1 vccd1 _15523_/CLK sky130_fd_sc_hd__clkbuf_16
X_07808_ _07810_/B _07807_/X _07816_/A vssd1 vssd1 vccd1 vccd1 _07808_/X sky130_fd_sc_hd__a21bo_1
XTAP_2904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08788_ _13322_/A0 _13814_/Q _08811_/S vssd1 vssd1 vccd1 vccd1 _13814_/D sky130_fd_sc_hd__mux2_1
XFILLER_72_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07739_ _13498_/Q _13497_/Q _07739_/C vssd1 vssd1 vccd1 vccd1 _07746_/C sky130_fd_sc_hd__and3_2
XTAP_2948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10750_ _15414_/Q _14782_/Q _10764_/S vssd1 vssd1 vccd1 vccd1 _14782_/D sky130_fd_sc_hd__mux2_1
XFILLER_25_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09409_ _15100_/Q _13130_/B1 _09408_/X _09450_/B1 vssd1 vssd1 vccd1 vccd1 _09409_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_158_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10681_ _15015_/Q _10567_/Y _10718_/A2 _14983_/Q _10717_/C1 vssd1 vssd1 vccd1 vccd1
+ _10681_/X sky130_fd_sc_hd__a221o_1
XFILLER_71_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12420_ _15296_/Q _15264_/Q _15232_/Q _15163_/Q _12430_/S _12563_/A vssd1 vssd1 vccd1
+ vccd1 _12421_/B sky130_fd_sc_hd__mux4_1
XFILLER_187_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12351_ _15293_/Q _15261_/Q _15229_/Q _15160_/Q _12541_/S _12540_/A vssd1 vssd1 vccd1
+ vccd1 _12352_/B sky130_fd_sc_hd__mux4_1
X_11302_ _11302_/A _11344_/A vssd1 vssd1 vccd1 vccd1 _11303_/A sky130_fd_sc_hd__nand2_4
X_15070_ _15579_/CLK _15070_/D vssd1 vssd1 vccd1 vccd1 _15070_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_14_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12282_ _15290_/Q _15258_/Q _15226_/Q _15157_/Q _12568_/S _12567_/A vssd1 vssd1 vccd1
+ vccd1 _12283_/B sky130_fd_sc_hd__mux4_1
X_14021_ _15677_/CLK _14021_/D vssd1 vssd1 vccd1 vccd1 _14021_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_135_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11233_ _10470_/C _15021_/Q _11237_/S vssd1 vssd1 vccd1 vccd1 _15021_/D sky130_fd_sc_hd__mux2_1
XFILLER_106_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_278 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11164_ _14976_/Q _11163_/X _11164_/S vssd1 vssd1 vccd1 vccd1 _14976_/D sky130_fd_sc_hd__mux2_1
XFILLER_96_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10115_ _14501_/Q _14749_/Q _10124_/S vssd1 vssd1 vccd1 vccd1 _14501_/D sky130_fd_sc_hd__mux2_1
XFILLER_67_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11095_ _11115_/S _10964_/X _11094_/Y vssd1 vssd1 vccd1 vccd1 _11096_/B sky130_fd_sc_hd__a21o_1
X_10046_ _14403_/Q _13078_/B2 _10059_/S vssd1 vssd1 vccd1 vccd1 _14403_/D sky130_fd_sc_hd__mux2_1
X_14923_ _15208_/CLK _14923_/D vssd1 vssd1 vccd1 vccd1 _14923_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_49_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_211_clk clkbuf_5_16_0_clk/X vssd1 vssd1 vccd1 vccd1 _15130_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_48_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14854_ _15518_/CLK _14854_/D vssd1 vssd1 vccd1 vccd1 _14854_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13805_ _14863_/CLK _13805_/D vssd1 vssd1 vccd1 vccd1 _13805_/Q sky130_fd_sc_hd__dfxtp_2
X_14785_ _15453_/CLK _14785_/D vssd1 vssd1 vccd1 vccd1 _14785_/Q sky130_fd_sc_hd__dfxtp_1
X_11997_ _12273_/A1 _11996_/X _11995_/X _12503_/C1 vssd1 vssd1 vccd1 vccd1 _11998_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_21_1095 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10948_ _11626_/A _10948_/B vssd1 vssd1 vccd1 vccd1 _10948_/Y sky130_fd_sc_hd__nand2_1
XFILLER_17_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13736_ _15540_/CLK _13736_/D vssd1 vssd1 vccd1 vccd1 _13736_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13667_ _14774_/CLK _13667_/D vssd1 vssd1 vccd1 vccd1 _13667_/Q sky130_fd_sc_hd__dfxtp_1
X_10879_ _14911_/Q _15542_/Q _13134_/A vssd1 vssd1 vccd1 vccd1 _14911_/D sky130_fd_sc_hd__mux2_1
X_15406_ _15591_/CLK _15406_/D vssd1 vssd1 vccd1 vccd1 _15406_/Q sky130_fd_sc_hd__dfxtp_2
X_12618_ _12618_/A1 _12617_/X _12616_/X _12618_/C1 vssd1 vssd1 vccd1 vccd1 _12619_/C
+ sky130_fd_sc_hd__a211o_1
X_13598_ _15354_/CLK _13598_/D vssd1 vssd1 vccd1 vccd1 _13598_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_169_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_714 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12549_ _12618_/A1 _12548_/X _12547_/X _12618_/C1 vssd1 vssd1 vccd1 vccd1 _12550_/C
+ sky130_fd_sc_hd__a211o_1
X_15337_ _15676_/CLK _15337_/D vssd1 vssd1 vccd1 vccd1 _15337_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_144_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_1 _07202_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15268_ _15544_/CLK _15268_/D vssd1 vssd1 vccd1 vccd1 _15268_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_172_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14219_ _15336_/CLK _14219_/D vssd1 vssd1 vccd1 vccd1 _14219_/Q sky130_fd_sc_hd__dfxtp_1
X_15199_ _15199_/CLK _15199_/D vssd1 vssd1 vccd1 vccd1 _15199_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_141_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout508 _14711_/Q vssd1 vssd1 vccd1 vccd1 _07498_/B sky130_fd_sc_hd__buf_8
Xfanout519 _09435_/A vssd1 vssd1 vccd1 vccd1 _09221_/A sky130_fd_sc_hd__buf_12
XFILLER_140_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09760_ _14128_/Q _13348_/A0 _09762_/S vssd1 vssd1 vccd1 vccd1 _14128_/D sky130_fd_sc_hd__mux2_1
X_06972_ _06710_/Y _13498_/Q _14506_/Q _06713_/Y vssd1 vssd1 vccd1 vccd1 _06972_/X
+ sky130_fd_sc_hd__o2bb2a_1
XTAP_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08711_ _13514_/Q _08750_/A2 _08750_/B1 _13617_/Q vssd1 vssd1 vccd1 vccd1 _08711_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09691_ _14062_/Q _13346_/A0 _09695_/S vssd1 vssd1 vccd1 vccd1 _14062_/D sky130_fd_sc_hd__mux2_1
XFILLER_55_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_202_clk clkbuf_5_16_0_clk/X vssd1 vssd1 vccd1 vccd1 _15081_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_82_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08642_ _13428_/Q _08690_/B1 _08693_/A2 _14501_/Q vssd1 vssd1 vccd1 vccd1 _08642_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_27_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08573_ _13780_/Q _08572_/X _08573_/S vssd1 vssd1 vccd1 vccd1 _13780_/D sky130_fd_sc_hd__mux2_1
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07524_ _14754_/Q _13433_/Q _07535_/S vssd1 vssd1 vccd1 vccd1 _13433_/D sky130_fd_sc_hd__mux2_1
XFILLER_41_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07455_ _13669_/Q _07483_/A2 _07483_/B1 _14697_/Q _07454_/X vssd1 vssd1 vccd1 vccd1
+ _07455_/X sky130_fd_sc_hd__a221o_1
XFILLER_50_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07386_ _14648_/Q _07498_/B _07498_/C vssd1 vssd1 vccd1 vccd1 _07386_/X sky130_fd_sc_hd__and3_1
XFILLER_22_399 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09125_ _13886_/Q _09231_/A2 _09403_/B1 _14401_/Q _09445_/C1 vssd1 vssd1 vccd1 vccd1
+ _09125_/X sky130_fd_sc_hd__a221o_1
XFILLER_157_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09056_ _13947_/Q _13689_/Q _09230_/S vssd1 vssd1 vccd1 vccd1 _09056_/X sky130_fd_sc_hd__mux2_1
XFILLER_151_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08007_ _13567_/Q _13566_/Q _08006_/D _13568_/Q vssd1 vssd1 vccd1 vccd1 _08007_/Y
+ sky130_fd_sc_hd__a31oi_1
XFILLER_135_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xmax_cap281 _07907_/A vssd1 vssd1 vccd1 vccd1 _07660_/B sky130_fd_sc_hd__buf_2
XFILLER_103_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09958_ _13104_/B2 _14318_/Q _09958_/S vssd1 vssd1 vccd1 vccd1 _14318_/D sky130_fd_sc_hd__mux2_1
XFILLER_106_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08909_ _14229_/Q _14261_/Q _14293_/Q _14325_/Q _09469_/S _09546_/S1 vssd1 vssd1
+ vccd1 vccd1 _08909_/X sky130_fd_sc_hd__mux4_1
XFILLER_100_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09889_ _13098_/B2 _14251_/Q _09897_/S vssd1 vssd1 vccd1 vccd1 _14251_/D sky130_fd_sc_hd__mux2_1
XFILLER_85_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11920_ _13876_/Q _14391_/Q _12522_/S vssd1 vssd1 vccd1 vccd1 _11920_/X sky130_fd_sc_hd__mux2_1
XFILLER_131_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11851_ _11851_/A _11851_/B vssd1 vssd1 vccd1 vccd1 _11851_/Y sky130_fd_sc_hd__nor2_8
XTAP_3479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_108 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10802_ _14834_/Q _07322_/X _10868_/S vssd1 vssd1 vccd1 vccd1 _14834_/D sky130_fd_sc_hd__mux2_1
XTAP_2767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14570_ _15293_/CLK _14570_/D vssd1 vssd1 vccd1 vccd1 _14570_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11782_ _15206_/Q _10892_/B _11781_/A _13810_/Q vssd1 vssd1 vccd1 vccd1 _15206_/D
+ sky130_fd_sc_hd__a22o_1
XTAP_2789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13521_ _15381_/CLK _13521_/D vssd1 vssd1 vccd1 vccd1 _13521_/Q sky130_fd_sc_hd__dfxtp_1
X_10733_ _14993_/Q _10733_/A2 _10733_/B1 _14961_/Q _10732_/X vssd1 vssd1 vccd1 vccd1
+ _10733_/X sky130_fd_sc_hd__a221o_1
XFILLER_159_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13452_ _15375_/CLK _13452_/D vssd1 vssd1 vccd1 vccd1 _13452_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_9_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10664_ _15060_/Q _10714_/A2 _10661_/X _10663_/X vssd1 vssd1 vccd1 vccd1 _10664_/X
+ sky130_fd_sc_hd__o22a_4
XFILLER_9_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12403_ _13897_/Q _14412_/Q _12407_/S vssd1 vssd1 vccd1 vccd1 _12403_/X sky130_fd_sc_hd__mux2_1
XFILLER_90_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13383_ _15649_/CLK _13383_/D vssd1 vssd1 vccd1 vccd1 _13383_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_167_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10595_ _14737_/Q _10594_/X _10615_/S vssd1 vssd1 vccd1 vccd1 _14737_/D sky130_fd_sc_hd__mux2_1
XFILLER_51_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12334_ _13894_/Q _14409_/Q _12543_/S vssd1 vssd1 vccd1 vccd1 _12334_/X sky130_fd_sc_hd__mux2_1
X_15122_ _15658_/CLK _15122_/D vssd1 vssd1 vccd1 vccd1 _15122_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_182_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15053_ _15054_/CLK _15053_/D vssd1 vssd1 vccd1 vccd1 _15053_/Q sky130_fd_sc_hd__dfxtp_4
X_12265_ _13891_/Q _14406_/Q _12269_/S vssd1 vssd1 vccd1 vccd1 _12265_/X sky130_fd_sc_hd__mux2_1
XFILLER_114_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14004_ _15125_/CLK _14004_/D vssd1 vssd1 vccd1 vccd1 _14004_/Q sky130_fd_sc_hd__dfxtp_1
X_11216_ _10382_/C _15005_/Q _11232_/S vssd1 vssd1 vccd1 vccd1 _15005_/D sky130_fd_sc_hd__mux2_1
XFILLER_141_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12196_ _13888_/Q _14403_/Q _12499_/S vssd1 vssd1 vccd1 vccd1 _12196_/X sky130_fd_sc_hd__mux2_1
XFILLER_123_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput60 _07166_/X vssd1 vssd1 vccd1 vccd1 ext_address[4] sky130_fd_sc_hd__clkbuf_2
XFILLER_122_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput71 _07127_/X vssd1 vssd1 vccd1 vccd1 ext_write_data[13] sky130_fd_sc_hd__clkbuf_2
Xoutput82 _07147_/X vssd1 vssd1 vccd1 vccd1 ext_write_data[23] sky130_fd_sc_hd__clkbuf_2
XFILLER_1_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput93 _07112_/X vssd1 vssd1 vccd1 vccd1 ext_write_data[4] sky130_fd_sc_hd__clkbuf_2
XFILLER_123_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11147_ _11077_/X _11086_/X _11298_/A vssd1 vssd1 vccd1 vccd1 _11147_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11078_ _13251_/A _11362_/C _11362_/B vssd1 vssd1 vccd1 vccd1 _11363_/B sky130_fd_sc_hd__o21ai_4
XFILLER_64_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10029_ _11883_/A1 _14387_/Q _10029_/S vssd1 vssd1 vccd1 vccd1 _14387_/D sky130_fd_sc_hd__mux2_1
X_14906_ _15540_/CLK _14906_/D vssd1 vssd1 vccd1 vccd1 _14906_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_63_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14837_ _15501_/CLK _14837_/D vssd1 vssd1 vccd1 vccd1 _14837_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_3980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14768_ _15619_/CLK _14768_/D vssd1 vssd1 vccd1 vccd1 _14768_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_108_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13719_ _15042_/CLK _13719_/D vssd1 vssd1 vccd1 vccd1 _13719_/Q sky130_fd_sc_hd__dfxtp_1
X_14699_ _15624_/CLK _14699_/D vssd1 vssd1 vccd1 vccd1 _14699_/Q sky130_fd_sc_hd__dfxtp_1
X_07240_ _15326_/Q _15482_/Q _07335_/S vssd1 vssd1 vccd1 vccd1 _07241_/A sky130_fd_sc_hd__mux2_8
XFILLER_108_1078 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07171_ _15345_/Q _15052_/Q _07188_/S vssd1 vssd1 vccd1 vccd1 _07171_/X sky130_fd_sc_hd__mux2_8
XFILLER_9_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_780 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout305 _13339_/A0 vssd1 vssd1 vccd1 vccd1 _11872_/A1 sky130_fd_sc_hd__buf_6
Xfanout316 _07440_/X vssd1 vssd1 vccd1 vccd1 _13335_/A0 sky130_fd_sc_hd__buf_4
XFILLER_98_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09812_ _14178_/Q _13334_/A0 _09823_/S vssd1 vssd1 vccd1 vccd1 _14178_/D sky130_fd_sc_hd__mux2_1
XFILLER_101_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout327 _13072_/B2 vssd1 vssd1 vccd1 vccd1 _13329_/A0 sky130_fd_sc_hd__buf_6
Xfanout338 _13324_/A0 vssd1 vssd1 vccd1 vccd1 _11649_/A0 sky130_fd_sc_hd__clkbuf_4
XFILLER_99_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout349 _07376_/X vssd1 vssd1 vccd1 vccd1 _13319_/A0 sky130_fd_sc_hd__buf_6
XFILLER_115_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06955_ _06944_/A _06941_/B _06934_/X vssd1 vssd1 vccd1 vccd1 _06955_/X sky130_fd_sc_hd__a21bo_1
X_09743_ _14111_/Q _13331_/A0 _09757_/S vssd1 vssd1 vccd1 vccd1 _14111_/D sky130_fd_sc_hd__mux2_1
XFILLER_67_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09674_ _14045_/Q _13072_/B2 _09690_/S vssd1 vssd1 vccd1 vccd1 _14045_/D sky130_fd_sc_hd__mux2_1
X_06886_ _15394_/Q _06701_/Y _06702_/Y _13470_/Q vssd1 vssd1 vccd1 vccd1 _06888_/A
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_36_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08625_ _15386_/Q _08748_/A2 _08622_/X _08623_/X _08624_/X vssd1 vssd1 vccd1 vccd1
+ _08625_/X sky130_fd_sc_hd__a2111o_2
XTAP_2019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_108 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08556_ _15396_/Q _08748_/A2 _08736_/A2 _13441_/Q vssd1 vssd1 vccd1 vccd1 _08556_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_42_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07507_ _14737_/Q _13416_/Q _07535_/S vssd1 vssd1 vccd1 vccd1 _13416_/D sky130_fd_sc_hd__mux2_1
XFILLER_52_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08487_ _08487_/A _08487_/B vssd1 vssd1 vccd1 vccd1 _08487_/X sky130_fd_sc_hd__and2_1
XFILLER_146_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07438_ _14661_/Q _07474_/B _07482_/C vssd1 vssd1 vccd1 vccd1 _07438_/X sky130_fd_sc_hd__and3_1
XFILLER_183_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_628 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07369_ _14712_/Q _14713_/Q _08817_/B vssd1 vssd1 vccd1 vccd1 _11710_/A sky130_fd_sc_hd__nand3_4
X_09108_ _14013_/Q _13981_/Q _09425_/S vssd1 vssd1 vccd1 vccd1 _09108_/X sky130_fd_sc_hd__mux2_1
XFILLER_136_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10380_ _11457_/A _11475_/B vssd1 vssd1 vccd1 vccd1 _10381_/B sky130_fd_sc_hd__or2_1
XFILLER_109_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09039_ _15280_/Q _15248_/Q _15216_/Q _15147_/Q _09225_/S0 _09225_/S1 vssd1 vssd1
+ vccd1 vccd1 _09039_/X sky130_fd_sc_hd__mux4_1
XFILLER_105_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12050_ _12046_/X _12047_/X _12260_/A vssd1 vssd1 vccd1 vccd1 _12050_/X sky130_fd_sc_hd__mux2_1
XFILLER_123_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11001_ _11362_/B _11000_/X _10997_/X _10996_/Y vssd1 vssd1 vccd1 vccd1 _11001_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_131_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_712 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12952_ _07384_/X _13039_/A2 _12951_/X _12944_/A vssd1 vssd1 vccd1 vccd1 _12952_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_73_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11903_ _11896_/X _11898_/X _11900_/X _11902_/X _12501_/C1 vssd1 vssd1 vccd1 vccd1
+ _11903_/X sky130_fd_sc_hd__o221a_1
XTAP_3265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15671_ _15679_/CLK _15671_/D vssd1 vssd1 vccd1 vccd1 _15671_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12883_ _15411_/Q _15596_/Q _12917_/S vssd1 vssd1 vccd1 vccd1 _15411_/D sky130_fd_sc_hd__mux2_1
XTAP_3276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14622_ _15628_/CLK _14622_/D vssd1 vssd1 vccd1 vccd1 _14622_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11834_ _15256_/Q _13334_/A0 _11849_/S vssd1 vssd1 vccd1 vccd1 _15256_/D sky130_fd_sc_hd__mux2_1
XTAP_2564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14553_ _15212_/CLK _14553_/D vssd1 vssd1 vccd1 vccd1 _14553_/Q sky130_fd_sc_hd__dfxtp_1
X_11765_ _11873_/A1 _15193_/Q _11775_/S vssd1 vssd1 vccd1 vccd1 _15193_/D sky130_fd_sc_hd__mux2_1
XFILLER_187_934 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10716_ _15581_/Q _10731_/B vssd1 vssd1 vccd1 vccd1 _10716_/X sky130_fd_sc_hd__and2_1
X_13504_ _14513_/CLK _13504_/D vssd1 vssd1 vccd1 vccd1 _13504_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_186_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11696_ _13338_/A0 _15127_/Q _11708_/S vssd1 vssd1 vccd1 vccd1 _15127_/D sky130_fd_sc_hd__mux2_1
X_14484_ _15672_/CLK _14484_/D vssd1 vssd1 vccd1 vccd1 _14484_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_187_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10647_ _15008_/Q _10717_/A2 _10652_/B _13727_/Q _10717_/C1 vssd1 vssd1 vccd1 vccd1
+ _10647_/X sky130_fd_sc_hd__a221o_1
X_13435_ _15393_/CLK _13435_/D vssd1 vssd1 vccd1 vccd1 _13435_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_139_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13366_ _14469_/Q vssd1 vssd1 vccd1 vccd1 _14469_/D sky130_fd_sc_hd__clkbuf_2
X_10578_ _07146_/S _10734_/A2 _10572_/X _10577_/X vssd1 vssd1 vccd1 vccd1 _10578_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_154_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15105_ _15226_/CLK _15105_/D vssd1 vssd1 vccd1 vccd1 _15105_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_155_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12317_ _12310_/X _12312_/X _12314_/X _12316_/X _12616_/C1 vssd1 vssd1 vccd1 vccd1
+ _12317_/X sky130_fd_sc_hd__o221a_1
X_13297_ _12703_/X _15629_/Q _13300_/S vssd1 vssd1 vccd1 vccd1 _15629_/D sky130_fd_sc_hd__mux2_1
XFILLER_177_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15036_ _15041_/CLK _15036_/D vssd1 vssd1 vccd1 vccd1 _15036_/Q sky130_fd_sc_hd__dfxtp_1
X_12248_ _12241_/X _12243_/X _12245_/X _12247_/X _12455_/C1 vssd1 vssd1 vccd1 vccd1
+ _12248_/X sky130_fd_sc_hd__o221a_1
XFILLER_96_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12179_ _12172_/X _12174_/X _12176_/X _12178_/X _12455_/C1 vssd1 vssd1 vccd1 vccd1
+ _12179_/X sky130_fd_sc_hd__o221a_1
XFILLER_111_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_306 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06740_ _14492_/Q vssd1 vssd1 vccd1 vccd1 _06740_/Y sky130_fd_sc_hd__inv_2
XFILLER_114_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06671_ _06671_/A vssd1 vssd1 vccd1 vccd1 _06671_/Y sky130_fd_sc_hd__inv_4
XFILLER_36_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_1006 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08410_ _14597_/Q _14595_/Q vssd1 vssd1 vccd1 vccd1 _08410_/Y sky130_fd_sc_hd__nand2_1
XFILLER_97_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09390_ _14380_/Q _15196_/Q _13835_/Q _14574_/Q _09407_/S _09406_/S1 vssd1 vssd1
+ vccd1 vccd1 _09391_/B sky130_fd_sc_hd__mux4_1
XFILLER_145_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_439 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08341_ _11037_/A _11440_/A vssd1 vssd1 vccd1 vccd1 _11033_/B sky130_fd_sc_hd__and2_1
XFILLER_149_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08272_ _11349_/B _13165_/B vssd1 vssd1 vccd1 vccd1 _11041_/A sky130_fd_sc_hd__nor2_1
XFILLER_165_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07223_ _15336_/Q _15492_/Q _07340_/S vssd1 vssd1 vccd1 vccd1 _07227_/A sky130_fd_sc_hd__mux2_8
XFILLER_121_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07154_ _14857_/Q _14849_/Q _14841_/Q _14833_/Q _07146_/S _07104_/C vssd1 vssd1 vccd1
+ vccd1 _07155_/B sky130_fd_sc_hd__mux4_2
XFILLER_118_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07085_ _07084_/X _13607_/Q _12662_/S vssd1 vssd1 vccd1 vccd1 _07085_/X sky130_fd_sc_hd__mux2_1
XFILLER_106_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout113 _13041_/Y vssd1 vssd1 vccd1 vccd1 _13105_/B1 sky130_fd_sc_hd__buf_12
XFILLER_87_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout124 fanout138/X vssd1 vssd1 vccd1 vccd1 _13119_/S sky130_fd_sc_hd__clkbuf_16
XFILLER_99_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout135 fanout138/X vssd1 vssd1 vccd1 vccd1 _13149_/S sky130_fd_sc_hd__buf_8
Xfanout146 _12904_/S vssd1 vssd1 vccd1 vccd1 _13134_/A sky130_fd_sc_hd__clkbuf_16
Xfanout157 _08573_/S vssd1 vssd1 vccd1 vccd1 _12932_/S sky130_fd_sc_hd__buf_12
Xfanout168 _11851_/Y vssd1 vssd1 vccd1 vccd1 _11883_/S sky130_fd_sc_hd__buf_12
XFILLER_102_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07987_ _14755_/Q _07971_/A _07986_/Y _07987_/C1 vssd1 vssd1 vccd1 vccd1 _13562_/D
+ sky130_fd_sc_hd__o211a_1
Xfanout179 _11643_/X vssd1 vssd1 vccd1 vccd1 _11670_/S sky130_fd_sc_hd__buf_12
XFILLER_87_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06938_ _14496_/Q _06732_/Y _06734_/Y _13486_/Q vssd1 vssd1 vccd1 vccd1 _06941_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_09726_ _11881_/A1 _14096_/Q _09728_/S vssd1 vssd1 vccd1 vccd1 _14096_/D sky130_fd_sc_hd__mux2_1
XFILLER_41_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09657_ _14030_/Q _13346_/A0 _09661_/S vssd1 vssd1 vccd1 vccd1 _14030_/D sky130_fd_sc_hd__mux2_1
X_06869_ _14511_/Q _06703_/Y _14510_/Q _06705_/Y vssd1 vssd1 vccd1 vccd1 _06879_/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_28_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08608_ _13600_/Q _08691_/A2 _08685_/A2 _13561_/Q _08607_/X vssd1 vssd1 vccd1 vccd1
+ _08612_/B sky130_fd_sc_hd__a221o_1
XTAP_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09588_ _13964_/Q _13344_/A0 _09589_/S vssd1 vssd1 vccd1 vccd1 _13964_/D sky130_fd_sc_hd__mux2_1
XTAP_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08539_ _13775_/Q _08573_/S _08527_/X _08534_/X vssd1 vssd1 vccd1 vccd1 _13775_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_42_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11550_ _11549_/Y _15063_/Q _11614_/S vssd1 vssd1 vccd1 vccd1 _15063_/D sky130_fd_sc_hd__mux2_1
XFILLER_11_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10501_ _13220_/B vssd1 vssd1 vccd1 vccd1 _11555_/A sky130_fd_sc_hd__inv_2
XFILLER_10_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11481_ _11502_/A _11481_/B vssd1 vssd1 vccd1 vccd1 _11505_/C sky130_fd_sc_hd__nor2_2
XFILLER_10_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13220_ _13236_/A _13220_/B vssd1 vssd1 vccd1 vccd1 _13220_/Y sky130_fd_sc_hd__nor2_1
X_10432_ _07202_/X _08225_/Y _10431_/X vssd1 vssd1 vccd1 vccd1 _11616_/A sky130_fd_sc_hd__a21oi_4
XFILLER_6_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13151_ _14611_/Q _15549_/Q _13154_/S vssd1 vssd1 vccd1 vccd1 _15549_/D sky130_fd_sc_hd__mux2_1
X_10363_ _13202_/B _11496_/B vssd1 vssd1 vccd1 vccd1 _10418_/B sky130_fd_sc_hd__nand2_1
XFILLER_136_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12102_ _13948_/Q _13690_/Q _12246_/S vssd1 vssd1 vccd1 vccd1 _12103_/B sky130_fd_sc_hd__mux2_1
XFILLER_152_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13082_ _12990_/X _13104_/A2 _13104_/B1 _13082_/B2 vssd1 vssd1 vccd1 vccd1 _13082_/X
+ sky130_fd_sc_hd__a22o_1
X_10294_ _14679_/Q _14864_/Q _10735_/S vssd1 vssd1 vccd1 vccd1 _14679_/D sky130_fd_sc_hd__mux2_1
X_12033_ _13945_/Q _13687_/Q _12591_/S vssd1 vssd1 vccd1 vccd1 _12034_/B sky130_fd_sc_hd__mux2_1
XFILLER_2_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13984_ _15659_/CLK _13984_/D vssd1 vssd1 vccd1 vccd1 _13984_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_74_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12935_ _12379_/A _08406_/B _12934_/Y vssd1 vssd1 vccd1 vccd1 _12935_/Y sky130_fd_sc_hd__o21ai_1
XTAP_3051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15654_ _15654_/CLK _15654_/D vssd1 vssd1 vccd1 vccd1 _15654_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12866_ _14760_/Q _15394_/Q _12866_/S vssd1 vssd1 vccd1 vccd1 _15394_/D sky130_fd_sc_hd__mux2_1
XFILLER_33_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14605_ _15613_/CLK _14605_/D vssd1 vssd1 vccd1 vccd1 _14605_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_21_409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11817_ _15240_/Q _13350_/A0 _11817_/S vssd1 vssd1 vccd1 vccd1 _15240_/D sky130_fd_sc_hd__mux2_1
XTAP_2394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15585_ _15617_/CLK _15585_/D vssd1 vssd1 vccd1 vccd1 _15585_/Q sky130_fd_sc_hd__dfxtp_1
X_12797_ _15362_/Q _13309_/B vssd1 vssd1 vccd1 vccd1 _12798_/B sky130_fd_sc_hd__or2_1
XTAP_1671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_5_21_0_clk clkbuf_5_21_0_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_5_21_0_clk/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_18_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14536_ _15667_/CLK _14536_/D vssd1 vssd1 vccd1 vccd1 _14536_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11748_ _13323_/A0 _15176_/Q _11774_/S vssd1 vssd1 vccd1 vccd1 _15176_/D sky130_fd_sc_hd__mux2_1
XFILLER_14_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14467_ _15235_/CLK _14467_/D vssd1 vssd1 vccd1 vccd1 _14467_/Q sky130_fd_sc_hd__dfxtp_1
X_11679_ _13321_/A0 _15110_/Q _11708_/S vssd1 vssd1 vccd1 vccd1 _15110_/D sky130_fd_sc_hd__mux2_1
X_13418_ _14493_/CLK _13418_/D vssd1 vssd1 vccd1 vccd1 _13418_/Q sky130_fd_sc_hd__dfxtp_1
X_14398_ _15657_/CLK _14398_/D vssd1 vssd1 vccd1 vccd1 _14398_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13349_ _13349_/A0 _15679_/Q _13350_/S vssd1 vssd1 vccd1 vccd1 _15679_/D sky130_fd_sc_hd__mux2_1
XFILLER_52_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15019_ _15020_/CLK _15019_/D vssd1 vssd1 vccd1 vccd1 _15019_/Q sky130_fd_sc_hd__dfxtp_1
X_07910_ _13542_/Q _07910_/B vssd1 vssd1 vccd1 vccd1 _07911_/B sky130_fd_sc_hd__xor2_1
X_08890_ _14454_/Q _14422_/Q _13843_/Q _14196_/Q _09225_/S0 _09225_/S1 vssd1 vssd1
+ vccd1 vccd1 _08890_/X sky130_fd_sc_hd__mux4_1
XFILLER_25_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07841_ _13524_/Q _07847_/D vssd1 vssd1 vccd1 vccd1 _07841_/X sky130_fd_sc_hd__or2_1
XFILLER_56_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07772_ _13507_/Q _07776_/C vssd1 vssd1 vccd1 vccd1 _07773_/B sky130_fd_sc_hd__xnor2_1
XFILLER_37_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06723_ _13460_/Q vssd1 vssd1 vccd1 vccd1 _07595_/A sky130_fd_sc_hd__inv_2
X_09511_ _14547_/Q _14160_/Q _14192_/Q _14128_/Q _09512_/S _09511_/S1 vssd1 vssd1
+ vccd1 vccd1 _09511_/X sky130_fd_sc_hd__mux4_1
XFILLER_83_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09442_ _14093_/Q _09445_/A2 _09522_/B1 _14061_/Q _09435_/A vssd1 vssd1 vccd1 vccd1
+ _09442_/X sky130_fd_sc_hd__a221o_1
XFILLER_92_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09373_ _14251_/Q _14283_/Q _14315_/Q _14347_/Q _09535_/S _08494_/B vssd1 vssd1 vccd1
+ vccd1 _09373_/X sky130_fd_sc_hd__mux4_1
XFILLER_24_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08324_ _08244_/A _13765_/Q _15407_/Q _08244_/B vssd1 vssd1 vccd1 vccd1 _08324_/X
+ sky130_fd_sc_hd__a22o_2
XFILLER_177_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08255_ _11356_/C _10895_/B vssd1 vssd1 vccd1 vccd1 _11360_/A sky130_fd_sc_hd__nor2_1
XFILLER_137_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07206_ _13932_/Q _15519_/Q _07339_/S vssd1 vssd1 vccd1 vccd1 _07206_/X sky130_fd_sc_hd__mux2_8
XFILLER_137_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08186_ _13680_/Q _10610_/S _08155_/X _08185_/X vssd1 vssd1 vccd1 vccd1 _13680_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_119_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07137_ _14832_/Q _07104_/X _07136_/X _07131_/A vssd1 vssd1 vccd1 vccd1 _07137_/X
+ sky130_fd_sc_hd__a22o_2
XFILLER_119_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07068_ _07067_/X _14755_/Q _07077_/S vssd1 vssd1 vccd1 vccd1 _13601_/D sky130_fd_sc_hd__mux2_1
XFILLER_106_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_2_2_1_clk clkbuf_2_2_1_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_5_0_clk/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09709_ _11689_/A0 _14079_/Q _09723_/S vssd1 vssd1 vccd1 vccd1 _14079_/D sky130_fd_sc_hd__mux2_1
X_10981_ _10973_/Y _10980_/Y _11252_/A vssd1 vssd1 vccd1 vccd1 _10981_/X sky130_fd_sc_hd__mux2_1
XFILLER_62_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12720_ _13428_/Q _12719_/X _12728_/S vssd1 vssd1 vccd1 vccd1 _12721_/B sky130_fd_sc_hd__mux2_1
XFILLER_15_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12651_ _15342_/Q _12657_/C vssd1 vssd1 vccd1 vccd1 _12651_/X sky130_fd_sc_hd__xor2_1
XFILLER_31_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11602_ _13236_/B _11602_/B vssd1 vssd1 vccd1 vccd1 _11603_/B sky130_fd_sc_hd__nor2_1
X_12582_ _12582_/A _12582_/B vssd1 vssd1 vccd1 vccd1 _12582_/X sky130_fd_sc_hd__or2_1
X_15370_ _15543_/CLK _15370_/D vssd1 vssd1 vccd1 vccd1 _15370_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_184_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14321_ _15526_/CLK _14321_/D vssd1 vssd1 vccd1 vccd1 _14321_/Q sky130_fd_sc_hd__dfxtp_1
X_11533_ _11530_/X _11533_/B vssd1 vssd1 vccd1 vccd1 _11544_/B sky130_fd_sc_hd__nand2b_1
XFILLER_23_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_424 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11464_ _11505_/A _11464_/B _11464_/C vssd1 vssd1 vccd1 vccd1 _11465_/C sky130_fd_sc_hd__nor3_1
XFILLER_7_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14252_ _14542_/CLK _14252_/D vssd1 vssd1 vccd1 vccd1 _14252_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10415_ _13189_/B _11476_/A _10387_/X _10414_/X _10389_/B vssd1 vssd1 vccd1 vccd1
+ _10415_/X sky130_fd_sc_hd__o221a_1
X_13203_ _13233_/A _13202_/B _13214_/B vssd1 vssd1 vccd1 vccd1 _13203_/Y sky130_fd_sc_hd__a21oi_1
X_14183_ _15096_/CLK _14183_/D vssd1 vssd1 vccd1 vccd1 _14183_/Q sky130_fd_sc_hd__dfxtp_1
X_11395_ _11394_/Y _15048_/Q _11641_/S vssd1 vssd1 vccd1 vccd1 _15048_/D sky130_fd_sc_hd__mux2_1
XFILLER_87_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13134_ _13134_/A _13134_/B _13134_/C vssd1 vssd1 vccd1 vccd1 _13134_/X sky130_fd_sc_hd__and3_1
X_10346_ _08240_/A _13775_/Q _13743_/Q _08237_/A vssd1 vssd1 vccd1 vccd1 _10346_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_151_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13065_ _15500_/Q _13139_/S _13105_/B1 _13064_/X vssd1 vssd1 vccd1 vccd1 _15500_/D
+ sky130_fd_sc_hd__a22o_1
X_10277_ _14662_/Q _14815_/Q _10665_/S vssd1 vssd1 vccd1 vccd1 _14662_/D sky130_fd_sc_hd__mux2_1
X_12016_ _14072_/Q _14040_/Q _12407_/S vssd1 vssd1 vccd1 vccd1 _12016_/X sky130_fd_sc_hd__mux2_1
XFILLER_2_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13967_ _15259_/CLK _13967_/D vssd1 vssd1 vccd1 vccd1 _13967_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12918_ _15446_/Q _15632_/Q _12918_/S vssd1 vssd1 vccd1 vccd1 _15446_/D sky130_fd_sc_hd__mux2_1
XFILLER_73_180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13898_ _15527_/CLK _13898_/D vssd1 vssd1 vccd1 vccd1 _13898_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15637_ _15637_/CLK _15637_/D vssd1 vssd1 vccd1 vccd1 _15637_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12849_ _14743_/Q _15377_/Q _12866_/S vssd1 vssd1 vccd1 vccd1 _15377_/D sky130_fd_sc_hd__mux2_1
XFILLER_34_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15568_ _15572_/CLK _15568_/D vssd1 vssd1 vccd1 vccd1 _15568_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14519_ _15650_/CLK _14519_/D vssd1 vssd1 vccd1 vccd1 _14519_/Q sky130_fd_sc_hd__dfxtp_1
X_15499_ _15499_/CLK _15499_/D vssd1 vssd1 vccd1 vccd1 _15499_/Q sky130_fd_sc_hd__dfxtp_1
X_08040_ _12839_/B _14717_/Q _08074_/A vssd1 vssd1 vccd1 vccd1 _08040_/X sky130_fd_sc_hd__or3b_4
XFILLER_31_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_973 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09991_ _13104_/B2 _14350_/Q _09991_/S vssd1 vssd1 vccd1 vccd1 _14350_/D sky130_fd_sc_hd__mux2_1
XFILLER_103_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08942_ _09523_/A1 _08940_/X _08941_/X vssd1 vssd1 vccd1 vccd1 _08943_/C sky130_fd_sc_hd__a21o_1
XFILLER_88_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08873_ _13894_/Q _13338_/A0 _08885_/S vssd1 vssd1 vccd1 vccd1 _13894_/D sky130_fd_sc_hd__mux2_1
XFILLER_96_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_572 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_103 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07824_ _14744_/Q _07830_/A _07823_/Y _12788_/C1 vssd1 vssd1 vccd1 vccd1 _13519_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_3809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07755_ _14759_/Q _07750_/A _07754_/Y _08012_/C1 vssd1 vssd1 vccd1 vccd1 _13502_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_44_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06706_ _15391_/Q vssd1 vssd1 vccd1 vccd1 _06918_/A sky130_fd_sc_hd__inv_2
X_07686_ _13484_/Q _07686_/B vssd1 vssd1 vccd1 vccd1 _07686_/Y sky130_fd_sc_hd__nor2_1
XFILLER_44_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09425_ _13964_/Q _13706_/Q _09425_/S vssd1 vssd1 vccd1 vccd1 _09425_/X sky130_fd_sc_hd__mux2_1
XFILLER_13_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09356_ _08668_/D _09352_/X _09355_/X _09351_/X vssd1 vssd1 vccd1 vccd1 _09356_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_178_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08307_ _11362_/B _08307_/B vssd1 vssd1 vccd1 vccd1 _08307_/X sky130_fd_sc_hd__or2_1
XFILLER_138_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09287_ _14247_/Q _14279_/Q _14311_/Q _14343_/Q _09484_/S _08519_/A vssd1 vssd1 vccd1
+ vccd1 _09287_/X sky130_fd_sc_hd__mux4_1
XFILLER_20_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08238_ _08240_/A _13805_/Q _07327_/A _10457_/A2 _08237_/X vssd1 vssd1 vccd1 vccd1
+ _08238_/Y sky130_fd_sc_hd__a221oi_4
XFILLER_181_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08169_ _08185_/A _08169_/B vssd1 vssd1 vccd1 vccd1 _08169_/X sky130_fd_sc_hd__and2_1
XFILLER_109_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10200_ input23/X _14585_/Q _13284_/S vssd1 vssd1 vccd1 vccd1 _14585_/D sky130_fd_sc_hd__mux2_1
X_11180_ _14982_/Q _11202_/A _11170_/X _11179_/Y vssd1 vssd1 vccd1 vccd1 _14982_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_106_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_206 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10131_ _14517_/Q _14765_/Q _10131_/S vssd1 vssd1 vccd1 vccd1 _14517_/D sky130_fd_sc_hd__mux2_1
XFILLER_134_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10062_ _14419_/Q _11881_/A1 _10064_/S vssd1 vssd1 vccd1 vccd1 _14419_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14870_ _15607_/CLK _14870_/D vssd1 vssd1 vccd1 vccd1 _14870_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13821_ _15298_/CLK _13821_/D vssd1 vssd1 vccd1 vccd1 _13821_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_72 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13752_ _14703_/CLK _13752_/D vssd1 vssd1 vccd1 vccd1 _13752_/Q sky130_fd_sc_hd__dfxtp_1
X_10964_ _10960_/X _10963_/Y _11259_/S vssd1 vssd1 vccd1 vccd1 _10964_/X sky130_fd_sc_hd__mux2_1
XFILLER_141_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12703_ _12710_/B _12703_/B vssd1 vssd1 vccd1 vccd1 _12703_/X sky130_fd_sc_hd__and2b_1
XFILLER_43_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13683_ _15275_/CLK _13683_/D vssd1 vssd1 vccd1 vccd1 _13683_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10895_ _11349_/B _10895_/B vssd1 vssd1 vccd1 vccd1 _10895_/X sky130_fd_sc_hd__or2_1
X_15422_ _15422_/CLK _15422_/D vssd1 vssd1 vccd1 vccd1 _15422_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12634_ _15339_/Q _12759_/B _12633_/X _12832_/C1 vssd1 vssd1 vccd1 vccd1 _15339_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_34_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_180_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15353_ _15634_/CLK _15353_/D vssd1 vssd1 vccd1 vccd1 _15353_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_141_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_520 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12565_ _12592_/A1 _12564_/X _12594_/S vssd1 vssd1 vccd1 vccd1 _12565_/X sky130_fd_sc_hd__a21o_1
X_14304_ _15184_/CLK _14304_/D vssd1 vssd1 vccd1 vccd1 _14304_/Q sky130_fd_sc_hd__dfxtp_1
X_11516_ _11516_/A _11546_/B vssd1 vssd1 vccd1 vccd1 _11516_/X sky130_fd_sc_hd__xor2_1
XFILLER_8_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_1018 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15284_ _15284_/CLK _15284_/D vssd1 vssd1 vccd1 vccd1 _15284_/Q sky130_fd_sc_hd__dfxtp_1
X_12496_ _12500_/A1 _12495_/X _12490_/A vssd1 vssd1 vccd1 vccd1 _12496_/X sky130_fd_sc_hd__a21o_1
XFILLER_184_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14235_ _15660_/CLK _14235_/D vssd1 vssd1 vccd1 vccd1 _14235_/Q sky130_fd_sc_hd__dfxtp_1
X_11447_ _11476_/A _11447_/B vssd1 vssd1 vccd1 vccd1 _11449_/B sky130_fd_sc_hd__xnor2_1
XFILLER_171_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14166_ _15276_/CLK _14166_/D vssd1 vssd1 vccd1 vccd1 _14166_/Q sky130_fd_sc_hd__dfxtp_1
X_11378_ _11378_/A _11378_/B vssd1 vssd1 vccd1 vccd1 _11378_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_124_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13117_ _07335_/S _12904_/S _13116_/X vssd1 vssd1 vccd1 vccd1 _15526_/D sky130_fd_sc_hd__o21ba_1
X_10329_ _14907_/Q _14714_/Q _10566_/B vssd1 vssd1 vccd1 vccd1 _14714_/D sky130_fd_sc_hd__mux2_1
XTAP_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14097_ _14420_/CLK _14097_/D vssd1 vssd1 vccd1 vccd1 _14097_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13048_ _08508_/B _08852_/B _11743_/C _09382_/A vssd1 vssd1 vccd1 vccd1 _13048_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_38_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14999_ _15558_/CLK _14999_/D vssd1 vssd1 vccd1 vccd1 _14999_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07540_ _14734_/Q _07644_/A _07539_/Y _08084_/C1 vssd1 vssd1 vccd1 vccd1 _13445_/D
+ sky130_fd_sc_hd__o211a_1
X_07471_ _13673_/Q _07483_/A2 _07483_/B1 _14701_/Q _07470_/X vssd1 vssd1 vccd1 vccd1
+ _07471_/X sky130_fd_sc_hd__a221o_1
XFILLER_90_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09210_ _14082_/Q _09445_/A2 _09522_/B1 _14050_/Q _09221_/A vssd1 vssd1 vccd1 vccd1
+ _09210_/X sky130_fd_sc_hd__a221o_1
XFILLER_148_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09141_ _09445_/C1 _09140_/X _09139_/X _09130_/A vssd1 vssd1 vccd1 vccd1 _09141_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_175_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09072_ _14236_/Q _14268_/Q _14300_/Q _14332_/Q _09073_/S _09530_/S1 vssd1 vssd1
+ vccd1 vccd1 _09072_/X sky130_fd_sc_hd__mux4_1
XFILLER_163_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08023_ _08022_/B _08021_/Y _08022_/Y input35/X vssd1 vssd1 vccd1 vccd1 _13572_/D
+ sky130_fd_sc_hd__a211oi_1
XFILLER_147_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_759 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09974_ _11861_/A1 _14333_/Q _09991_/S vssd1 vssd1 vccd1 vccd1 _14333_/D sky130_fd_sc_hd__mux2_1
XFILLER_118_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08925_ _08507_/Y _08921_/X _08924_/X _08920_/X vssd1 vssd1 vccd1 vccd1 _08926_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_58_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08856_ _13877_/Q _11854_/A1 _08885_/S vssd1 vssd1 vccd1 vccd1 _13877_/D sky130_fd_sc_hd__mux2_1
XTAP_3606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07807_ _13515_/Q _07813_/D vssd1 vssd1 vccd1 vccd1 _07807_/X sky130_fd_sc_hd__or2_1
XTAP_3639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08787_ _11854_/A1 _13813_/Q _08816_/S vssd1 vssd1 vccd1 vccd1 _13813_/D sky130_fd_sc_hd__mux2_1
XFILLER_84_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_832 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07738_ _13497_/Q _07739_/C _13498_/Q vssd1 vssd1 vccd1 vccd1 _07738_/Y sky130_fd_sc_hd__a21oi_1
XTAP_2938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07669_ _07777_/A _07669_/B vssd1 vssd1 vccd1 vccd1 _07669_/Y sky130_fd_sc_hd__nand2_1
XFILLER_111_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09408_ _15132_/Q _09536_/A2 _08520_/B _09407_/X vssd1 vssd1 vccd1 vccd1 _09408_/X
+ sky130_fd_sc_hd__a22o_1
X_10680_ _14754_/Q _10679_/X _10715_/S vssd1 vssd1 vccd1 vccd1 _14754_/D sky130_fd_sc_hd__mux2_1
XFILLER_185_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09339_ _09546_/S1 _09337_/X _09338_/X vssd1 vssd1 vccd1 vccd1 _09340_/C sky130_fd_sc_hd__a21o_1
XFILLER_40_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12350_ _14376_/Q _15192_/Q _13831_/Q _14570_/Q _12541_/S _12540_/A vssd1 vssd1 vccd1
+ vccd1 _12350_/X sky130_fd_sc_hd__mux4_1
XFILLER_166_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11301_ _15034_/Q _08232_/A _11300_/X vssd1 vssd1 vccd1 vccd1 _15034_/D sky130_fd_sc_hd__a21o_1
XFILLER_153_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12281_ _14373_/Q _15189_/Q _13828_/Q _14567_/Q _12430_/S _12563_/A vssd1 vssd1 vccd1
+ vccd1 _12281_/X sky130_fd_sc_hd__mux4_1
XFILLER_181_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11232_ _10470_/A _15020_/Q _11232_/S vssd1 vssd1 vccd1 vccd1 _15020_/D sky130_fd_sc_hd__mux2_1
X_14020_ _15668_/CLK _14020_/D vssd1 vssd1 vccd1 vccd1 _14020_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11163_ _11199_/A _11199_/B _11161_/Y _11162_/X vssd1 vssd1 vccd1 vccd1 _11163_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_96_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_931 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10114_ _14500_/Q _14748_/Q _10124_/S vssd1 vssd1 vccd1 vccd1 _14500_/D sky130_fd_sc_hd__mux2_1
X_11094_ _11115_/S _11129_/B vssd1 vssd1 vccd1 vccd1 _11094_/Y sky130_fd_sc_hd__nor2_2
XFILLER_96_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10045_ _14402_/Q _11689_/A0 _10059_/S vssd1 vssd1 vccd1 vccd1 _14402_/D sky130_fd_sc_hd__mux2_1
X_14922_ _15618_/CLK _14922_/D vssd1 vssd1 vccd1 vccd1 _14922_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14853_ _14861_/CLK _14853_/D vssd1 vssd1 vccd1 vccd1 _14853_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13804_ _15372_/CLK _13804_/D vssd1 vssd1 vccd1 vccd1 _13804_/Q sky130_fd_sc_hd__dfxtp_4
X_14784_ _15354_/CLK _14784_/D vssd1 vssd1 vccd1 vccd1 _14784_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11996_ _11979_/X _11980_/X _12260_/A vssd1 vssd1 vccd1 vccd1 _11996_/X sky130_fd_sc_hd__mux2_1
XFILLER_32_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13735_ _15537_/CLK _13735_/D vssd1 vssd1 vccd1 vccd1 _13735_/Q sky130_fd_sc_hd__dfxtp_1
X_10947_ _14958_/Q _10948_/B _10946_/Y _13242_/B vssd1 vssd1 vccd1 vccd1 _14958_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_45_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13666_ _15641_/CLK _13666_/D vssd1 vssd1 vccd1 vccd1 _13666_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10878_ _14910_/Q _15541_/Q _13134_/A vssd1 vssd1 vccd1 vccd1 _14910_/D sky130_fd_sc_hd__mux2_1
X_15405_ _15646_/CLK _15405_/D vssd1 vssd1 vccd1 vccd1 _15405_/Q sky130_fd_sc_hd__dfxtp_2
XPHY_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12617_ _12600_/X _12601_/X _12617_/S vssd1 vssd1 vccd1 vccd1 _12617_/X sky130_fd_sc_hd__mux2_1
X_13597_ _15354_/CLK _13597_/D vssd1 vssd1 vccd1 vccd1 _13597_/Q sky130_fd_sc_hd__dfxtp_2
Xclkbuf_4_14_0_clk clkbuf_3_7_0_clk/X vssd1 vssd1 vccd1 vccd1 clkbuf_5_29_0_clk/A
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_129_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15336_ _15336_/CLK _15336_/D vssd1 vssd1 vccd1 vccd1 _15336_/Q sky130_fd_sc_hd__dfxtp_1
X_12548_ _12531_/X _12532_/X _12548_/S vssd1 vssd1 vccd1 vccd1 _12548_/X sky130_fd_sc_hd__mux2_1
XFILLER_129_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15267_ _15267_/CLK _15267_/D vssd1 vssd1 vccd1 vccd1 _15267_/Q sky130_fd_sc_hd__dfxtp_1
X_12479_ _12462_/X _12463_/X _12490_/A vssd1 vssd1 vccd1 vccd1 _12479_/X sky130_fd_sc_hd__mux2_1
XANTENNA_2 _07319_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14218_ _15679_/CLK _14218_/D vssd1 vssd1 vccd1 vccd1 _14218_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_172_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15198_ _15675_/CLK _15198_/D vssd1 vssd1 vccd1 vccd1 _15198_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14149_ _15667_/CLK _14149_/D vssd1 vssd1 vccd1 vccd1 _14149_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout509 _07498_/C vssd1 vssd1 vccd1 vccd1 _07482_/C sky130_fd_sc_hd__buf_8
XFILLER_101_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06971_ _06708_/Y _13499_/Q _06710_/Y _13498_/Q vssd1 vssd1 vccd1 vccd1 _06971_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_100_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_1013 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08710_ _13800_/Q _12878_/S _08709_/X vssd1 vssd1 vccd1 vccd1 _13800_/D sky130_fd_sc_hd__o21a_1
XTAP_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09690_ _14061_/Q _13104_/B2 _09690_/S vssd1 vssd1 vccd1 vccd1 _14061_/D sky130_fd_sc_hd__mux2_1
XFILLER_117_1091 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08641_ _13524_/Q _08683_/A2 _08691_/B1 _13492_/Q _08640_/X vssd1 vssd1 vccd1 vccd1
+ _08645_/B sky130_fd_sc_hd__a221o_1
XFILLER_66_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08572_ _14512_/Q _08748_/B1 _08569_/X _08570_/X _08571_/X vssd1 vssd1 vccd1 vccd1
+ _08572_/X sky130_fd_sc_hd__a2111o_1
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_187_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07523_ _14753_/Q _13432_/Q _07529_/S vssd1 vssd1 vccd1 vccd1 _13432_/D sky130_fd_sc_hd__mux2_1
XFILLER_41_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_179_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07454_ _14665_/Q _07490_/B _14710_/Q vssd1 vssd1 vccd1 vccd1 _07454_/X sky130_fd_sc_hd__and3_1
XFILLER_34_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_520 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07385_ _11854_/A1 _13385_/Q _07501_/S vssd1 vssd1 vccd1 vccd1 _13385_/D sky130_fd_sc_hd__mux2_1
XFILLER_22_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09124_ _13950_/Q _13692_/Q _09230_/S vssd1 vssd1 vccd1 vccd1 _09124_/X sky130_fd_sc_hd__mux2_1
XFILLER_182_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09055_ _13914_/Q _09054_/X _13138_/S vssd1 vssd1 vccd1 vccd1 _13914_/D sky130_fd_sc_hd__mux2_1
XFILLER_135_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08006_ _13568_/Q _13567_/Q _13566_/Q _08006_/D vssd1 vssd1 vccd1 vccd1 _08017_/D
+ sky130_fd_sc_hd__and4_2
XFILLER_151_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09957_ _11877_/A1 _14317_/Q _09958_/S vssd1 vssd1 vccd1 vccd1 _14317_/D sky130_fd_sc_hd__mux2_1
XFILLER_103_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_1090 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08908_ _13123_/A _08907_/X _08906_/X _09382_/A vssd1 vssd1 vccd1 vccd1 _08908_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09888_ _11874_/A1 _14250_/Q _09897_/S vssd1 vssd1 vccd1 vccd1 _14250_/D sky130_fd_sc_hd__mux2_1
XFILLER_58_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_607 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08839_ _13862_/Q _11838_/A1 _08851_/S vssd1 vssd1 vccd1 vccd1 _13862_/D sky130_fd_sc_hd__mux2_1
XFILLER_79_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11850_ _15272_/Q _11883_/A1 _11850_/S vssd1 vssd1 vccd1 vccd1 _15272_/D sky130_fd_sc_hd__mux2_1
XTAP_2724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10801_ _14833_/Q _07339_/X _12481_/A vssd1 vssd1 vccd1 vccd1 _14833_/D sky130_fd_sc_hd__mux2_1
XTAP_2757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11781_ _11781_/A vssd1 vssd1 vccd1 vccd1 _11781_/Y sky130_fd_sc_hd__inv_2
XTAP_2779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13520_ _15379_/CLK _13520_/D vssd1 vssd1 vccd1 vccd1 _13520_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10732_ _15025_/Q _10569_/B _10602_/B _15042_/Q _10732_/C1 vssd1 vssd1 vccd1 vccd1
+ _10732_/X sky130_fd_sc_hd__a221o_1
XFILLER_158_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13451_ _15374_/CLK _13451_/D vssd1 vssd1 vccd1 vccd1 _13451_/Q sky130_fd_sc_hd__dfxtp_2
X_10663_ _15028_/Q _10602_/B _10662_/X vssd1 vssd1 vccd1 vccd1 _10663_/X sky130_fd_sc_hd__a21o_1
XFILLER_139_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12402_ _12406_/A _12402_/B vssd1 vssd1 vccd1 vccd1 _12402_/X sky130_fd_sc_hd__and2_1
XFILLER_40_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13382_ _14485_/Q vssd1 vssd1 vccd1 vccd1 _14485_/D sky130_fd_sc_hd__clkbuf_2
X_10594_ _10591_/X _10592_/X _10593_/X _10734_/A2 _15046_/Q vssd1 vssd1 vccd1 vccd1
+ _10594_/X sky130_fd_sc_hd__o32a_2
XFILLER_127_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15121_ _15659_/CLK _15121_/D vssd1 vssd1 vccd1 vccd1 _15121_/Q sky130_fd_sc_hd__dfxtp_1
X_12333_ _12544_/A _12333_/B vssd1 vssd1 vccd1 vccd1 _12333_/X sky130_fd_sc_hd__and2_1
XFILLER_182_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_3_3_0_clk clkbuf_3_3_0_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_7_0_clk/A sky130_fd_sc_hd__clkbuf_8
X_15052_ _15054_/CLK _15052_/D vssd1 vssd1 vccd1 vccd1 _15052_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_154_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12264_ _12268_/A _12264_/B vssd1 vssd1 vccd1 vccd1 _12264_/X sky130_fd_sc_hd__and2_1
XFILLER_141_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14003_ _14470_/CLK _14003_/D vssd1 vssd1 vccd1 vccd1 _14003_/Q sky130_fd_sc_hd__dfxtp_1
X_11215_ _10390_/C _15004_/Q _11232_/S vssd1 vssd1 vccd1 vccd1 _15004_/D sky130_fd_sc_hd__mux2_1
X_12195_ _12498_/A _12195_/B vssd1 vssd1 vccd1 vccd1 _12195_/X sky130_fd_sc_hd__and2_1
Xoutput50 _07186_/X vssd1 vssd1 vccd1 vccd1 ext_address[24] sky130_fd_sc_hd__clkbuf_2
XFILLER_134_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput61 _07167_/X vssd1 vssd1 vccd1 vccd1 ext_address[5] sky130_fd_sc_hd__clkbuf_2
Xoutput72 _07129_/X vssd1 vssd1 vccd1 vccd1 ext_write_data[14] sky130_fd_sc_hd__clkbuf_2
X_11146_ _11199_/A _11193_/B vssd1 vssd1 vccd1 vccd1 _11146_/Y sky130_fd_sc_hd__nand2_1
Xoutput83 _07149_/X vssd1 vssd1 vccd1 vccd1 ext_write_data[24] sky130_fd_sc_hd__clkbuf_2
Xoutput94 _07113_/X vssd1 vssd1 vccd1 vccd1 ext_write_data[5] sky130_fd_sc_hd__clkbuf_2
XFILLER_150_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11077_ _11074_/X _11076_/X _11362_/B vssd1 vssd1 vccd1 vccd1 _11077_/X sky130_fd_sc_hd__mux2_1
X_10028_ _11816_/A1 _14386_/Q _10028_/S vssd1 vssd1 vccd1 vccd1 _14386_/D sky130_fd_sc_hd__mux2_1
XFILLER_48_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14905_ _15499_/CLK _14905_/D vssd1 vssd1 vccd1 vccd1 _14905_/Q sky130_fd_sc_hd__dfxtp_2
Xclkbuf_leaf_196_clk clkbuf_5_17_0_clk/X vssd1 vssd1 vccd1 vccd1 _14373_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_64_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14836_ _15536_/CLK _14836_/D vssd1 vssd1 vccd1 vccd1 _14836_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_91_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14767_ _14861_/CLK _14767_/D vssd1 vssd1 vccd1 vccd1 _14767_/Q sky130_fd_sc_hd__dfxtp_4
X_11979_ _14522_/Q _14135_/Q _14167_/Q _14103_/Q _11993_/S _11992_/A vssd1 vssd1 vccd1
+ vccd1 _11979_/X sky130_fd_sc_hd__mux4_1
XFILLER_17_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13718_ _14997_/CLK _13718_/D vssd1 vssd1 vccd1 vccd1 _13718_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_177_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14698_ _15624_/CLK _14698_/D vssd1 vssd1 vccd1 vccd1 _14698_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_177_637 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13649_ _15434_/CLK _13649_/D vssd1 vssd1 vccd1 vccd1 _13649_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07170_ _15344_/Q _15051_/Q _07188_/S vssd1 vssd1 vccd1 vccd1 _07170_/X sky130_fd_sc_hd__mux2_8
XFILLER_173_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15319_ _15332_/CLK _15319_/D vssd1 vssd1 vccd1 vccd1 _15319_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_120_clk clkbuf_5_30_0_clk/X vssd1 vssd1 vccd1 vccd1 _15389_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_172_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_792 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout306 _13092_/B2 vssd1 vssd1 vccd1 vccd1 _13339_/A0 sky130_fd_sc_hd__clkbuf_4
XFILLER_114_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09811_ _14177_/Q _13333_/A0 _09823_/S vssd1 vssd1 vccd1 vccd1 _14177_/D sky130_fd_sc_hd__mux2_1
XFILLER_87_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout317 _13082_/B2 vssd1 vssd1 vccd1 vccd1 _13334_/A0 sky130_fd_sc_hd__buf_6
XFILLER_154_1055 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout328 _07416_/X vssd1 vssd1 vccd1 vccd1 _13072_/B2 sky130_fd_sc_hd__clkbuf_16
Xfanout339 _07396_/X vssd1 vssd1 vccd1 vccd1 _13324_/A0 sky130_fd_sc_hd__buf_6
XFILLER_140_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_103 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09742_ _14110_/Q _13074_/B2 _09757_/S vssd1 vssd1 vccd1 vccd1 _14110_/D sky130_fd_sc_hd__mux2_1
X_06954_ _06892_/X _06932_/X _06945_/Y _06951_/X _06953_/X vssd1 vssd1 vccd1 vccd1
+ _06954_/X sky130_fd_sc_hd__a2111o_2
X_09673_ _14044_/Q _13328_/A0 _09690_/S vssd1 vssd1 vccd1 vccd1 _14044_/D sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_187_clk clkbuf_5_21_0_clk/X vssd1 vssd1 vccd1 vccd1 _15669_/CLK sky130_fd_sc_hd__clkbuf_16
X_06885_ _15396_/Q _06696_/Y _15395_/Q _06699_/Y vssd1 vssd1 vccd1 vccd1 _06929_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_27_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08624_ _13431_/Q _08736_/A2 _08748_/B1 _14504_/Q vssd1 vssd1 vccd1 vccd1 _08624_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_43_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08555_ _13537_/Q _08750_/A2 _08747_/B1 _13505_/Q _08554_/X vssd1 vssd1 vccd1 vccd1
+ _08559_/B sky130_fd_sc_hd__a221o_1
X_07506_ _14736_/Q _13415_/Q _07535_/S vssd1 vssd1 vccd1 vccd1 _13415_/D sky130_fd_sc_hd__mux2_1
X_08486_ _13772_/Q _08485_/X _12906_/S vssd1 vssd1 vccd1 vccd1 _13772_/D sky130_fd_sc_hd__mux2_1
XFILLER_51_974 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07437_ _13334_/A0 _13398_/Q _07481_/S vssd1 vssd1 vccd1 vccd1 _13398_/D sky130_fd_sc_hd__mux2_1
XFILLER_50_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07368_ _14713_/Q _08817_/B vssd1 vssd1 vccd1 vccd1 _08852_/B sky130_fd_sc_hd__nand2_4
XFILLER_149_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09107_ _09427_/A1 _09105_/X _09106_/X vssd1 vssd1 vccd1 vccd1 _09107_/X sky130_fd_sc_hd__a21o_1
XFILLER_182_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_111_clk _15447_/CLK vssd1 vssd1 vccd1 vccd1 _15354_/CLK sky130_fd_sc_hd__clkbuf_16
X_07299_ _07294_/Y _07295_/X _07297_/Y _07298_/X vssd1 vssd1 vccd1 vccd1 _07350_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_109_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09038_ _09221_/A _09038_/B vssd1 vssd1 vccd1 vccd1 _09038_/X sky130_fd_sc_hd__or2_1
XFILLER_163_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11000_ _10998_/Y _10999_/Y _11088_/S vssd1 vssd1 vccd1 vccd1 _11000_/X sky130_fd_sc_hd__mux2_1
XFILLER_117_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_795 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12951_ _10589_/X _14864_/Q _13038_/S vssd1 vssd1 vccd1 vccd1 _12951_/X sky130_fd_sc_hd__mux2_2
XTAP_3211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_178_clk clkbuf_5_22_0_clk/X vssd1 vssd1 vccd1 vccd1 _15324_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_3222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11902_ _12500_/A1 _11901_/X _12500_/B1 vssd1 vssd1 vccd1 vccd1 _11902_/X sky130_fd_sc_hd__a21o_1
XFILLER_93_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15670_ _15670_/CLK _15670_/D vssd1 vssd1 vccd1 vccd1 _15670_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12882_ _15410_/Q _15595_/Q _12885_/S vssd1 vssd1 vccd1 vccd1 _15410_/D sky130_fd_sc_hd__mux2_1
XTAP_3255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14621_ _14774_/CLK _14621_/D vssd1 vssd1 vccd1 vccd1 _14621_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_93_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11833_ _15255_/Q _13080_/B2 _11849_/S vssd1 vssd1 vccd1 vccd1 _15255_/D sky130_fd_sc_hd__mux2_1
XTAP_2554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14552_ _15275_/CLK _14552_/D vssd1 vssd1 vccd1 vccd1 _14552_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11764_ _13339_/A0 _15192_/Q _11775_/S vssd1 vssd1 vccd1 vccd1 _15192_/D sky130_fd_sc_hd__mux2_1
XTAP_1864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13503_ _14513_/CLK _13503_/D vssd1 vssd1 vccd1 vccd1 _13503_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_14_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10715_ _14761_/Q _10714_/X _10715_/S vssd1 vssd1 vccd1 vccd1 _14761_/D sky130_fd_sc_hd__mux2_1
XFILLER_13_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14483_ _15650_/CLK _14483_/D vssd1 vssd1 vccd1 vccd1 _14483_/Q sky130_fd_sc_hd__dfxtp_1
X_11695_ _13337_/A0 _15126_/Q _11708_/S vssd1 vssd1 vccd1 vccd1 _15126_/D sky130_fd_sc_hd__mux2_1
X_13434_ _14495_/CLK _13434_/D vssd1 vssd1 vccd1 vccd1 _13434_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10646_ _15567_/Q _10706_/B vssd1 vssd1 vccd1 vccd1 _10646_/X sky130_fd_sc_hd__and2_1
XFILLER_155_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_102_clk clkbuf_5_26_0_clk/X vssd1 vssd1 vccd1 vccd1 _15452_/CLK sky130_fd_sc_hd__clkbuf_16
X_13365_ _14468_/Q vssd1 vssd1 vccd1 vccd1 _14468_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_182_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10577_ _14962_/Q _10733_/A2 _10733_/B1 _14930_/Q _10574_/X vssd1 vssd1 vccd1 vccd1
+ _10577_/X sky130_fd_sc_hd__a221o_1
XFILLER_6_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15104_ _15259_/CLK _15104_/D vssd1 vssd1 vccd1 vccd1 _15104_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_170_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12316_ _12592_/A1 _12315_/X _12615_/B1 vssd1 vssd1 vccd1 vccd1 _12316_/X sky130_fd_sc_hd__a21o_1
XFILLER_142_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13296_ _12695_/X _15628_/Q _13300_/S vssd1 vssd1 vccd1 vccd1 _15628_/D sky130_fd_sc_hd__mux2_1
XFILLER_138_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15035_ _15041_/CLK _15035_/D vssd1 vssd1 vccd1 vccd1 _15035_/Q sky130_fd_sc_hd__dfxtp_1
X_12247_ _12477_/A1 _12246_/X _12468_/A1 vssd1 vssd1 vccd1 vccd1 _12247_/X sky130_fd_sc_hd__a21o_1
XFILLER_123_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12178_ _12477_/A1 _12177_/X _12468_/A1 vssd1 vssd1 vccd1 vccd1 _12178_/X sky130_fd_sc_hd__a21o_1
XFILLER_69_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11129_ _11129_/A _11129_/B vssd1 vssd1 vccd1 vccd1 _11129_/Y sky130_fd_sc_hd__nor2_4
XFILLER_95_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_169_clk clkbuf_5_23_0_clk/X vssd1 vssd1 vccd1 vccd1 _15161_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_95_189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06670_ _06670_/A vssd1 vssd1 vccd1 vccd1 _06670_/Y sky130_fd_sc_hd__inv_2
XFILLER_37_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1018 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14819_ _15638_/CLK _14819_/D vssd1 vssd1 vccd1 vccd1 _14819_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08340_ _13723_/Q _11346_/A2 _11351_/C1 _08339_/X vssd1 vssd1 vccd1 vccd1 _13723_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_177_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08271_ _07341_/A _10481_/B _08270_/X vssd1 vssd1 vccd1 vccd1 _13165_/B sky130_fd_sc_hd__a21oi_4
XFILLER_165_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07222_ _07206_/X _07208_/Y _07219_/X _07221_/Y _07218_/Y vssd1 vssd1 vccd1 vccd1
+ _07231_/B sky130_fd_sc_hd__a221o_1
XFILLER_165_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07153_ _07163_/A _07153_/B vssd1 vssd1 vccd1 vccd1 _07153_/X sky130_fd_sc_hd__and2_4
XFILLER_173_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07084_ _14640_/Q _14672_/Q _07096_/S vssd1 vssd1 vccd1 vccd1 _07084_/X sky130_fd_sc_hd__mux2_1
XFILLER_173_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout103 _12759_/B vssd1 vssd1 vccd1 vccd1 _12765_/B sky130_fd_sc_hd__clkbuf_16
Xfanout114 _13041_/Y vssd1 vssd1 vccd1 vccd1 _13042_/A sky130_fd_sc_hd__buf_8
Xfanout125 fanout138/X vssd1 vssd1 vccd1 vccd1 _13139_/S sky130_fd_sc_hd__buf_6
Xfanout136 _10765_/S vssd1 vssd1 vccd1 vccd1 _08722_/A sky130_fd_sc_hd__buf_12
XFILLER_59_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout147 _12320_/A vssd1 vssd1 vccd1 vccd1 _12904_/S sky130_fd_sc_hd__buf_12
Xfanout158 _08573_/S vssd1 vssd1 vccd1 vccd1 _12933_/S sky130_fd_sc_hd__clkbuf_16
X_07986_ _07995_/D _07985_/Y _07964_/A vssd1 vssd1 vccd1 vccd1 _07986_/Y sky130_fd_sc_hd__o21ai_1
Xfanout169 _11818_/Y vssd1 vssd1 vccd1 vccd1 _11849_/S sky130_fd_sc_hd__buf_12
X_09725_ _13347_/A0 _14095_/Q _09728_/S vssd1 vssd1 vccd1 vccd1 _14095_/D sky130_fd_sc_hd__mux2_1
X_06937_ _06736_/Y _13485_/Q _06738_/Y _13484_/Q _06936_/Y vssd1 vssd1 vccd1 vccd1
+ _06943_/A sky130_fd_sc_hd__o221a_1
XFILLER_80_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09656_ _14029_/Q _13104_/B2 _09660_/S vssd1 vssd1 vccd1 vccd1 _14029_/D sky130_fd_sc_hd__mux2_1
XFILLER_55_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06868_ _06872_/A _13508_/Q _06874_/A _13507_/Q vssd1 vssd1 vccd1 vccd1 _06882_/C
+ sky130_fd_sc_hd__a22o_1
X_08607_ _13465_/Q _08684_/A2 _08683_/A2 _13529_/Q vssd1 vssd1 vccd1 vccd1 _08607_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09587_ _13963_/Q _13343_/A0 _09589_/S vssd1 vssd1 vccd1 vccd1 _13963_/D sky130_fd_sc_hd__mux2_1
XTAP_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_226 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06799_ _06799_/A _08477_/C vssd1 vssd1 vccd1 vccd1 _08773_/A sky130_fd_sc_hd__or2_2
XFILLER_179_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08538_ _08538_/A _08538_/B vssd1 vssd1 vccd1 vccd1 _08538_/Y sky130_fd_sc_hd__nor2_4
XFILLER_23_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_771 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08469_ _08469_/A _08765_/D vssd1 vssd1 vccd1 vccd1 _08487_/B sky130_fd_sc_hd__or2_2
XFILLER_169_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10500_ _07244_/A _10523_/A2 _10499_/X vssd1 vssd1 vccd1 vccd1 _13220_/B sky130_fd_sc_hd__a21o_4
XFILLER_183_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11480_ _13199_/B _11480_/B vssd1 vssd1 vccd1 vccd1 _11481_/B sky130_fd_sc_hd__and2_1
XFILLER_155_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10431_ _10520_/A1 _13778_/Q _13746_/Q _10520_/B2 vssd1 vssd1 vccd1 vccd1 _10431_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_12_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13150_ _14610_/Q _15548_/Q _13154_/S vssd1 vssd1 vccd1 vccd1 _15548_/D sky130_fd_sc_hd__mux2_1
X_10362_ _14767_/Q _13791_/Q _13759_/Q _14766_/Q _10360_/X vssd1 vssd1 vccd1 vccd1
+ _10362_/X sky130_fd_sc_hd__a221o_4
X_12101_ _12273_/A1 _12096_/X _12099_/X _12100_/X _08449_/A vssd1 vssd1 vccd1 vccd1
+ _12113_/B sky130_fd_sc_hd__a221o_1
XFILLER_128_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13081_ _15508_/Q _13081_/A2 _13105_/B1 _13080_/X vssd1 vssd1 vccd1 vccd1 _15508_/D
+ sky130_fd_sc_hd__a22o_1
X_10293_ _14678_/Q _14863_/Q _10730_/S vssd1 vssd1 vccd1 vccd1 _14678_/D sky130_fd_sc_hd__mux2_1
XFILLER_152_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12032_ _12595_/A1 _12027_/X _12030_/X _12031_/X _08405_/D vssd1 vssd1 vccd1 vccd1
+ _12044_/B sky130_fd_sc_hd__a221o_1
XFILLER_2_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13983_ _15510_/CLK _13983_/D vssd1 vssd1 vccd1 vccd1 _13983_/Q sky130_fd_sc_hd__dfxtp_1
X_12934_ _14923_/Q _14902_/Q vssd1 vssd1 vccd1 vccd1 _12934_/Y sky130_fd_sc_hd__nand2_1
XTAP_3030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_565 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15653_ _15660_/CLK _15653_/D vssd1 vssd1 vccd1 vccd1 _15653_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12865_ _14759_/Q _15393_/Q _12866_/S vssd1 vssd1 vccd1 vccd1 _15393_/D sky130_fd_sc_hd__mux2_1
XTAP_3085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14604_ _15587_/CLK _14604_/D vssd1 vssd1 vccd1 vccd1 _14604_/Q sky130_fd_sc_hd__dfxtp_1
X_11816_ _15239_/Q _11816_/A1 _11816_/S vssd1 vssd1 vccd1 vccd1 _15239_/D sky130_fd_sc_hd__mux2_1
XTAP_2384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15584_ _15584_/CLK _15584_/D vssd1 vssd1 vccd1 vccd1 _15584_/Q sky130_fd_sc_hd__dfxtp_1
X_12796_ _15362_/Q _13309_/B vssd1 vssd1 vccd1 vccd1 _12810_/C sky130_fd_sc_hd__and2_2
XTAP_2395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_434 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14535_ _15125_/CLK _14535_/D vssd1 vssd1 vccd1 vccd1 _14535_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11747_ _13322_/A0 _15175_/Q _11774_/S vssd1 vssd1 vccd1 vccd1 _15175_/D sky130_fd_sc_hd__mux2_1
XFILLER_30_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_467 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14466_ _14525_/CLK _14466_/D vssd1 vssd1 vccd1 vccd1 _14466_/Q sky130_fd_sc_hd__dfxtp_1
X_11678_ _11853_/A1 _15109_/Q _11708_/S vssd1 vssd1 vccd1 vccd1 _15109_/D sky130_fd_sc_hd__mux2_1
XFILLER_146_128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13417_ _13803_/CLK _13417_/D vssd1 vssd1 vccd1 vccd1 _13417_/Q sky130_fd_sc_hd__dfxtp_2
X_10629_ _15053_/Q _10714_/A2 _10626_/X _10628_/X vssd1 vssd1 vccd1 vccd1 _10629_/X
+ sky130_fd_sc_hd__o22a_2
X_14397_ _15652_/CLK _14397_/D vssd1 vssd1 vccd1 vccd1 _14397_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_155_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13348_ _13348_/A0 _15678_/Q _13350_/S vssd1 vssd1 vccd1 vccd1 _15678_/D sky130_fd_sc_hd__mux2_1
XFILLER_115_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13279_ _15363_/Q _15610_/Q _13309_/A vssd1 vssd1 vccd1 vccd1 _15610_/D sky130_fd_sc_hd__mux2_1
XFILLER_5_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15018_ _15020_/CLK _15018_/D vssd1 vssd1 vccd1 vccd1 _15018_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_97_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07840_ _13524_/Q _07847_/D vssd1 vssd1 vccd1 vccd1 _07844_/B sky130_fd_sc_hd__nand2_1
XFILLER_110_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07771_ _14763_/Q _07777_/A _07770_/Y _08012_/C1 vssd1 vssd1 vccd1 vccd1 _13506_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_110_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09510_ _09524_/A _09510_/B _09510_/C vssd1 vssd1 vccd1 vccd1 _09510_/X sky130_fd_sc_hd__and3_1
XFILLER_65_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06722_ _13492_/Q vssd1 vssd1 vccd1 vccd1 _06936_/B sky130_fd_sc_hd__inv_2
XFILLER_92_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09441_ _14029_/Q _13997_/Q _09441_/S vssd1 vssd1 vccd1 vccd1 _09441_/X sky130_fd_sc_hd__mux2_1
XFILLER_80_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09372_ _06675_/Y _09369_/X _09371_/X _09382_/A vssd1 vssd1 vccd1 vccd1 _09372_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_178_710 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08323_ _11025_/A _11419_/A vssd1 vssd1 vccd1 vccd1 _11045_/B sky130_fd_sc_hd__nor2_1
XFILLER_20_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_607 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08254_ _07329_/A _10481_/B _08253_/X vssd1 vssd1 vccd1 vccd1 _13159_/B sky130_fd_sc_hd__a21o_4
X_07205_ _07228_/A _07228_/B _07202_/X _07204_/Y vssd1 vssd1 vccd1 vccd1 _07205_/X
+ sky130_fd_sc_hd__a22o_1
X_08185_ _08185_/A _08185_/B vssd1 vssd1 vccd1 vccd1 _08185_/X sky130_fd_sc_hd__and2_1
XFILLER_180_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07136_ _14848_/Q _14840_/Q _07146_/S vssd1 vssd1 vccd1 vccd1 _07136_/X sky130_fd_sc_hd__mux2_1
XFILLER_106_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07067_ _07066_/X _13601_/Q _12764_/S vssd1 vssd1 vccd1 vccd1 _07067_/X sky130_fd_sc_hd__mux2_1
XFILLER_133_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07969_ _14750_/Q _07971_/A _07968_/X _07987_/C1 vssd1 vssd1 vccd1 vccd1 _13557_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_87_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09708_ _13074_/B2 _14078_/Q _09723_/S vssd1 vssd1 vccd1 vccd1 _14078_/D sky130_fd_sc_hd__mux2_1
X_10980_ _11356_/B _10978_/X _10979_/X vssd1 vssd1 vccd1 vccd1 _10980_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_83_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09639_ _14012_/Q _13328_/A0 _09660_/S vssd1 vssd1 vccd1 vccd1 _14012_/D sky130_fd_sc_hd__mux2_1
XFILLER_167_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12650_ _15341_/Q _12759_/B _12649_/X _12832_/C1 vssd1 vssd1 vccd1 vccd1 _15341_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_70_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_64 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11601_ _13236_/B _11602_/B vssd1 vssd1 vccd1 vccd1 _11611_/A sky130_fd_sc_hd__and2_1
X_12581_ _15303_/Q _15271_/Q _15239_/Q _15170_/Q _12453_/S _12452_/A vssd1 vssd1 vccd1
+ vccd1 _12582_/B sky130_fd_sc_hd__mux4_1
XFILLER_169_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14320_ _15291_/CLK _14320_/D vssd1 vssd1 vccd1 vccd1 _14320_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11532_ _13215_/B _11532_/B vssd1 vssd1 vccd1 vccd1 _11533_/B sky130_fd_sc_hd__or2_1
XFILLER_184_724 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_183_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14251_ _15527_/CLK _14251_/D vssd1 vssd1 vccd1 vccd1 _14251_/Q sky130_fd_sc_hd__dfxtp_1
X_11463_ _11464_/B _11464_/C _11505_/A vssd1 vssd1 vccd1 vccd1 _11472_/B sky130_fd_sc_hd__o21a_1
XFILLER_139_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13202_ _13233_/A _13202_/B vssd1 vssd1 vccd1 vccd1 _13202_/X sky130_fd_sc_hd__or2_1
X_10414_ _08313_/Y _11436_/A _10382_/B _11436_/B _13183_/B vssd1 vssd1 vccd1 vccd1
+ _10414_/X sky130_fd_sc_hd__o32a_1
XFILLER_137_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14182_ _14537_/CLK _14182_/D vssd1 vssd1 vccd1 vccd1 _14182_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_104_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11394_ _11394_/A _11394_/B vssd1 vssd1 vccd1 vccd1 _11394_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_99_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13133_ _14608_/Q _14609_/Q _13133_/C vssd1 vssd1 vccd1 vccd1 _13134_/C sky130_fd_sc_hd__nor3_1
XFILLER_136_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10345_ _14929_/D _14928_/D _14927_/D vssd1 vssd1 vccd1 vccd1 _10560_/S sky130_fd_sc_hd__and3b_1
XFILLER_87_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13064_ _12963_/X _13118_/A2 _13104_/B1 _07400_/X vssd1 vssd1 vccd1 vccd1 _13064_/X
+ sky130_fd_sc_hd__a22o_1
X_10276_ _14661_/Q _14814_/Q _10650_/S vssd1 vssd1 vccd1 vccd1 _14661_/D sky130_fd_sc_hd__mux2_1
XFILLER_79_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12015_ _12590_/A _12015_/B vssd1 vssd1 vccd1 vccd1 _12015_/X sky130_fd_sc_hd__and2_1
XFILLER_94_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13966_ _15334_/CLK _13966_/D vssd1 vssd1 vccd1 vccd1 _13966_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_46_351 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12917_ _15445_/Q _15631_/Q _12917_/S vssd1 vssd1 vccd1 vccd1 _15445_/D sky130_fd_sc_hd__mux2_1
XFILLER_34_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13897_ _15130_/CLK _13897_/D vssd1 vssd1 vccd1 vccd1 _13897_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_192 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15636_ _15636_/CLK _15636_/D vssd1 vssd1 vccd1 vccd1 _15636_/Q sky130_fd_sc_hd__dfxtp_1
X_12848_ _14742_/Q _15376_/Q _12866_/S vssd1 vssd1 vccd1 vccd1 _15376_/D sky130_fd_sc_hd__mux2_1
XTAP_2170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15567_ _15569_/CLK _15567_/D vssd1 vssd1 vccd1 vccd1 _15567_/Q sky130_fd_sc_hd__dfxtp_1
X_12779_ _15066_/Q _12792_/B vssd1 vssd1 vccd1 vccd1 _12779_/X sky130_fd_sc_hd__or2_1
XTAP_1480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14518_ _15108_/CLK _14518_/D vssd1 vssd1 vccd1 vccd1 _14518_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_148_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15498_ _15507_/CLK _15498_/D vssd1 vssd1 vccd1 vccd1 _15498_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14449_ _15199_/CLK _14449_/D vssd1 vssd1 vccd1 vccd1 _14449_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09990_ _11877_/A1 _14349_/Q _09991_/S vssd1 vssd1 vccd1 vccd1 _14349_/D sky130_fd_sc_hd__mux2_1
XFILLER_170_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_171_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08941_ _14069_/Q _13123_/B _08512_/B _14037_/Q _09543_/A vssd1 vssd1 vccd1 vccd1
+ _08941_/X sky130_fd_sc_hd__a221o_1
XFILLER_142_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08872_ _13893_/Q _13337_/A0 _08885_/S vssd1 vssd1 vccd1 vccd1 _13893_/D sky130_fd_sc_hd__mux2_1
XFILLER_57_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07823_ _07821_/X _07822_/Y _07830_/A vssd1 vssd1 vccd1 vccd1 _07823_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_28_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_115 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07754_ _07752_/Y _07756_/B _07750_/A vssd1 vssd1 vccd1 vccd1 _07754_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_25_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06705_ _13501_/Q vssd1 vssd1 vccd1 vccd1 _06705_/Y sky130_fd_sc_hd__inv_2
X_07685_ _14740_/Q _07676_/A _07684_/Y _07938_/C1 vssd1 vssd1 vccd1 vccd1 _13483_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_52_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_91_clk clkbuf_5_13_0_clk/X vssd1 vssd1 vccd1 vccd1 _15434_/CLK sky130_fd_sc_hd__clkbuf_16
X_09424_ _09427_/A1 _09422_/X _09423_/X vssd1 vssd1 vccd1 vccd1 _09424_/X sky130_fd_sc_hd__a21o_1
XFILLER_52_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09355_ _14476_/Q _09558_/A2 _09354_/X _13049_/A1 vssd1 vssd1 vccd1 vccd1 _09355_/X
+ sky130_fd_sc_hd__a211o_1
X_08306_ _08288_/X _08305_/X _11088_/S vssd1 vssd1 vccd1 vccd1 _08307_/B sky130_fd_sc_hd__mux2_1
XFILLER_165_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09286_ _13123_/A _09285_/X _09284_/X _09554_/A vssd1 vssd1 vccd1 vccd1 _09286_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_60_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08237_ _08237_/A _13773_/Q vssd1 vssd1 vccd1 vccd1 _08237_/X sky130_fd_sc_hd__and2_2
XFILLER_119_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08168_ _13671_/Q _10695_/S _08155_/X _08167_/X vssd1 vssd1 vccd1 vccd1 _13671_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_146_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07119_ _07131_/A _07119_/B vssd1 vssd1 vccd1 vccd1 _07119_/X sky130_fd_sc_hd__and2_4
X_08099_ input12/X input32/X input9/X input18/X _08150_/S _08151_/S vssd1 vssd1 vccd1
+ vccd1 _08099_/X sky130_fd_sc_hd__mux4_1
XFILLER_109_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10130_ _14516_/Q _14764_/Q _10131_/S vssd1 vssd1 vccd1 vccd1 _14516_/D sky130_fd_sc_hd__mux2_1
XFILLER_106_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10061_ _14418_/Q _13347_/A0 _10064_/S vssd1 vssd1 vccd1 vccd1 _14418_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_5_20_0_clk clkbuf_5_21_0_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_5_20_0_clk/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_134_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13820_ _15218_/CLK _13820_/D vssd1 vssd1 vccd1 vccd1 _13820_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13751_ _14703_/CLK _13751_/D vssd1 vssd1 vccd1 vccd1 _13751_/Q sky130_fd_sc_hd__dfxtp_1
X_10963_ _10963_/A _10963_/B vssd1 vssd1 vccd1 vccd1 _10963_/Y sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_82_clk clkbuf_5_15_0_clk/X vssd1 vssd1 vccd1 vccd1 _15422_/CLK sky130_fd_sc_hd__clkbuf_16
X_12702_ _15348_/Q _15347_/Q _12688_/B _15349_/Q vssd1 vssd1 vccd1 vccd1 _12703_/B
+ sky130_fd_sc_hd__a31o_1
X_13682_ _15334_/CLK _13682_/D vssd1 vssd1 vccd1 vccd1 _13682_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10894_ _14927_/D _14928_/D _14929_/D vssd1 vssd1 vccd1 vccd1 _10894_/X sky130_fd_sc_hd__and3b_4
XFILLER_188_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15421_ _15606_/CLK _15421_/D vssd1 vssd1 vccd1 vccd1 _15421_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_70_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12633_ _12743_/A _12633_/B vssd1 vssd1 vccd1 vccd1 _12633_/X sky130_fd_sc_hd__or2_1
XFILLER_141_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15352_ _15630_/CLK _15352_/D vssd1 vssd1 vccd1 vccd1 _15352_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_8_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12564_ _13904_/Q _14419_/Q _12568_/S vssd1 vssd1 vccd1 vccd1 _12564_/X sky130_fd_sc_hd__mux2_1
XFILLER_180_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14303_ _15181_/CLK _14303_/D vssd1 vssd1 vccd1 vccd1 _14303_/Q sky130_fd_sc_hd__dfxtp_1
X_11515_ _11512_/X _11515_/B vssd1 vssd1 vccd1 vccd1 _11546_/B sky130_fd_sc_hd__and2b_1
XFILLER_7_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15283_ _15662_/CLK _15283_/D vssd1 vssd1 vccd1 vccd1 _15283_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_184_565 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12495_ _13901_/Q _14416_/Q _12499_/S vssd1 vssd1 vccd1 vccd1 _12495_/X sky130_fd_sc_hd__mux2_1
X_14234_ _15178_/CLK _14234_/D vssd1 vssd1 vccd1 vccd1 _14234_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11446_ _11476_/B _11476_/C _13229_/A vssd1 vssd1 vccd1 vccd1 _11447_/B sky130_fd_sc_hd__a21oi_1
XFILLER_50_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_171_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14165_ _15654_/CLK _14165_/D vssd1 vssd1 vccd1 vccd1 _14165_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_166_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11377_ _11377_/A _11377_/B vssd1 vssd1 vccd1 vccd1 _11378_/B sky130_fd_sc_hd__nor2_1
XFILLER_153_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13116_ _12944_/A _13116_/B _13116_/C vssd1 vssd1 vccd1 vccd1 _13116_/X sky130_fd_sc_hd__and3b_1
XTAP_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10328_ _14906_/Q _14713_/Q _10566_/B vssd1 vssd1 vccd1 vccd1 _14713_/D sky130_fd_sc_hd__mux2_1
XFILLER_113_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14096_ _15226_/CLK _14096_/D vssd1 vssd1 vccd1 vccd1 _14096_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13047_ _13049_/A1 _13318_/C _09662_/B _08910_/S vssd1 vssd1 vccd1 vccd1 _13050_/B
+ sky130_fd_sc_hd__a22oi_1
X_10259_ _14644_/Q _14797_/Q _10343_/S vssd1 vssd1 vccd1 vccd1 _14644_/D sky130_fd_sc_hd__mux2_1
XFILLER_79_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14998_ _15556_/CLK _14998_/D vssd1 vssd1 vccd1 vccd1 _14998_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_693 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13949_ _15331_/CLK _13949_/D vssd1 vssd1 vccd1 vccd1 _13949_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_73_clk clkbuf_5_14_0_clk/X vssd1 vssd1 vccd1 vccd1 _15592_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_62_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07470_ _14669_/Q _07474_/B _07482_/C vssd1 vssd1 vccd1 vccd1 _07470_/X sky130_fd_sc_hd__and3_1
XFILLER_62_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_151 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_2_1_1_clk clkbuf_2_1_1_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_3_0_clk/A sky130_fd_sc_hd__clkbuf_8
X_15619_ _15619_/CLK _15619_/D vssd1 vssd1 vccd1 vccd1 _15619_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_882 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09140_ _15285_/Q _15253_/Q _15221_/Q _15152_/Q _09132_/S _09427_/A1 vssd1 vssd1
+ vccd1 vccd1 _09140_/X sky130_fd_sc_hd__mux4_1
XFILLER_148_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09071_ _09445_/C1 _09068_/X _09070_/X _09130_/A vssd1 vssd1 vccd1 vccd1 _09071_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_147_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08022_ _14765_/Q _08022_/B vssd1 vssd1 vccd1 vccd1 _08022_/Y sky130_fd_sc_hd__nor2_1
XFILLER_135_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_771 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09973_ _11860_/A1 _14332_/Q _09991_/S vssd1 vssd1 vccd1 vccd1 _14332_/D sky130_fd_sc_hd__mux2_1
XFILLER_103_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08924_ _15109_/Q _09558_/A2 _08540_/B _15077_/Q _08923_/X vssd1 vssd1 vccd1 vccd1
+ _08924_/X sky130_fd_sc_hd__a221o_1
XFILLER_162_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08855_ _13876_/Q _11853_/A1 _08885_/S vssd1 vssd1 vccd1 vccd1 _13876_/D sky130_fd_sc_hd__mux2_1
XTAP_3607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07806_ _13515_/Q _07813_/D vssd1 vssd1 vccd1 vccd1 _07810_/B sky130_fd_sc_hd__nand2_1
XTAP_3629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08786_ _13320_/A0 _13812_/Q _08816_/S vssd1 vssd1 vccd1 vccd1 _13812_/D sky130_fd_sc_hd__mux2_1
XTAP_2906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07737_ _14754_/Q _07736_/A _07736_/Y _08002_/C1 vssd1 vssd1 vccd1 vccd1 _13497_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_2928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_64_clk clkbuf_5_11_0_clk/X vssd1 vssd1 vccd1 vccd1 _15570_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_53_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07668_ _13479_/Q _07672_/C vssd1 vssd1 vccd1 vccd1 _07669_/B sky130_fd_sc_hd__xnor2_1
XFILLER_13_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09407_ _15673_/Q _13407_/Q _09407_/S vssd1 vssd1 vccd1 vccd1 _09407_/X sky130_fd_sc_hd__mux2_1
XFILLER_186_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07599_ _13461_/Q _07599_/B vssd1 vssd1 vccd1 vccd1 _07600_/B sky130_fd_sc_hd__xnor2_1
XFILLER_187_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_99 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09338_ _14088_/Q _13123_/B _08512_/B _14056_/Q _09466_/A vssd1 vssd1 vccd1 vccd1
+ _09338_/X sky130_fd_sc_hd__a221o_1
XFILLER_21_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09269_ _13957_/Q _13699_/Q _09557_/S vssd1 vssd1 vccd1 vccd1 _09269_/X sky130_fd_sc_hd__mux2_1
XFILLER_166_565 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11300_ _11414_/A _08309_/Y _11298_/Y _11299_/Y wire438/X vssd1 vssd1 vccd1 vccd1
+ _11300_/X sky130_fd_sc_hd__o221a_1
XFILLER_154_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12280_ _12276_/X _12277_/X _12536_/A vssd1 vssd1 vccd1 vccd1 _12280_/X sky130_fd_sc_hd__mux2_1
XFILLER_181_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11231_ _10470_/D _15019_/Q _11232_/S vssd1 vssd1 vccd1 vccd1 _15019_/D sky130_fd_sc_hd__mux2_1
XFILLER_101_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_985 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11162_ _11371_/A _11112_/X _11199_/A vssd1 vssd1 vccd1 vccd1 _11162_/X sky130_fd_sc_hd__a21o_1
XFILLER_45_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10113_ _14499_/Q _14747_/Q _10124_/S vssd1 vssd1 vccd1 vccd1 _14499_/D sky130_fd_sc_hd__mux2_1
XFILLER_1_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11093_ _10959_/Y _10980_/Y _11115_/S vssd1 vssd1 vccd1 vccd1 _11093_/X sky130_fd_sc_hd__mux2_2
X_10044_ _14401_/Q _13074_/B2 _10059_/S vssd1 vssd1 vccd1 vccd1 _14401_/D sky130_fd_sc_hd__mux2_1
X_14921_ _15552_/CLK _14921_/D vssd1 vssd1 vccd1 vccd1 _14921_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14852_ _15500_/CLK _14852_/D vssd1 vssd1 vccd1 vccd1 _14852_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_1080 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13803_ _13803_/CLK _13803_/D vssd1 vssd1 vccd1 vccd1 _13803_/Q sky130_fd_sc_hd__dfxtp_2
X_14783_ _15634_/CLK _14783_/D vssd1 vssd1 vccd1 vccd1 _14783_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11995_ _11988_/X _11990_/X _11992_/X _11994_/X _12501_/C1 vssd1 vssd1 vccd1 vccd1
+ _11995_/X sky130_fd_sc_hd__o221a_1
XFILLER_63_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_55_clk clkbuf_5_11_0_clk/X vssd1 vssd1 vccd1 vccd1 _15582_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_16_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13734_ _15530_/CLK _13734_/D vssd1 vssd1 vccd1 vccd1 _13734_/Q sky130_fd_sc_hd__dfxtp_1
X_10946_ _11616_/A _10948_/B vssd1 vssd1 vccd1 vccd1 _10946_/Y sky130_fd_sc_hd__nand2_1
XFILLER_16_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_663 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13665_ _15606_/CLK _13665_/D vssd1 vssd1 vccd1 vccd1 _13665_/Q sky130_fd_sc_hd__dfxtp_1
X_10877_ _13729_/Q _14909_/Q _10877_/S vssd1 vssd1 vccd1 vccd1 _14909_/D sky130_fd_sc_hd__mux2_1
XFILLER_188_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12616_ _12609_/X _12611_/X _12613_/X _12615_/X _12616_/C1 vssd1 vssd1 vccd1 vccd1
+ _12616_/X sky130_fd_sc_hd__o221a_1
X_15404_ _15589_/CLK _15404_/D vssd1 vssd1 vccd1 vccd1 _15404_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_169_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13596_ _15630_/CLK _13596_/D vssd1 vssd1 vccd1 vccd1 _13596_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_185_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15335_ _15335_/CLK _15335_/D vssd1 vssd1 vccd1 vccd1 _15335_/Q sky130_fd_sc_hd__dfxtp_2
X_12547_ _12540_/X _12542_/X _12544_/X _12546_/X _12616_/C1 vssd1 vssd1 vccd1 vccd1
+ _12547_/X sky130_fd_sc_hd__o221a_1
XFILLER_184_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15266_ _15298_/CLK _15266_/D vssd1 vssd1 vccd1 vccd1 _15266_/Q sky130_fd_sc_hd__dfxtp_1
X_12478_ _12471_/X _12473_/X _12475_/X _12477_/X _12501_/C1 vssd1 vssd1 vccd1 vccd1
+ _12478_/X sky130_fd_sc_hd__o221a_1
XANTENNA_3 _08659_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14217_ _14485_/CLK _14217_/D vssd1 vssd1 vccd1 vccd1 _14217_/Q sky130_fd_sc_hd__dfxtp_1
X_11429_ _11431_/A _11431_/B vssd1 vssd1 vccd1 vccd1 _11432_/A sky130_fd_sc_hd__nor2_1
XFILLER_6_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_963 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15197_ _15286_/CLK _15197_/D vssd1 vssd1 vccd1 vccd1 _15197_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14148_ _14225_/CLK _14148_/D vssd1 vssd1 vccd1 vccd1 _14148_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_140_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06970_ _14509_/Q _06707_/Y _06708_/Y _13499_/Q vssd1 vssd1 vccd1 vccd1 _06974_/B
+ sky130_fd_sc_hd__a2bb2o_1
X_14079_ _15233_/CLK _14079_/D vssd1 vssd1 vccd1 vccd1 _14079_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_79_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08640_ _13460_/Q _08684_/A2 _08691_/A2 _13595_/Q vssd1 vssd1 vccd1 vccd1 _08640_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_55_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08571_ _13606_/Q _08749_/A2 _08750_/B1 _13638_/Q vssd1 vssd1 vccd1 vccd1 _08571_/X
+ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_46_clk clkbuf_5_9_0_clk/X vssd1 vssd1 vccd1 vccd1 _15306_/CLK sky130_fd_sc_hd__clkbuf_16
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07522_ _14752_/Q _13431_/Q _07529_/S vssd1 vssd1 vccd1 vccd1 _13431_/D sky130_fd_sc_hd__mux2_1
XFILLER_35_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07453_ _13338_/A0 _13402_/Q _07501_/S vssd1 vssd1 vccd1 vccd1 _13402_/D sky130_fd_sc_hd__mux2_1
XFILLER_179_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07384_ _14736_/Q _07383_/X _07500_/S vssd1 vssd1 vccd1 vccd1 _07384_/X sky130_fd_sc_hd__mux2_8
X_09123_ _09449_/A1 _09121_/X _09122_/X _09449_/B2 _06676_/A vssd1 vssd1 vccd1 vccd1
+ _09123_/X sky130_fd_sc_hd__a221o_1
XFILLER_124_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09054_ _06676_/A _09043_/X _09052_/X _09053_/X vssd1 vssd1 vccd1 vccd1 _09054_/X
+ sky130_fd_sc_hd__o22a_2
XFILLER_68_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08005_ _14760_/Q _08022_/B _08004_/Y vssd1 vssd1 vccd1 vccd1 _13567_/D sky130_fd_sc_hd__o21a_1
XFILLER_163_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_218 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09956_ _11876_/A1 _14316_/Q _09958_/S vssd1 vssd1 vccd1 vccd1 _14316_/D sky130_fd_sc_hd__mux2_1
XFILLER_44_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08907_ _15274_/Q _15242_/Q _15210_/Q _15141_/Q _09469_/S _09546_/S1 vssd1 vssd1
+ vccd1 vccd1 _08907_/X sky130_fd_sc_hd__mux4_1
XFILLER_98_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09887_ _11873_/A1 _14249_/Q _09897_/S vssd1 vssd1 vccd1 vccd1 _14249_/D sky130_fd_sc_hd__mux2_1
XTAP_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08838_ _13861_/Q _13337_/A0 _08851_/S vssd1 vssd1 vccd1 vccd1 _13861_/D sky130_fd_sc_hd__mux2_1
XTAP_3415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08769_ _14612_/Q _08769_/B vssd1 vssd1 vccd1 vccd1 _08769_/X sky130_fd_sc_hd__and2_1
XTAP_2725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_37_clk clkbuf_5_12_0_clk/X vssd1 vssd1 vccd1 vccd1 _14863_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_2736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10800_ _14832_/Q _07337_/A _10871_/S vssd1 vssd1 vccd1 vccd1 _14832_/D sky130_fd_sc_hd__mux2_1
XTAP_2747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11780_ _13807_/Q _10891_/X _12904_/S vssd1 vssd1 vccd1 vccd1 _11781_/A sky130_fd_sc_hd__o21a_1
XTAP_2769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10731_ _15584_/Q _10731_/B vssd1 vssd1 vccd1 vccd1 _10731_/X sky130_fd_sc_hd__and2_1
XFILLER_80_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13450_ _15399_/CLK _13450_/D vssd1 vssd1 vccd1 vccd1 _13450_/Q sky130_fd_sc_hd__dfxtp_2
X_10662_ _15570_/Q _10706_/B _10722_/B1 _14947_/Q vssd1 vssd1 vccd1 vccd1 _10662_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_139_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12401_ _13961_/Q _13703_/Q _12407_/S vssd1 vssd1 vccd1 vccd1 _12402_/B sky130_fd_sc_hd__mux2_1
XFILLER_167_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13381_ _14484_/Q vssd1 vssd1 vccd1 vccd1 _14484_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_167_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10593_ _15556_/Q _10731_/B _10733_/A2 _14965_/Q vssd1 vssd1 vccd1 vccd1 _10593_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_182_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15120_ _15233_/CLK _15120_/D vssd1 vssd1 vccd1 vccd1 _15120_/Q sky130_fd_sc_hd__dfxtp_1
X_12332_ _13958_/Q _13700_/Q _12541_/S vssd1 vssd1 vccd1 vccd1 _12333_/B sky130_fd_sc_hd__mux2_1
XFILLER_5_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15051_ _15054_/CLK _15051_/D vssd1 vssd1 vccd1 vccd1 _15051_/Q sky130_fd_sc_hd__dfxtp_4
X_12263_ _13955_/Q _13697_/Q _12269_/S vssd1 vssd1 vccd1 vccd1 _12264_/B sky130_fd_sc_hd__mux2_1
X_14002_ _15324_/CLK _14002_/D vssd1 vssd1 vccd1 vccd1 _14002_/Q sky130_fd_sc_hd__dfxtp_1
X_11214_ _10382_/B _15003_/Q _11232_/S vssd1 vssd1 vccd1 vccd1 _15003_/D sky130_fd_sc_hd__mux2_1
X_12194_ _13952_/Q _13694_/Q _12499_/S vssd1 vssd1 vccd1 vccd1 _12195_/B sky130_fd_sc_hd__mux2_1
XFILLER_122_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput40 _07176_/X vssd1 vssd1 vccd1 vccd1 ext_address[14] sky130_fd_sc_hd__clkbuf_2
Xoutput51 _07187_/X vssd1 vssd1 vccd1 vccd1 ext_address[25] sky130_fd_sc_hd__clkbuf_2
Xoutput62 _07168_/X vssd1 vssd1 vccd1 vccd1 ext_address[6] sky130_fd_sc_hd__clkbuf_2
X_11145_ _11129_/A _11082_/A _11129_/Y vssd1 vssd1 vccd1 vccd1 _11193_/B sky130_fd_sc_hd__a21oi_1
Xoutput73 _07131_/X vssd1 vssd1 vccd1 vccd1 ext_write_data[15] sky130_fd_sc_hd__clkbuf_2
Xoutput84 _07151_/X vssd1 vssd1 vccd1 vccd1 ext_write_data[25] sky130_fd_sc_hd__clkbuf_2
XFILLER_95_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput95 _07114_/X vssd1 vssd1 vccd1 vccd1 ext_write_data[6] sky130_fd_sc_hd__clkbuf_2
X_11076_ _11259_/S _11024_/X _11075_/X vssd1 vssd1 vccd1 vccd1 _11076_/X sky130_fd_sc_hd__a21o_1
XFILLER_95_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10027_ _13348_/A0 _14385_/Q _10029_/S vssd1 vssd1 vccd1 vccd1 _14385_/D sky130_fd_sc_hd__mux2_1
X_14904_ _15530_/CLK _14904_/D vssd1 vssd1 vccd1 vccd1 _14904_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14835_ _15536_/CLK _14835_/D vssd1 vssd1 vccd1 vccd1 _14835_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_3960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_28_clk clkbuf_5_6_0_clk/X vssd1 vssd1 vccd1 vccd1 _15507_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_3971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11978_ _14458_/Q _14426_/Q _13847_/Q _14200_/Q _12154_/S _12253_/S1 vssd1 vssd1
+ vccd1 vccd1 _11978_/X sky130_fd_sc_hd__mux4_1
XFILLER_63_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14766_ _14861_/CLK _14766_/D vssd1 vssd1 vccd1 vccd1 _14766_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_91_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10929_ _11536_/C _10929_/B vssd1 vssd1 vccd1 vccd1 _10929_/Y sky130_fd_sc_hd__nand2_1
X_13717_ _14997_/CLK _13717_/D vssd1 vssd1 vccd1 vccd1 _13717_/Q sky130_fd_sc_hd__dfxtp_1
X_14697_ _15452_/CLK _14697_/D vssd1 vssd1 vccd1 vccd1 _14697_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13648_ _15372_/CLK _13648_/D vssd1 vssd1 vccd1 vccd1 _13648_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13579_ _14493_/CLK _13579_/D vssd1 vssd1 vccd1 vccd1 _13579_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_157_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_390 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15318_ _15661_/CLK _15318_/D vssd1 vssd1 vccd1 vccd1 _15318_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_172_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15249_ _15281_/CLK _15249_/D vssd1 vssd1 vccd1 vccd1 _15249_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09810_ _14176_/Q _13332_/A0 _09823_/S vssd1 vssd1 vccd1 vccd1 _14176_/D sky130_fd_sc_hd__mux2_1
Xfanout307 _07456_/X vssd1 vssd1 vccd1 vccd1 _13092_/B2 sky130_fd_sc_hd__buf_6
XFILLER_87_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout318 _07436_/X vssd1 vssd1 vccd1 vccd1 _13082_/B2 sky130_fd_sc_hd__buf_8
Xfanout329 _13328_/A0 vssd1 vssd1 vccd1 vccd1 _11861_/A1 sky130_fd_sc_hd__buf_6
XFILLER_115_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09741_ _14109_/Q _13329_/A0 _09757_/S vssd1 vssd1 vccd1 vccd1 _14109_/D sky130_fd_sc_hd__mux2_1
XFILLER_100_115 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06953_ _14486_/Q _06756_/Y _06947_/X _06963_/A _06952_/X vssd1 vssd1 vccd1 vccd1
+ _06953_/X sky130_fd_sc_hd__a2111o_1
XFILLER_95_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_243 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09672_ _14043_/Q _13327_/A0 _09690_/S vssd1 vssd1 vccd1 vccd1 _14043_/D sky130_fd_sc_hd__mux2_1
X_06884_ _15397_/Q _06694_/Y _15396_/Q _06696_/Y vssd1 vssd1 vccd1 vccd1 _06884_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_94_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08623_ _13559_/Q _08685_/A2 _08691_/B1 _13495_/Q vssd1 vssd1 vccd1 vccd1 _08623_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_36_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_19_clk clkbuf_5_3_0_clk/X vssd1 vssd1 vccd1 vccd1 _15332_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_1309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08554_ _13473_/Q _08746_/A2 _08750_/B1 _13640_/Q vssd1 vssd1 vccd1 vccd1 _08554_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_42_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07505_ _14718_/Q _08037_/C _08025_/C _14717_/Q vssd1 vssd1 vccd1 vccd1 _07505_/X
+ sky130_fd_sc_hd__or4b_4
XFILLER_35_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08485_ _08453_/A _08477_/X _08484_/X vssd1 vssd1 vccd1 vccd1 _08485_/X sky130_fd_sc_hd__a21o_1
XFILLER_22_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07436_ _14749_/Q _07435_/X _07480_/S vssd1 vssd1 vccd1 vccd1 _07436_/X sky130_fd_sc_hd__mux2_8
XFILLER_51_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07367_ _14712_/Q _08817_/B vssd1 vssd1 vccd1 vccd1 _09662_/B sky130_fd_sc_hd__nand2_8
XFILLER_109_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09106_ _13885_/Q _09445_/A2 _09522_/B1 _14400_/Q _09437_/A1 vssd1 vssd1 vccd1 vccd1
+ _09106_/X sky130_fd_sc_hd__a221o_1
XFILLER_108_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07298_ _15317_/Q _15473_/Q _07340_/S vssd1 vssd1 vccd1 vccd1 _07298_/X sky130_fd_sc_hd__mux2_8
XFILLER_108_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09037_ _14363_/Q _15179_/Q _13818_/Q _14557_/Q _09225_/S0 _09225_/S1 vssd1 vssd1
+ vccd1 vccd1 _09038_/B sky130_fd_sc_hd__mux4_1
XFILLER_163_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09939_ _12967_/A1 _14299_/Q _09958_/S vssd1 vssd1 vccd1 vccd1 _14299_/D sky130_fd_sc_hd__mux2_1
XFILLER_58_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_4_13_0_clk clkbuf_3_6_0_clk/X vssd1 vssd1 vccd1 vccd1 clkbuf_5_27_0_clk/A
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_58_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12950_ _15463_/Q _13139_/S _13116_/C _12949_/X vssd1 vssd1 vccd1 vccd1 _15463_/D
+ sky130_fd_sc_hd__a22o_1
XTAP_3201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_75 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11901_ _14067_/Q _14035_/Q _12269_/S vssd1 vssd1 vccd1 vccd1 _11901_/X sky130_fd_sc_hd__mux2_1
XTAP_3234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12881_ _15409_/Q _15594_/Q _12885_/S vssd1 vssd1 vccd1 vccd1 _15409_/D sky130_fd_sc_hd__mux2_1
XTAP_3245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11832_ _15254_/Q _13332_/A0 _11849_/S vssd1 vssd1 vccd1 vccd1 _15254_/D sky130_fd_sc_hd__mux2_1
XFILLER_93_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14620_ _15623_/CLK _14620_/D vssd1 vssd1 vccd1 vccd1 _14620_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14551_ _14606_/CLK _14551_/D vssd1 vssd1 vccd1 vccd1 _14551_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11763_ _11838_/A1 _15191_/Q _11775_/S vssd1 vssd1 vccd1 vccd1 _15191_/D sky130_fd_sc_hd__mux2_1
XTAP_1854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10714_ _15070_/Q _10714_/A2 _10711_/X _10713_/X vssd1 vssd1 vccd1 vccd1 _10714_/X
+ sky130_fd_sc_hd__o22a_4
X_13502_ _14511_/CLK _13502_/D vssd1 vssd1 vccd1 vccd1 _13502_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_1887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14482_ _14482_/CLK _14482_/D vssd1 vssd1 vccd1 vccd1 _14482_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11694_ _13336_/A0 _15125_/Q _11708_/S vssd1 vssd1 vccd1 vccd1 _15125_/D sky130_fd_sc_hd__mux2_1
X_13433_ _15389_/CLK _13433_/D vssd1 vssd1 vccd1 vccd1 _13433_/Q sky130_fd_sc_hd__dfxtp_1
X_10645_ _14747_/Q _10644_/X _10650_/S vssd1 vssd1 vccd1 vccd1 _14747_/D sky130_fd_sc_hd__mux2_1
XFILLER_167_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13364_ _14467_/Q vssd1 vssd1 vccd1 vccd1 _14467_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_158_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10576_ _14927_/Q _14928_/Q _14929_/Q vssd1 vssd1 vccd1 vccd1 _10576_/X sky130_fd_sc_hd__and3b_2
X_12315_ _14085_/Q _14053_/Q _12614_/S vssd1 vssd1 vccd1 vccd1 _12315_/X sky130_fd_sc_hd__mux2_1
X_15103_ _15670_/CLK _15103_/D vssd1 vssd1 vccd1 vccd1 _15103_/Q sky130_fd_sc_hd__dfxtp_1
X_13295_ _12689_/Y _15627_/Q _13300_/S vssd1 vssd1 vccd1 vccd1 _15627_/D sky130_fd_sc_hd__mux2_1
XFILLER_154_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15034_ _15042_/CLK _15034_/D vssd1 vssd1 vccd1 vccd1 _15034_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_142_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12246_ _14082_/Q _14050_/Q _12246_/S vssd1 vssd1 vccd1 vccd1 _12246_/X sky130_fd_sc_hd__mux2_1
XFILLER_177_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12177_ _14079_/Q _14047_/Q _12246_/S vssd1 vssd1 vccd1 vccd1 _12177_/X sky130_fd_sc_hd__mux2_1
XFILLER_122_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_327 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11128_ _14969_/Q _11202_/A _11127_/X vssd1 vssd1 vccd1 vccd1 _14969_/D sky130_fd_sc_hd__o21ba_1
XFILLER_1_581 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11059_ _10972_/B _10978_/X _11330_/A vssd1 vssd1 vccd1 vccd1 _11059_/X sky130_fd_sc_hd__mux2_1
XFILLER_49_574 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14818_ _15636_/CLK _14818_/D vssd1 vssd1 vccd1 vccd1 _14818_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_184_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14749_ _15608_/CLK _14749_/D vssd1 vssd1 vccd1 vccd1 _14749_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_33_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08270_ _10507_/A1 _13771_/Q _15401_/Q _10515_/B2 vssd1 vssd1 vccd1 vccd1 _08270_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_149_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07221_ _07221_/A vssd1 vssd1 vccd1 vccd1 _07221_/Y sky130_fd_sc_hd__inv_2
XFILLER_146_800 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07152_ _14856_/Q _14848_/Q _14840_/Q _14832_/Q _07146_/S _07104_/C vssd1 vssd1 vccd1
+ vccd1 _07153_/B sky130_fd_sc_hd__mux4_1
XFILLER_118_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_1044 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07083_ _07082_/X _14760_/Q _07098_/S vssd1 vssd1 vccd1 vccd1 _13606_/D sky130_fd_sc_hd__mux2_1
XFILLER_106_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_8_clk clkbuf_5_3_0_clk/X vssd1 vssd1 vccd1 vccd1 _15133_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_133_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout104 _12622_/X vssd1 vssd1 vccd1 vccd1 _12759_/B sky130_fd_sc_hd__buf_12
Xfanout115 _12946_/Y vssd1 vssd1 vccd1 vccd1 _13025_/B1 sky130_fd_sc_hd__clkbuf_16
XFILLER_102_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout126 _13140_/S vssd1 vssd1 vccd1 vccd1 _13120_/S sky130_fd_sc_hd__clkbuf_16
XFILLER_102_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout137 fanout138/X vssd1 vssd1 vccd1 vccd1 _10765_/S sky130_fd_sc_hd__buf_12
Xfanout148 _06781_/X vssd1 vssd1 vccd1 vccd1 _12320_/A sky130_fd_sc_hd__buf_12
X_07985_ _13561_/Q _13560_/Q _07984_/D _13562_/Q vssd1 vssd1 vccd1 vccd1 _07985_/Y
+ sky130_fd_sc_hd__a31oi_1
XFILLER_101_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout159 _06781_/X vssd1 vssd1 vccd1 vccd1 _08573_/S sky130_fd_sc_hd__buf_12
XFILLER_101_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09724_ _13346_/A0 _14094_/Q _09728_/S vssd1 vssd1 vccd1 vccd1 _14094_/D sky130_fd_sc_hd__mux2_1
X_06936_ _14501_/Q _06936_/B vssd1 vssd1 vccd1 vccd1 _06936_/Y sky130_fd_sc_hd__nand2_1
XFILLER_170_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_1034 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09655_ _14028_/Q _13344_/A0 _09660_/S vssd1 vssd1 vccd1 vccd1 _14028_/D sky130_fd_sc_hd__mux2_1
XFILLER_67_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06867_ _06697_/Y _13504_/Q _06700_/Y _13503_/Q vssd1 vssd1 vccd1 vccd1 _06882_/B
+ sky130_fd_sc_hd__a22o_1
X_08606_ _13785_/Q _08626_/S _08605_/X vssd1 vssd1 vccd1 vccd1 _13785_/D sky130_fd_sc_hd__o21a_1
XFILLER_15_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09586_ _13962_/Q _13342_/A0 _09594_/S vssd1 vssd1 vccd1 vccd1 _13962_/D sky130_fd_sc_hd__mux2_1
XFILLER_83_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_3_2_0_clk clkbuf_3_3_0_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_5_0_clk/A sky130_fd_sc_hd__clkbuf_8
XTAP_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06798_ _14589_/Q _14587_/Q _06798_/C vssd1 vssd1 vccd1 vccd1 _08477_/C sky130_fd_sc_hd__and3_4
XTAP_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08537_ _08537_/A _08538_/B vssd1 vssd1 vccd1 vccd1 _08537_/Y sky130_fd_sc_hd__nor2_4
XFILLER_179_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08468_ _13763_/Q _08467_/X _12900_/S vssd1 vssd1 vccd1 vccd1 _13763_/D sky130_fd_sc_hd__mux2_1
XFILLER_51_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07419_ _13660_/Q _07499_/A2 _07499_/B1 _14688_/Q _07418_/X vssd1 vssd1 vccd1 vccd1
+ _07419_/X sky130_fd_sc_hd__a221o_1
X_08399_ _13733_/Q _13140_/S _08394_/X hold5/X vssd1 vssd1 vccd1 vccd1 _13733_/D sky130_fd_sc_hd__a22o_1
XFILLER_149_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10430_ _11639_/A _10430_/B vssd1 vssd1 vccd1 vccd1 _10537_/A sky130_fd_sc_hd__or2_1
XFILLER_183_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10361_ _08240_/A _13791_/Q _13759_/Q _08237_/A _10360_/X vssd1 vssd1 vccd1 vccd1
+ _11496_/B sky130_fd_sc_hd__a221oi_4
XFILLER_136_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12100_ _12500_/B1 _12097_/X _12501_/C1 vssd1 vssd1 vccd1 vccd1 _12100_/X sky130_fd_sc_hd__o21a_1
X_13080_ _12987_/X _13104_/A2 _13104_/B1 _13080_/B2 vssd1 vssd1 vccd1 vccd1 _13080_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_163_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10292_ _14677_/Q _14862_/Q _10615_/S vssd1 vssd1 vccd1 vccd1 _14677_/D sky130_fd_sc_hd__mux2_1
XFILLER_152_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12031_ _06670_/A _12028_/X _06671_/A vssd1 vssd1 vccd1 vccd1 _12031_/X sky130_fd_sc_hd__o21a_1
XFILLER_104_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_722 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13982_ _15285_/CLK _13982_/D vssd1 vssd1 vccd1 vccd1 _13982_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12933_ _15461_/Q _15647_/Q _12933_/S vssd1 vssd1 vccd1 vccd1 _15461_/D sky130_fd_sc_hd__mux2_1
XTAP_3031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15652_ _15652_/CLK _15652_/D vssd1 vssd1 vccd1 vccd1 _15652_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12864_ _14758_/Q _15392_/Q _12866_/S vssd1 vssd1 vccd1 vccd1 _15392_/D sky130_fd_sc_hd__mux2_1
XTAP_3086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14603_ _15622_/CLK _14603_/D vssd1 vssd1 vccd1 vccd1 _14603_/Q sky130_fd_sc_hd__dfxtp_1
X_11815_ _15238_/Q _11881_/A1 _11817_/S vssd1 vssd1 vccd1 vccd1 _15238_/D sky130_fd_sc_hd__mux2_1
XTAP_2374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12795_ _15361_/Q _12765_/B _12794_/X _12809_/C1 vssd1 vssd1 vccd1 vccd1 _15361_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_15_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15583_ _15613_/CLK _15583_/D vssd1 vssd1 vccd1 vccd1 _15583_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14534_ _15212_/CLK _14534_/D vssd1 vssd1 vccd1 vccd1 _14534_/Q sky130_fd_sc_hd__dfxtp_1
X_11746_ _11854_/A1 _15174_/Q _11775_/S vssd1 vssd1 vccd1 vccd1 _15174_/D sky130_fd_sc_hd__mux2_1
XFILLER_186_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11677_ _13319_/A0 _15108_/Q _11703_/S vssd1 vssd1 vccd1 vccd1 _15108_/D sky130_fd_sc_hd__mux2_1
X_14465_ _15663_/CLK _14465_/D vssd1 vssd1 vccd1 vccd1 _14465_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_800 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10628_ _14972_/Q _10718_/A2 _10722_/B1 _14940_/Q _10627_/X vssd1 vssd1 vccd1 vccd1
+ _10628_/X sky130_fd_sc_hd__a221o_1
X_13416_ _15429_/CLK _13416_/D vssd1 vssd1 vccd1 vccd1 _13416_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_139_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14396_ _15178_/CLK _14396_/D vssd1 vssd1 vccd1 vccd1 _14396_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_183_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13347_ _13347_/A0 _15677_/Q _13350_/S vssd1 vssd1 vccd1 vccd1 _15677_/D sky130_fd_sc_hd__mux2_1
XFILLER_115_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10559_ _10420_/A _11239_/B _11240_/A vssd1 vssd1 vccd1 vccd1 _10559_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_128_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_493 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13278_ _15362_/Q _15609_/Q _13309_/A vssd1 vssd1 vccd1 vccd1 _15609_/D sky130_fd_sc_hd__mux2_1
X_15017_ _15017_/CLK _15017_/D vssd1 vssd1 vccd1 vccd1 _15017_/Q sky130_fd_sc_hd__dfxtp_1
X_12229_ _15320_/Q _13105_/A2 _12228_/X vssd1 vssd1 vccd1 vccd1 _15320_/D sky130_fd_sc_hd__a21o_1
XFILLER_97_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07770_ _07768_/Y _07776_/C _07676_/A vssd1 vssd1 vccd1 vccd1 _07770_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_65_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06721_ _15384_/Q vssd1 vssd1 vccd1 vccd1 _06919_/A sky130_fd_sc_hd__inv_2
XFILLER_49_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09440_ _09449_/A1 _09438_/X _09439_/X _09449_/B2 _09437_/X vssd1 vssd1 vccd1 vccd1
+ _09440_/X sky130_fd_sc_hd__a221o_1
XFILLER_65_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09371_ _09532_/A _09371_/B vssd1 vssd1 vccd1 vccd1 _09371_/X sky130_fd_sc_hd__or2_1
XFILLER_17_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08322_ _13721_/Q _11346_/A2 _11351_/C1 _08321_/X vssd1 vssd1 vccd1 vccd1 _13721_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_33_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_271 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08253_ _10507_/A1 _13773_/Q _15431_/Q _10515_/B2 vssd1 vssd1 vccd1 vccd1 _08253_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_138_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07204_ _07204_/A vssd1 vssd1 vccd1 vccd1 _07204_/Y sky130_fd_sc_hd__inv_2
XFILLER_165_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08184_ _13679_/Q _10730_/S _08155_/X _08183_/X vssd1 vssd1 vccd1 vccd1 _13679_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_174_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07135_ _14831_/Q _07104_/X _07134_/X _07131_/A vssd1 vssd1 vccd1 vccd1 _07135_/X
+ sky130_fd_sc_hd__a22o_4
XFILLER_118_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_460 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07066_ _14634_/Q _14666_/Q _07096_/S vssd1 vssd1 vccd1 vccd1 _07066_/X sky130_fd_sc_hd__mux2_1
XFILLER_134_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_250_clk clkbuf_5_1_0_clk/X vssd1 vssd1 vccd1 vccd1 _15649_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_75_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07968_ _07970_/B _07967_/X _07971_/A vssd1 vssd1 vccd1 vccd1 _07968_/X sky130_fd_sc_hd__a21bo_1
X_06919_ _06919_/A _13461_/Q vssd1 vssd1 vccd1 vccd1 _06921_/A sky130_fd_sc_hd__nor2_1
XFILLER_28_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09707_ _13072_/B2 _14077_/Q _09723_/S vssd1 vssd1 vccd1 vccd1 _14077_/D sky130_fd_sc_hd__mux2_1
XFILLER_56_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07899_ _14764_/Q _07903_/A _07898_/Y _08016_/C1 vssd1 vssd1 vccd1 vccd1 _13539_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_28_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09638_ _14011_/Q _13327_/A0 _09660_/S vssd1 vssd1 vccd1 vccd1 _14011_/D sky130_fd_sc_hd__mux2_1
XFILLER_71_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09569_ _13945_/Q _13325_/A0 _09594_/S vssd1 vssd1 vccd1 vccd1 _13945_/D sky130_fd_sc_hd__mux2_1
XFILLER_130_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11600_ _11600_/A _11600_/B vssd1 vssd1 vccd1 vccd1 _11602_/B sky130_fd_sc_hd__xnor2_1
XFILLER_130_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12580_ _14386_/Q _15202_/Q _13841_/Q _14580_/Q _12591_/S _12590_/A vssd1 vssd1 vccd1
+ vccd1 _12580_/X sky130_fd_sc_hd__mux4_1
XFILLER_142_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11531_ _11531_/A _11531_/B vssd1 vssd1 vccd1 vccd1 _11534_/A sky130_fd_sc_hd__nand2_1
XFILLER_157_928 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_736 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14250_ _15295_/CLK _14250_/D vssd1 vssd1 vccd1 vccd1 _14250_/Q sky130_fd_sc_hd__dfxtp_1
X_11462_ _11442_/Y _11460_/C _11461_/X _11450_/A vssd1 vssd1 vccd1 vccd1 _11464_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_184_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13201_ _13219_/S _13199_/X _13200_/Y _13198_/X vssd1 vssd1 vccd1 vccd1 _15567_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_104_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10413_ _10395_/B _10411_/X _10412_/X _10558_/A vssd1 vssd1 vccd1 vccd1 _10413_/X
+ sky130_fd_sc_hd__a31o_2
XFILLER_183_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14181_ _14439_/CLK _14181_/D vssd1 vssd1 vccd1 vccd1 _14181_/Q sky130_fd_sc_hd__dfxtp_1
X_11393_ _11423_/A _11423_/B _11401_/A _11384_/A vssd1 vssd1 vccd1 vccd1 _11394_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_152_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13132_ _14612_/Q _14611_/Q _13130_/X _13131_/Y vssd1 vssd1 vccd1 vccd1 _13134_/B
+ sky130_fd_sc_hd__a2bb2o_1
X_10344_ _14922_/Q _14729_/Q _10344_/S vssd1 vssd1 vccd1 vccd1 _14729_/D sky130_fd_sc_hd__mux2_1
XFILLER_174_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13063_ _15499_/Q _13119_/S _13042_/A _13062_/X vssd1 vssd1 vccd1 vccd1 _15499_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_112_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10275_ _14660_/Q _14813_/Q _10710_/S vssd1 vssd1 vccd1 vccd1 _14660_/D sky130_fd_sc_hd__mux2_1
XFILLER_2_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12014_ _14008_/Q _13976_/Q _12407_/S vssd1 vssd1 vccd1 vccd1 _12015_/B sky130_fd_sc_hd__mux2_1
XFILLER_2_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_241_clk clkbuf_5_5_0_clk/X vssd1 vssd1 vccd1 vccd1 _15281_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_78_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout490 _07104_/C vssd1 vssd1 vccd1 vccd1 _08151_/S sky130_fd_sc_hd__clkbuf_16
X_13965_ _14405_/CLK _13965_/D vssd1 vssd1 vccd1 vccd1 _13965_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12916_ _15444_/Q _15630_/Q _12928_/S vssd1 vssd1 vccd1 vccd1 _15444_/D sky130_fd_sc_hd__mux2_1
XFILLER_46_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13896_ _15680_/CLK _13896_/D vssd1 vssd1 vccd1 vccd1 _13896_/Q sky130_fd_sc_hd__dfxtp_1
X_15635_ _15635_/CLK _15635_/D vssd1 vssd1 vccd1 vccd1 _15635_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12847_ _14741_/Q _15375_/Q _12871_/S vssd1 vssd1 vccd1 vccd1 _15375_/D sky130_fd_sc_hd__mux2_1
XFILLER_61_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15566_ _15580_/CLK _15566_/D vssd1 vssd1 vccd1 vccd1 _15566_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12778_ _12828_/A _12778_/B vssd1 vssd1 vccd1 vccd1 _12778_/X sky130_fd_sc_hd__or2_1
XFILLER_15_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14517_ _14517_/CLK _14517_/D vssd1 vssd1 vccd1 vccd1 _14517_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11729_ _15158_/Q _11870_/A1 _11742_/S vssd1 vssd1 vccd1 vccd1 _15158_/D sky130_fd_sc_hd__mux2_1
X_15497_ _15497_/CLK _15497_/D vssd1 vssd1 vccd1 vccd1 _15497_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_174_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14448_ _15556_/CLK _14448_/D vssd1 vssd1 vccd1 vccd1 _14448_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14379_ _15336_/CLK _14379_/D vssd1 vssd1 vccd1 vccd1 _14379_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_142_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08940_ _14005_/Q _13973_/Q _09484_/S vssd1 vssd1 vccd1 vccd1 _08940_/X sky130_fd_sc_hd__mux2_1
XFILLER_124_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_496 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08871_ _13892_/Q _11761_/A0 _08885_/S vssd1 vssd1 vccd1 vccd1 _13892_/D sky130_fd_sc_hd__mux2_1
X_07822_ _13518_/Q _07825_/D _13519_/Q vssd1 vssd1 vccd1 vccd1 _07822_/Y sky130_fd_sc_hd__a21oi_1
Xclkbuf_leaf_232_clk clkbuf_5_4_0_clk/X vssd1 vssd1 vccd1 vccd1 _15656_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_57_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_127 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07753_ _13502_/Q _13501_/Q _07757_/D vssd1 vssd1 vccd1 vccd1 _07756_/B sky130_fd_sc_hd__and3_1
XFILLER_38_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06704_ _15392_/Q vssd1 vssd1 vccd1 vccd1 _06704_/Y sky130_fd_sc_hd__inv_2
X_07684_ _07682_/Y _07686_/B _07676_/A vssd1 vssd1 vccd1 vccd1 _07684_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_25_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09423_ _14092_/Q _09445_/A2 _08508_/Y _14060_/Q _09221_/A vssd1 vssd1 vccd1 vccd1
+ _09423_/X sky130_fd_sc_hd__a221o_1
XFILLER_53_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09354_ _14444_/Q _08540_/B _08520_/B _09353_/X vssd1 vssd1 vccd1 vccd1 _09354_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_178_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08305_ _11044_/B _11045_/A vssd1 vssd1 vccd1 vccd1 _08305_/X sky130_fd_sc_hd__or2_1
XFILLER_127_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09285_ _15292_/Q _15260_/Q _15228_/Q _15159_/Q _09484_/S _08519_/A vssd1 vssd1 vccd1
+ vccd1 _09285_/X sky130_fd_sc_hd__mux4_1
X_08236_ _07337_/A _10457_/A2 _08234_/X vssd1 vssd1 vccd1 vccd1 _08236_/X sky130_fd_sc_hd__a21o_4
XFILLER_165_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08167_ _08185_/A _08167_/B vssd1 vssd1 vccd1 vccd1 _08167_/X sky130_fd_sc_hd__and2_1
XFILLER_134_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_696 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07118_ _14839_/Q _14831_/Q _08094_/S vssd1 vssd1 vccd1 vccd1 _07119_/B sky130_fd_sc_hd__mux2_1
XFILLER_133_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08098_ input9/X input18/X _08133_/S vssd1 vssd1 vccd1 vccd1 _08157_/B sky130_fd_sc_hd__mux2_1
XFILLER_118_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07049_ _07048_/X _13595_/Q _12728_/S vssd1 vssd1 vccd1 vccd1 _07049_/X sky130_fd_sc_hd__mux2_1
XFILLER_134_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10060_ _14417_/Q _13346_/A0 _10064_/S vssd1 vssd1 vccd1 vccd1 _14417_/D sky130_fd_sc_hd__mux2_1
XFILLER_102_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_850 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_679 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_223_clk clkbuf_5_7_0_clk/X vssd1 vssd1 vccd1 vccd1 _15536_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_88_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_108 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10962_ _11023_/A _13242_/B vssd1 vssd1 vccd1 vccd1 _10963_/B sky130_fd_sc_hd__nand2_1
XFILLER_29_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13750_ _14868_/CLK _13750_/D vssd1 vssd1 vccd1 vccd1 _13750_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_43_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12701_ _15349_/Q _15348_/Q _12701_/C vssd1 vssd1 vccd1 vccd1 _12710_/B sky130_fd_sc_hd__and3_1
XFILLER_44_856 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13681_ _15665_/CLK _13681_/D vssd1 vssd1 vccd1 vccd1 _13681_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10893_ _14924_/Q _12904_/S _10892_/X vssd1 vssd1 vccd1 vccd1 _14924_/D sky130_fd_sc_hd__o21a_1
XFILLER_70_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15420_ _15638_/CLK _15420_/D vssd1 vssd1 vccd1 vccd1 _15420_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_70_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12632_ _13416_/Q _12631_/X _12640_/S vssd1 vssd1 vccd1 vccd1 _12633_/B sky130_fd_sc_hd__mux2_1
X_15351_ _15630_/CLK _15351_/D vssd1 vssd1 vccd1 vccd1 _15351_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_15_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12563_ _12563_/A _12563_/B vssd1 vssd1 vccd1 vccd1 _12563_/X sky130_fd_sc_hd__and2_1
XFILLER_184_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11514_ _10483_/A _10483_/B _11512_/B vssd1 vssd1 vccd1 vccd1 _11515_/B sky130_fd_sc_hd__o21bai_1
X_14302_ _14468_/CLK _14302_/D vssd1 vssd1 vccd1 vccd1 _14302_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15282_ _15674_/CLK _15282_/D vssd1 vssd1 vccd1 vccd1 _15282_/Q sky130_fd_sc_hd__dfxtp_1
X_12494_ _12498_/A _12494_/B vssd1 vssd1 vccd1 vccd1 _12494_/X sky130_fd_sc_hd__and2_1
XFILLER_8_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11445_ _11443_/Y _11444_/X _15053_/Q _11474_/S vssd1 vssd1 vccd1 vccd1 _15053_/D
+ sky130_fd_sc_hd__a2bb2o_1
X_14233_ _15211_/CLK _14233_/D vssd1 vssd1 vccd1 vccd1 _14233_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_171_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14164_ _15650_/CLK _14164_/D vssd1 vssd1 vccd1 vccd1 _14164_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_153_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11376_ _11368_/A _11368_/B _11377_/B _11363_/X vssd1 vssd1 vccd1 vccd1 _11423_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_4_952 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13115_ _15525_/Q _13129_/A _13042_/A _13114_/X vssd1 vssd1 vccd1 vccd1 _15525_/D
+ sky130_fd_sc_hd__a22o_1
X_10327_ _14905_/Q _14712_/Q _10566_/B vssd1 vssd1 vccd1 vccd1 _14712_/D sky130_fd_sc_hd__mux2_1
XFILLER_152_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14095_ _15677_/CLK _14095_/D vssd1 vssd1 vccd1 vccd1 _14095_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_112_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_152_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13046_ _08910_/S _09662_/B _08852_/B _08508_/B _13045_/Y vssd1 vssd1 vccd1 vccd1
+ _13050_/A sky130_fd_sc_hd__o221a_1
XFILLER_105_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10258_ _14643_/Q _14796_/Q _10615_/S vssd1 vssd1 vccd1 vccd1 _14643_/D sky130_fd_sc_hd__mux2_1
XFILLER_39_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_214_clk clkbuf_5_18_0_clk/X vssd1 vssd1 vccd1 vccd1 _15335_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_94_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10189_ _13098_/B2 _14573_/Q _10197_/S vssd1 vssd1 vccd1 vccd1 _14573_/D sky130_fd_sc_hd__mux2_1
XFILLER_67_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14997_ _14997_/CLK _14997_/D vssd1 vssd1 vccd1 vccd1 _14997_/Q sky130_fd_sc_hd__dfxtp_1
X_13948_ _14530_/CLK _13948_/D vssd1 vssd1 vccd1 vccd1 _13948_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13879_ _15108_/CLK _13879_/D vssd1 vssd1 vccd1 vccd1 _13879_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15618_ _15618_/CLK _15618_/D vssd1 vssd1 vccd1 vccd1 _15618_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15549_ _15552_/CLK _15549_/D vssd1 vssd1 vccd1 vccd1 _15549_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_188_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09070_ _09391_/A _09070_/B vssd1 vssd1 vccd1 vccd1 _09070_/X sky130_fd_sc_hd__or2_1
XFILLER_163_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08021_ _13572_/Q _08021_/B vssd1 vssd1 vccd1 vccd1 _08021_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_129_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09972_ _12967_/A1 _14331_/Q _09991_/S vssd1 vssd1 vccd1 vccd1 _14331_/D sky130_fd_sc_hd__mux2_1
XFILLER_116_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08923_ _09546_/S1 _08519_/B _08922_/X _08501_/A vssd1 vssd1 vccd1 vccd1 _08923_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_97_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_205_clk clkbuf_5_16_0_clk/X vssd1 vssd1 vccd1 vccd1 _15178_/CLK sky130_fd_sc_hd__clkbuf_16
X_08854_ _13875_/Q _13319_/A0 _08880_/S vssd1 vssd1 vccd1 vccd1 _13875_/D sky130_fd_sc_hd__mux2_1
XFILLER_57_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07805_ _14739_/Q _07816_/A _07804_/Y _08084_/C1 vssd1 vssd1 vccd1 vccd1 _13514_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_3619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08785_ _11852_/A1 _13811_/Q _08811_/S vssd1 vssd1 vccd1 vccd1 _13811_/D sky130_fd_sc_hd__mux2_1
XFILLER_44_108 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07736_ _07736_/A _07736_/B vssd1 vssd1 vccd1 vccd1 _07736_/Y sky130_fd_sc_hd__nand2_1
XFILLER_66_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_940 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07667_ _14735_/Q _07777_/A _07666_/Y _08016_/C1 vssd1 vssd1 vccd1 vccd1 _13478_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_111_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09406_ _14542_/Q _14155_/Q _14187_/Q _14123_/Q _09407_/S _09406_/S1 vssd1 vssd1
+ vccd1 vccd1 _09406_/X sky130_fd_sc_hd__mux4_1
X_07598_ _14749_/Q _07607_/A _07597_/Y _07965_/C1 vssd1 vssd1 vccd1 vccd1 _13460_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_71_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09337_ _14024_/Q _13992_/Q _09342_/S vssd1 vssd1 vccd1 vccd1 _09337_/X sky130_fd_sc_hd__mux2_1
XFILLER_179_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09268_ _08510_/B _09264_/X _09267_/X _09263_/X vssd1 vssd1 vccd1 vccd1 _09281_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_138_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08219_ _13710_/Q _11881_/A1 _08221_/S vssd1 vssd1 vccd1 vccd1 _13710_/D sky130_fd_sc_hd__mux2_1
XFILLER_14_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09199_ _15288_/Q _15256_/Q _15224_/Q _15155_/Q _09441_/S _09448_/S1 vssd1 vssd1
+ vccd1 vccd1 _09199_/X sky130_fd_sc_hd__mux4_1
XFILLER_119_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11230_ _10470_/B _15018_/Q _11232_/S vssd1 vssd1 vccd1 vccd1 _15018_/D sky130_fd_sc_hd__mux2_1
XFILLER_135_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11161_ _11347_/A _11161_/B vssd1 vssd1 vccd1 vccd1 _11161_/Y sky130_fd_sc_hd__nor2_1
XFILLER_84_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10112_ _14498_/Q _14746_/Q _10124_/S vssd1 vssd1 vccd1 vccd1 _14498_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11092_ _14965_/Q _10984_/Y _11090_/Y _11091_/Y vssd1 vssd1 vccd1 vccd1 _14965_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_1_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10043_ _14400_/Q _13072_/B2 _10059_/S vssd1 vssd1 vccd1 vccd1 _14400_/D sky130_fd_sc_hd__mux2_1
X_14920_ _15676_/CLK _14920_/D vssd1 vssd1 vccd1 vccd1 _14920_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14851_ _14851_/CLK _14851_/D vssd1 vssd1 vccd1 vccd1 _14851_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13802_ _15587_/CLK _13802_/D vssd1 vssd1 vccd1 vccd1 _13802_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14782_ _15596_/CLK _14782_/D vssd1 vssd1 vccd1 vccd1 _14782_/Q sky130_fd_sc_hd__dfxtp_1
X_11994_ _12500_/A1 _11993_/X _12500_/B1 vssd1 vssd1 vccd1 vccd1 _11994_/X sky130_fd_sc_hd__a21o_1
XFILLER_21_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13733_ _15530_/CLK _13733_/D vssd1 vssd1 vccd1 vccd1 _13733_/Q sky130_fd_sc_hd__dfxtp_2
X_10945_ _14957_/Q _10944_/B _10944_/Y _11610_/A vssd1 vssd1 vccd1 vccd1 _14957_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_43_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13664_ _15606_/CLK _13664_/D vssd1 vssd1 vccd1 vccd1 _13664_/Q sky130_fd_sc_hd__dfxtp_1
X_10876_ _13730_/Q _14908_/Q _10877_/S vssd1 vssd1 vccd1 vccd1 _14908_/D sky130_fd_sc_hd__mux2_1
X_15403_ _15588_/CLK _15403_/D vssd1 vssd1 vccd1 vccd1 _15403_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12615_ _12615_/A1 _12614_/X _12615_/B1 vssd1 vssd1 vccd1 vccd1 _12615_/X sky130_fd_sc_hd__a21o_1
XPHY_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13595_ _15630_/CLK _13595_/D vssd1 vssd1 vccd1 vccd1 _13595_/Q sky130_fd_sc_hd__dfxtp_2
XPHY_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15334_ _15334_/CLK _15334_/D vssd1 vssd1 vccd1 vccd1 _15334_/Q sky130_fd_sc_hd__dfxtp_2
X_12546_ _12615_/A1 _12545_/X _12615_/B1 vssd1 vssd1 vccd1 vccd1 _12546_/X sky130_fd_sc_hd__a21o_1
XFILLER_184_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15265_ _15518_/CLK _15265_/D vssd1 vssd1 vccd1 vccd1 _15265_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_177_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12477_ _12477_/A1 _12476_/X _12500_/B1 vssd1 vssd1 vccd1 vccd1 _12477_/X sky130_fd_sc_hd__a21o_1
XFILLER_144_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_4 _08688_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14216_ _15669_/CLK _14216_/D vssd1 vssd1 vccd1 vccd1 _14216_/Q sky130_fd_sc_hd__dfxtp_1
X_11428_ _11436_/B _11428_/B vssd1 vssd1 vccd1 vccd1 _11431_/B sky130_fd_sc_hd__xor2_2
X_15196_ _15652_/CLK _15196_/D vssd1 vssd1 vccd1 vccd1 _15196_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14147_ _15212_/CLK _14147_/D vssd1 vssd1 vccd1 vccd1 _14147_/Q sky130_fd_sc_hd__dfxtp_1
X_11359_ _11359_/A _11359_/B vssd1 vssd1 vccd1 vccd1 _11360_/B sky130_fd_sc_hd__nor2_1
XFILLER_113_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14078_ _15253_/CLK _14078_/D vssd1 vssd1 vccd1 vccd1 _14078_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_140_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13029_ _10719_/X _14890_/Q _13029_/S vssd1 vssd1 vccd1 vccd1 _13029_/X sky130_fd_sc_hd__mux2_4
XFILLER_6_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_553 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08570_ _15394_/Q _08748_/A2 _08736_/A2 _13439_/Q vssd1 vssd1 vccd1 vccd1 _08570_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_82_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07521_ _14751_/Q _13430_/Q _07529_/S vssd1 vssd1 vccd1 vccd1 _13430_/D sky130_fd_sc_hd__mux2_1
XFILLER_63_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07452_ _14753_/Q _07451_/X _07480_/S vssd1 vssd1 vccd1 vccd1 _07452_/X sky130_fd_sc_hd__mux2_8
XFILLER_34_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07383_ _13651_/Q _07499_/A2 _07499_/B1 _14679_/Q _07382_/X vssd1 vssd1 vccd1 vccd1
+ _07383_/X sky130_fd_sc_hd__a221o_1
XFILLER_188_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09122_ _14239_/Q _14271_/Q _14303_/Q _14335_/Q _09190_/S _09429_/S1 vssd1 vssd1
+ vccd1 vccd1 _09122_/X sky130_fd_sc_hd__mux4_1
XFILLER_148_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09053_ _09130_/A _09046_/X _09049_/X _09450_/B1 vssd1 vssd1 vccd1 vccd1 _09053_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_159_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_536 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08004_ _08022_/B _08003_/X input35/X vssd1 vssd1 vccd1 vccd1 _08004_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_163_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09955_ _13098_/B2 _14315_/Q _09963_/S vssd1 vssd1 vccd1 vccd1 _14315_/D sky130_fd_sc_hd__mux2_1
XFILLER_132_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08906_ _09466_/A _08906_/B vssd1 vssd1 vccd1 vccd1 _08906_/X sky130_fd_sc_hd__or2_1
XTAP_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09886_ _13339_/A0 _14248_/Q _09897_/S vssd1 vssd1 vccd1 vccd1 _14248_/D sky130_fd_sc_hd__mux2_1
XTAP_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08837_ _13860_/Q _11761_/A0 _08851_/S vssd1 vssd1 vccd1 vccd1 _13860_/D sky130_fd_sc_hd__mux2_1
XFILLER_57_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08768_ _13125_/B _14612_/Q _08769_/B _08530_/B vssd1 vssd1 vccd1 vccd1 _08772_/B
+ sky130_fd_sc_hd__o31a_1
XTAP_2715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07719_ _14749_/Q _07713_/A _07718_/Y _07949_/C1 vssd1 vssd1 vccd1 vccd1 _13492_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_2748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08699_ _13587_/Q _08749_/A2 _08537_/Y _14493_/Q vssd1 vssd1 vccd1 vccd1 _08699_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_53_472 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10730_ _14764_/Q _10729_/X _10730_/S vssd1 vssd1 vccd1 vccd1 _14764_/D sky130_fd_sc_hd__mux2_1
XFILLER_159_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_848 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_122 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10661_ _15011_/Q _10569_/B _10733_/A2 _14979_/Q _10732_/C1 vssd1 vssd1 vccd1 vccd1
+ _10661_/X sky130_fd_sc_hd__a221o_1
X_12400_ _12595_/A1 _12395_/X _12398_/X _12399_/X _08405_/D vssd1 vssd1 vccd1 vccd1
+ _12412_/B sky130_fd_sc_hd__a221o_1
XFILLER_185_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13380_ _14483_/Q vssd1 vssd1 vccd1 vccd1 _14483_/D sky130_fd_sc_hd__clkbuf_2
X_10592_ _13716_/Q _10602_/B vssd1 vssd1 vccd1 vccd1 _10592_/X sky130_fd_sc_hd__and2_1
XFILLER_166_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12331_ _12618_/A1 _12326_/X _12329_/X _12330_/X _08405_/D vssd1 vssd1 vccd1 vccd1
+ _12343_/B sky130_fd_sc_hd__a221o_1
XFILLER_154_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12262_ _12273_/A1 _12257_/X _12260_/X _12261_/X _08449_/A vssd1 vssd1 vccd1 vccd1
+ _12274_/B sky130_fd_sc_hd__a221o_1
X_15050_ _15587_/CLK _15050_/D vssd1 vssd1 vccd1 vccd1 _15050_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_108_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11213_ _10382_/A _15002_/Q _11232_/S vssd1 vssd1 vccd1 vccd1 _15002_/D sky130_fd_sc_hd__mux2_1
X_14001_ _14420_/CLK _14001_/D vssd1 vssd1 vccd1 vccd1 _14001_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_579 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12193_ _12503_/A1 _12188_/X _12191_/X _12192_/X _08449_/A vssd1 vssd1 vccd1 vccd1
+ _12205_/B sky130_fd_sc_hd__a221o_1
Xoutput41 _07177_/X vssd1 vssd1 vccd1 vccd1 ext_address[15] sky130_fd_sc_hd__clkbuf_2
Xoutput52 _07188_/X vssd1 vssd1 vccd1 vccd1 ext_address[26] sky130_fd_sc_hd__clkbuf_2
X_11144_ _14972_/Q _10984_/Y _11141_/Y _11143_/Y vssd1 vssd1 vccd1 vccd1 _14972_/D
+ sky130_fd_sc_hd__a22o_1
Xoutput63 _07169_/X vssd1 vssd1 vccd1 vccd1 ext_address[7] sky130_fd_sc_hd__clkbuf_2
XFILLER_123_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput74 _07133_/X vssd1 vssd1 vccd1 vccd1 ext_write_data[16] sky130_fd_sc_hd__clkbuf_2
Xclkbuf_2_0_1_clk clkbuf_2_0_1_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_1_0_clk/A sky130_fd_sc_hd__clkbuf_8
XFILLER_68_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput85 _07153_/X vssd1 vssd1 vccd1 vccd1 ext_write_data[26] sky130_fd_sc_hd__clkbuf_2
XFILLER_150_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput96 _07115_/X vssd1 vssd1 vccd1 vccd1 ext_write_data[7] sky130_fd_sc_hd__clkbuf_2
XFILLER_122_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11075_ _11330_/A _11312_/A _11324_/B vssd1 vssd1 vccd1 vccd1 _11075_/X sky130_fd_sc_hd__and3_1
XFILLER_23_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10026_ _11847_/A1 _14384_/Q _10029_/S vssd1 vssd1 vccd1 vccd1 _14384_/D sky130_fd_sc_hd__mux2_1
XFILLER_48_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14903_ _15537_/CLK _14903_/D vssd1 vssd1 vccd1 vccd1 _14903_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_102_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14834_ _15508_/CLK _14834_/D vssd1 vssd1 vccd1 vccd1 _14834_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_36_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_940 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14765_ _15646_/CLK _14765_/D vssd1 vssd1 vccd1 vccd1 _14765_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_3994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11977_ _14232_/Q _14264_/Q _14296_/Q _14328_/Q _12154_/S _12253_/S1 vssd1 vssd1
+ vccd1 vccd1 _11977_/X sky130_fd_sc_hd__mux4_1
XFILLER_16_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13716_ _14997_/CLK _13716_/D vssd1 vssd1 vccd1 vccd1 _13716_/Q sky130_fd_sc_hd__dfxtp_1
X_10928_ _14947_/Q _10929_/B _10927_/Y _13208_/B vssd1 vssd1 vccd1 vccd1 _14947_/D
+ sky130_fd_sc_hd__o22a_1
X_14696_ _15643_/CLK _14696_/D vssd1 vssd1 vccd1 vccd1 _14696_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13647_ _13803_/CLK _13647_/D vssd1 vssd1 vccd1 vccd1 _13647_/Q sky130_fd_sc_hd__dfxtp_1
X_10859_ _14891_/Q _13777_/Q _12933_/S vssd1 vssd1 vccd1 vccd1 _14891_/D sky130_fd_sc_hd__mux2_1
XFILLER_31_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13578_ _14493_/CLK _13578_/D vssd1 vssd1 vccd1 vccd1 _13578_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_185_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15317_ _15497_/CLK _15317_/D vssd1 vssd1 vccd1 vccd1 _15317_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12529_ _14256_/Q _14288_/Q _14320_/Q _14352_/Q _12612_/S _12613_/A vssd1 vssd1 vccd1
+ vccd1 _12529_/X sky130_fd_sc_hd__mux4_1
XFILLER_117_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15248_ _15284_/CLK _15248_/D vssd1 vssd1 vccd1 vccd1 _15248_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_172_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15179_ _15220_/CLK _15179_/D vssd1 vssd1 vccd1 vccd1 _15179_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout308 _13338_/A0 vssd1 vssd1 vccd1 vccd1 _11838_/A1 sky130_fd_sc_hd__buf_6
Xfanout319 _07432_/X vssd1 vssd1 vccd1 vccd1 _13333_/A0 sky130_fd_sc_hd__buf_6
XFILLER_113_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09740_ _14108_/Q _11861_/A1 _09757_/S vssd1 vssd1 vccd1 vccd1 _14108_/D sky130_fd_sc_hd__mux2_1
X_06952_ _14490_/Q _06746_/Y _14489_/Q _06748_/Y _06948_/X vssd1 vssd1 vccd1 vccd1
+ _06952_/X sky130_fd_sc_hd__a221o_1
.ends

