// This is the unpowered netlist.
module core (clk,
    ext_instruction,
    ext_ready,
    ext_valid,
    meip,
    reset,
    ext_address,
    ext_read_data,
    ext_write_data,
    ext_write_strobe);
 input clk;
 output ext_instruction;
 input ext_ready;
 output ext_valid;
 input meip;
 input reset;
 output [31:0] ext_address;
 input [31:0] ext_read_data;
 output [31:0] ext_write_data;
 output [3:0] ext_write_strobe;

 wire net648;
 wire net649;
 wire net650;
 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire _06506_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06530_;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire _06559_;
 wire _06560_;
 wire _06561_;
 wire _06562_;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire _06571_;
 wire _06572_;
 wire _06573_;
 wire _06574_;
 wire _06575_;
 wire _06576_;
 wire _06577_;
 wire _06578_;
 wire _06579_;
 wire _06580_;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire _06584_;
 wire _06585_;
 wire _06586_;
 wire _06587_;
 wire _06588_;
 wire _06589_;
 wire _06590_;
 wire _06591_;
 wire _06592_;
 wire _06593_;
 wire _06594_;
 wire _06595_;
 wire _06596_;
 wire _06597_;
 wire _06598_;
 wire _06599_;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire _06603_;
 wire _06604_;
 wire _06605_;
 wire _06606_;
 wire _06607_;
 wire _06608_;
 wire _06609_;
 wire _06610_;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire _06616_;
 wire _06617_;
 wire _06618_;
 wire _06619_;
 wire _06620_;
 wire _06621_;
 wire _06622_;
 wire _06623_;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire _06655_;
 wire _06656_;
 wire _06657_;
 wire clknet_0_clk;
 wire clknet_1_0_0_clk;
 wire clknet_1_0_1_clk;
 wire clknet_1_1_0_clk;
 wire clknet_1_1_1_clk;
 wire clknet_2_0_0_clk;
 wire clknet_2_0_1_clk;
 wire clknet_2_1_0_clk;
 wire clknet_2_1_1_clk;
 wire clknet_2_2_0_clk;
 wire clknet_2_2_1_clk;
 wire clknet_2_3_0_clk;
 wire clknet_2_3_1_clk;
 wire clknet_3_0_0_clk;
 wire clknet_3_1_0_clk;
 wire clknet_3_2_0_clk;
 wire clknet_3_3_0_clk;
 wire clknet_3_4_0_clk;
 wire clknet_3_5_0_clk;
 wire clknet_3_6_0_clk;
 wire clknet_3_7_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_5_0_0_clk;
 wire clknet_5_10_0_clk;
 wire clknet_5_11_0_clk;
 wire clknet_5_12_0_clk;
 wire clknet_5_13_0_clk;
 wire clknet_5_14_0_clk;
 wire clknet_5_15_0_clk;
 wire clknet_5_16_0_clk;
 wire clknet_5_17_0_clk;
 wire clknet_5_18_0_clk;
 wire clknet_5_19_0_clk;
 wire clknet_5_1_0_clk;
 wire clknet_5_20_0_clk;
 wire clknet_5_21_0_clk;
 wire clknet_5_22_0_clk;
 wire clknet_5_23_0_clk;
 wire clknet_5_24_0_clk;
 wire clknet_5_25_0_clk;
 wire clknet_5_26_0_clk;
 wire clknet_5_27_0_clk;
 wire clknet_5_28_0_clk;
 wire clknet_5_29_0_clk;
 wire clknet_5_2_0_clk;
 wire clknet_5_30_0_clk;
 wire clknet_5_31_0_clk;
 wire clknet_5_3_0_clk;
 wire clknet_5_4_0_clk;
 wire clknet_5_5_0_clk;
 wire clknet_5_6_0_clk;
 wire clknet_5_7_0_clk;
 wire clknet_5_8_0_clk;
 wire clknet_5_9_0_clk;
 wire clknet_leaf_0_clk;
 wire clknet_leaf_100_clk;
 wire clknet_leaf_101_clk;
 wire clknet_leaf_102_clk;
 wire clknet_leaf_103_clk;
 wire clknet_leaf_104_clk;
 wire clknet_leaf_105_clk;
 wire clknet_leaf_106_clk;
 wire clknet_leaf_107_clk;
 wire clknet_leaf_108_clk;
 wire clknet_leaf_109_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_110_clk;
 wire clknet_leaf_111_clk;
 wire clknet_leaf_113_clk;
 wire clknet_leaf_114_clk;
 wire clknet_leaf_115_clk;
 wire clknet_leaf_116_clk;
 wire clknet_leaf_117_clk;
 wire clknet_leaf_118_clk;
 wire clknet_leaf_119_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_120_clk;
 wire clknet_leaf_121_clk;
 wire clknet_leaf_122_clk;
 wire clknet_leaf_123_clk;
 wire clknet_leaf_124_clk;
 wire clknet_leaf_125_clk;
 wire clknet_leaf_126_clk;
 wire clknet_leaf_127_clk;
 wire clknet_leaf_128_clk;
 wire clknet_leaf_129_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_130_clk;
 wire clknet_leaf_131_clk;
 wire clknet_leaf_132_clk;
 wire clknet_leaf_133_clk;
 wire clknet_leaf_134_clk;
 wire clknet_leaf_135_clk;
 wire clknet_leaf_136_clk;
 wire clknet_leaf_137_clk;
 wire clknet_leaf_138_clk;
 wire clknet_leaf_139_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_140_clk;
 wire clknet_leaf_141_clk;
 wire clknet_leaf_142_clk;
 wire clknet_leaf_143_clk;
 wire clknet_leaf_144_clk;
 wire clknet_leaf_145_clk;
 wire clknet_leaf_146_clk;
 wire clknet_leaf_147_clk;
 wire clknet_leaf_148_clk;
 wire clknet_leaf_149_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_150_clk;
 wire clknet_leaf_151_clk;
 wire clknet_leaf_152_clk;
 wire clknet_leaf_153_clk;
 wire clknet_leaf_154_clk;
 wire clknet_leaf_155_clk;
 wire clknet_leaf_156_clk;
 wire clknet_leaf_157_clk;
 wire clknet_leaf_158_clk;
 wire clknet_leaf_159_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_160_clk;
 wire clknet_leaf_161_clk;
 wire clknet_leaf_162_clk;
 wire clknet_leaf_163_clk;
 wire clknet_leaf_164_clk;
 wire clknet_leaf_165_clk;
 wire clknet_leaf_166_clk;
 wire clknet_leaf_167_clk;
 wire clknet_leaf_168_clk;
 wire clknet_leaf_169_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_170_clk;
 wire clknet_leaf_171_clk;
 wire clknet_leaf_172_clk;
 wire clknet_leaf_173_clk;
 wire clknet_leaf_174_clk;
 wire clknet_leaf_175_clk;
 wire clknet_leaf_176_clk;
 wire clknet_leaf_177_clk;
 wire clknet_leaf_178_clk;
 wire clknet_leaf_179_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_180_clk;
 wire clknet_leaf_181_clk;
 wire clknet_leaf_182_clk;
 wire clknet_leaf_183_clk;
 wire clknet_leaf_184_clk;
 wire clknet_leaf_185_clk;
 wire clknet_leaf_186_clk;
 wire clknet_leaf_187_clk;
 wire clknet_leaf_188_clk;
 wire clknet_leaf_189_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_190_clk;
 wire clknet_leaf_191_clk;
 wire clknet_leaf_192_clk;
 wire clknet_leaf_193_clk;
 wire clknet_leaf_194_clk;
 wire clknet_leaf_195_clk;
 wire clknet_leaf_196_clk;
 wire clknet_leaf_197_clk;
 wire clknet_leaf_198_clk;
 wire clknet_leaf_199_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_200_clk;
 wire clknet_leaf_201_clk;
 wire clknet_leaf_202_clk;
 wire clknet_leaf_203_clk;
 wire clknet_leaf_204_clk;
 wire clknet_leaf_205_clk;
 wire clknet_leaf_206_clk;
 wire clknet_leaf_207_clk;
 wire clknet_leaf_208_clk;
 wire clknet_leaf_209_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_210_clk;
 wire clknet_leaf_211_clk;
 wire clknet_leaf_212_clk;
 wire clknet_leaf_213_clk;
 wire clknet_leaf_214_clk;
 wire clknet_leaf_215_clk;
 wire clknet_leaf_216_clk;
 wire clknet_leaf_217_clk;
 wire clknet_leaf_218_clk;
 wire clknet_leaf_219_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_220_clk;
 wire clknet_leaf_221_clk;
 wire clknet_leaf_222_clk;
 wire clknet_leaf_223_clk;
 wire clknet_leaf_224_clk;
 wire clknet_leaf_225_clk;
 wire clknet_leaf_226_clk;
 wire clknet_leaf_227_clk;
 wire clknet_leaf_228_clk;
 wire clknet_leaf_229_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_230_clk;
 wire clknet_leaf_231_clk;
 wire clknet_leaf_232_clk;
 wire clknet_leaf_233_clk;
 wire clknet_leaf_234_clk;
 wire clknet_leaf_235_clk;
 wire clknet_leaf_236_clk;
 wire clknet_leaf_237_clk;
 wire clknet_leaf_238_clk;
 wire clknet_leaf_239_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_240_clk;
 wire clknet_leaf_241_clk;
 wire clknet_leaf_242_clk;
 wire clknet_leaf_243_clk;
 wire clknet_leaf_244_clk;
 wire clknet_leaf_245_clk;
 wire clknet_leaf_246_clk;
 wire clknet_leaf_247_clk;
 wire clknet_leaf_248_clk;
 wire clknet_leaf_249_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_250_clk;
 wire clknet_leaf_251_clk;
 wire clknet_leaf_252_clk;
 wire clknet_leaf_253_clk;
 wire clknet_leaf_254_clk;
 wire clknet_leaf_255_clk;
 wire clknet_leaf_256_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_55_clk;
 wire clknet_leaf_56_clk;
 wire clknet_leaf_57_clk;
 wire clknet_leaf_58_clk;
 wire clknet_leaf_59_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_60_clk;
 wire clknet_leaf_61_clk;
 wire clknet_leaf_62_clk;
 wire clknet_leaf_63_clk;
 wire clknet_leaf_64_clk;
 wire clknet_leaf_65_clk;
 wire clknet_leaf_66_clk;
 wire clknet_leaf_67_clk;
 wire clknet_leaf_68_clk;
 wire clknet_leaf_69_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_70_clk;
 wire clknet_leaf_71_clk;
 wire clknet_leaf_72_clk;
 wire clknet_leaf_73_clk;
 wire clknet_leaf_74_clk;
 wire clknet_leaf_75_clk;
 wire clknet_leaf_76_clk;
 wire clknet_leaf_77_clk;
 wire clknet_leaf_78_clk;
 wire clknet_leaf_79_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_80_clk;
 wire clknet_leaf_81_clk;
 wire clknet_leaf_82_clk;
 wire clknet_leaf_83_clk;
 wire clknet_leaf_84_clk;
 wire clknet_leaf_85_clk;
 wire clknet_leaf_86_clk;
 wire clknet_leaf_87_clk;
 wire clknet_leaf_88_clk;
 wire clknet_leaf_89_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_90_clk;
 wire clknet_leaf_91_clk;
 wire clknet_leaf_92_clk;
 wire clknet_leaf_93_clk;
 wire clknet_leaf_94_clk;
 wire clknet_leaf_95_clk;
 wire clknet_leaf_96_clk;
 wire clknet_leaf_97_clk;
 wire clknet_leaf_98_clk;
 wire clknet_leaf_99_clk;
 wire clknet_leaf_9_clk;
 wire clknet_opt_1_0_clk;
 wire clknet_opt_2_0_clk;
 wire \core_busio.mem_address[0] ;
 wire \core_busio.mem_address[10] ;
 wire \core_busio.mem_address[11] ;
 wire \core_busio.mem_address[12] ;
 wire \core_busio.mem_address[13] ;
 wire \core_busio.mem_address[14] ;
 wire \core_busio.mem_address[15] ;
 wire \core_busio.mem_address[16] ;
 wire \core_busio.mem_address[17] ;
 wire \core_busio.mem_address[18] ;
 wire \core_busio.mem_address[19] ;
 wire \core_busio.mem_address[1] ;
 wire \core_busio.mem_address[20] ;
 wire \core_busio.mem_address[21] ;
 wire \core_busio.mem_address[22] ;
 wire \core_busio.mem_address[23] ;
 wire \core_busio.mem_address[24] ;
 wire \core_busio.mem_address[25] ;
 wire \core_busio.mem_address[26] ;
 wire \core_busio.mem_address[27] ;
 wire \core_busio.mem_address[28] ;
 wire \core_busio.mem_address[29] ;
 wire \core_busio.mem_address[2] ;
 wire \core_busio.mem_address[30] ;
 wire \core_busio.mem_address[31] ;
 wire \core_busio.mem_address[3] ;
 wire \core_busio.mem_address[4] ;
 wire \core_busio.mem_address[5] ;
 wire \core_busio.mem_address[6] ;
 wire \core_busio.mem_address[7] ;
 wire \core_busio.mem_address[8] ;
 wire \core_busio.mem_address[9] ;
 wire \core_busio.mem_signed ;
 wire \core_busio.mem_size[0] ;
 wire \core_busio.mem_size[1] ;
 wire \core_busio.mem_store_data[0] ;
 wire \core_busio.mem_store_data[10] ;
 wire \core_busio.mem_store_data[11] ;
 wire \core_busio.mem_store_data[12] ;
 wire \core_busio.mem_store_data[13] ;
 wire \core_busio.mem_store_data[14] ;
 wire \core_busio.mem_store_data[15] ;
 wire \core_busio.mem_store_data[16] ;
 wire \core_busio.mem_store_data[17] ;
 wire \core_busio.mem_store_data[18] ;
 wire \core_busio.mem_store_data[19] ;
 wire \core_busio.mem_store_data[1] ;
 wire \core_busio.mem_store_data[20] ;
 wire \core_busio.mem_store_data[21] ;
 wire \core_busio.mem_store_data[22] ;
 wire \core_busio.mem_store_data[23] ;
 wire \core_busio.mem_store_data[24] ;
 wire \core_busio.mem_store_data[25] ;
 wire \core_busio.mem_store_data[26] ;
 wire \core_busio.mem_store_data[27] ;
 wire \core_busio.mem_store_data[28] ;
 wire \core_busio.mem_store_data[29] ;
 wire \core_busio.mem_store_data[2] ;
 wire \core_busio.mem_store_data[30] ;
 wire \core_busio.mem_store_data[31] ;
 wire \core_busio.mem_store_data[3] ;
 wire \core_busio.mem_store_data[4] ;
 wire \core_busio.mem_store_data[5] ;
 wire \core_busio.mem_store_data[6] ;
 wire \core_busio.mem_store_data[7] ;
 wire \core_busio.mem_store_data[8] ;
 wire \core_busio.mem_store_data[9] ;
 wire \core_pipeline.csr_to_fetch_mret_vector[0] ;
 wire \core_pipeline.csr_to_fetch_mret_vector[10] ;
 wire \core_pipeline.csr_to_fetch_mret_vector[11] ;
 wire \core_pipeline.csr_to_fetch_mret_vector[12] ;
 wire \core_pipeline.csr_to_fetch_mret_vector[13] ;
 wire \core_pipeline.csr_to_fetch_mret_vector[14] ;
 wire \core_pipeline.csr_to_fetch_mret_vector[15] ;
 wire \core_pipeline.csr_to_fetch_mret_vector[16] ;
 wire \core_pipeline.csr_to_fetch_mret_vector[17] ;
 wire \core_pipeline.csr_to_fetch_mret_vector[18] ;
 wire \core_pipeline.csr_to_fetch_mret_vector[19] ;
 wire \core_pipeline.csr_to_fetch_mret_vector[1] ;
 wire \core_pipeline.csr_to_fetch_mret_vector[20] ;
 wire \core_pipeline.csr_to_fetch_mret_vector[21] ;
 wire \core_pipeline.csr_to_fetch_mret_vector[22] ;
 wire \core_pipeline.csr_to_fetch_mret_vector[23] ;
 wire \core_pipeline.csr_to_fetch_mret_vector[24] ;
 wire \core_pipeline.csr_to_fetch_mret_vector[25] ;
 wire \core_pipeline.csr_to_fetch_mret_vector[26] ;
 wire \core_pipeline.csr_to_fetch_mret_vector[27] ;
 wire \core_pipeline.csr_to_fetch_mret_vector[28] ;
 wire \core_pipeline.csr_to_fetch_mret_vector[29] ;
 wire \core_pipeline.csr_to_fetch_mret_vector[2] ;
 wire \core_pipeline.csr_to_fetch_mret_vector[30] ;
 wire \core_pipeline.csr_to_fetch_mret_vector[31] ;
 wire \core_pipeline.csr_to_fetch_mret_vector[3] ;
 wire \core_pipeline.csr_to_fetch_mret_vector[4] ;
 wire \core_pipeline.csr_to_fetch_mret_vector[5] ;
 wire \core_pipeline.csr_to_fetch_mret_vector[6] ;
 wire \core_pipeline.csr_to_fetch_mret_vector[7] ;
 wire \core_pipeline.csr_to_fetch_mret_vector[8] ;
 wire \core_pipeline.csr_to_fetch_mret_vector[9] ;
 wire \core_pipeline.csr_to_fetch_trap_vector[10] ;
 wire \core_pipeline.csr_to_fetch_trap_vector[11] ;
 wire \core_pipeline.csr_to_fetch_trap_vector[12] ;
 wire \core_pipeline.csr_to_fetch_trap_vector[13] ;
 wire \core_pipeline.csr_to_fetch_trap_vector[14] ;
 wire \core_pipeline.csr_to_fetch_trap_vector[15] ;
 wire \core_pipeline.csr_to_fetch_trap_vector[16] ;
 wire \core_pipeline.csr_to_fetch_trap_vector[17] ;
 wire \core_pipeline.csr_to_fetch_trap_vector[18] ;
 wire \core_pipeline.csr_to_fetch_trap_vector[19] ;
 wire \core_pipeline.csr_to_fetch_trap_vector[20] ;
 wire \core_pipeline.csr_to_fetch_trap_vector[21] ;
 wire \core_pipeline.csr_to_fetch_trap_vector[22] ;
 wire \core_pipeline.csr_to_fetch_trap_vector[23] ;
 wire \core_pipeline.csr_to_fetch_trap_vector[24] ;
 wire \core_pipeline.csr_to_fetch_trap_vector[25] ;
 wire \core_pipeline.csr_to_fetch_trap_vector[26] ;
 wire \core_pipeline.csr_to_fetch_trap_vector[27] ;
 wire \core_pipeline.csr_to_fetch_trap_vector[28] ;
 wire \core_pipeline.csr_to_fetch_trap_vector[29] ;
 wire \core_pipeline.csr_to_fetch_trap_vector[2] ;
 wire \core_pipeline.csr_to_fetch_trap_vector[30] ;
 wire \core_pipeline.csr_to_fetch_trap_vector[31] ;
 wire \core_pipeline.csr_to_fetch_trap_vector[3] ;
 wire \core_pipeline.csr_to_fetch_trap_vector[4] ;
 wire \core_pipeline.csr_to_fetch_trap_vector[5] ;
 wire \core_pipeline.csr_to_fetch_trap_vector[6] ;
 wire \core_pipeline.csr_to_fetch_trap_vector[7] ;
 wire \core_pipeline.csr_to_fetch_trap_vector[8] ;
 wire \core_pipeline.csr_to_fetch_trap_vector[9] ;
 wire \core_pipeline.decode_to_csr_read_address[0] ;
 wire \core_pipeline.decode_to_csr_read_address[10] ;
 wire \core_pipeline.decode_to_csr_read_address[11] ;
 wire \core_pipeline.decode_to_csr_read_address[1] ;
 wire \core_pipeline.decode_to_csr_read_address[2] ;
 wire \core_pipeline.decode_to_csr_read_address[3] ;
 wire \core_pipeline.decode_to_csr_read_address[4] ;
 wire \core_pipeline.decode_to_csr_read_address[5] ;
 wire \core_pipeline.decode_to_csr_read_address[6] ;
 wire \core_pipeline.decode_to_csr_read_address[7] ;
 wire \core_pipeline.decode_to_csr_read_address[8] ;
 wire \core_pipeline.decode_to_csr_read_address[9] ;
 wire \core_pipeline.decode_to_execute_alu_function[0] ;
 wire \core_pipeline.decode_to_execute_alu_function[1] ;
 wire \core_pipeline.decode_to_execute_alu_function[2] ;
 wire \core_pipeline.decode_to_execute_alu_function_modifier ;
 wire \core_pipeline.decode_to_execute_branch ;
 wire \core_pipeline.decode_to_execute_bypass_memory ;
 wire \core_pipeline.decode_to_execute_cmp_function[0] ;
 wire \core_pipeline.decode_to_execute_cmp_function[1] ;
 wire \core_pipeline.decode_to_execute_cmp_function[2] ;
 wire \core_pipeline.decode_to_execute_csr_address[0] ;
 wire \core_pipeline.decode_to_execute_csr_address[10] ;
 wire \core_pipeline.decode_to_execute_csr_address[11] ;
 wire \core_pipeline.decode_to_execute_csr_address[1] ;
 wire \core_pipeline.decode_to_execute_csr_address[2] ;
 wire \core_pipeline.decode_to_execute_csr_address[3] ;
 wire \core_pipeline.decode_to_execute_csr_address[4] ;
 wire \core_pipeline.decode_to_execute_csr_address[5] ;
 wire \core_pipeline.decode_to_execute_csr_address[6] ;
 wire \core_pipeline.decode_to_execute_csr_address[7] ;
 wire \core_pipeline.decode_to_execute_csr_address[8] ;
 wire \core_pipeline.decode_to_execute_csr_address[9] ;
 wire \core_pipeline.decode_to_execute_csr_data[0] ;
 wire \core_pipeline.decode_to_execute_csr_data[10] ;
 wire \core_pipeline.decode_to_execute_csr_data[11] ;
 wire \core_pipeline.decode_to_execute_csr_data[12] ;
 wire \core_pipeline.decode_to_execute_csr_data[13] ;
 wire \core_pipeline.decode_to_execute_csr_data[14] ;
 wire \core_pipeline.decode_to_execute_csr_data[15] ;
 wire \core_pipeline.decode_to_execute_csr_data[16] ;
 wire \core_pipeline.decode_to_execute_csr_data[17] ;
 wire \core_pipeline.decode_to_execute_csr_data[18] ;
 wire \core_pipeline.decode_to_execute_csr_data[19] ;
 wire \core_pipeline.decode_to_execute_csr_data[1] ;
 wire \core_pipeline.decode_to_execute_csr_data[20] ;
 wire \core_pipeline.decode_to_execute_csr_data[21] ;
 wire \core_pipeline.decode_to_execute_csr_data[22] ;
 wire \core_pipeline.decode_to_execute_csr_data[23] ;
 wire \core_pipeline.decode_to_execute_csr_data[24] ;
 wire \core_pipeline.decode_to_execute_csr_data[25] ;
 wire \core_pipeline.decode_to_execute_csr_data[26] ;
 wire \core_pipeline.decode_to_execute_csr_data[27] ;
 wire \core_pipeline.decode_to_execute_csr_data[28] ;
 wire \core_pipeline.decode_to_execute_csr_data[29] ;
 wire \core_pipeline.decode_to_execute_csr_data[2] ;
 wire \core_pipeline.decode_to_execute_csr_data[30] ;
 wire \core_pipeline.decode_to_execute_csr_data[31] ;
 wire \core_pipeline.decode_to_execute_csr_data[3] ;
 wire \core_pipeline.decode_to_execute_csr_data[4] ;
 wire \core_pipeline.decode_to_execute_csr_data[5] ;
 wire \core_pipeline.decode_to_execute_csr_data[6] ;
 wire \core_pipeline.decode_to_execute_csr_data[7] ;
 wire \core_pipeline.decode_to_execute_csr_data[8] ;
 wire \core_pipeline.decode_to_execute_csr_data[9] ;
 wire \core_pipeline.decode_to_execute_csr_read ;
 wire \core_pipeline.decode_to_execute_csr_readable ;
 wire \core_pipeline.decode_to_execute_csr_write ;
 wire \core_pipeline.decode_to_execute_csr_writeable ;
 wire \core_pipeline.decode_to_execute_ecause[0] ;
 wire \core_pipeline.decode_to_execute_ecause[1] ;
 wire \core_pipeline.decode_to_execute_ecause[3] ;
 wire \core_pipeline.decode_to_execute_exception ;
 wire \core_pipeline.decode_to_execute_imm_data[0] ;
 wire \core_pipeline.decode_to_execute_imm_data[10] ;
 wire \core_pipeline.decode_to_execute_imm_data[11] ;
 wire \core_pipeline.decode_to_execute_imm_data[12] ;
 wire \core_pipeline.decode_to_execute_imm_data[13] ;
 wire \core_pipeline.decode_to_execute_imm_data[14] ;
 wire \core_pipeline.decode_to_execute_imm_data[15] ;
 wire \core_pipeline.decode_to_execute_imm_data[16] ;
 wire \core_pipeline.decode_to_execute_imm_data[17] ;
 wire \core_pipeline.decode_to_execute_imm_data[18] ;
 wire \core_pipeline.decode_to_execute_imm_data[19] ;
 wire \core_pipeline.decode_to_execute_imm_data[1] ;
 wire \core_pipeline.decode_to_execute_imm_data[20] ;
 wire \core_pipeline.decode_to_execute_imm_data[21] ;
 wire \core_pipeline.decode_to_execute_imm_data[22] ;
 wire \core_pipeline.decode_to_execute_imm_data[23] ;
 wire \core_pipeline.decode_to_execute_imm_data[24] ;
 wire \core_pipeline.decode_to_execute_imm_data[25] ;
 wire \core_pipeline.decode_to_execute_imm_data[26] ;
 wire \core_pipeline.decode_to_execute_imm_data[27] ;
 wire \core_pipeline.decode_to_execute_imm_data[28] ;
 wire \core_pipeline.decode_to_execute_imm_data[29] ;
 wire \core_pipeline.decode_to_execute_imm_data[2] ;
 wire \core_pipeline.decode_to_execute_imm_data[30] ;
 wire \core_pipeline.decode_to_execute_imm_data[31] ;
 wire \core_pipeline.decode_to_execute_imm_data[3] ;
 wire \core_pipeline.decode_to_execute_imm_data[4] ;
 wire \core_pipeline.decode_to_execute_imm_data[5] ;
 wire \core_pipeline.decode_to_execute_imm_data[6] ;
 wire \core_pipeline.decode_to_execute_imm_data[7] ;
 wire \core_pipeline.decode_to_execute_imm_data[8] ;
 wire \core_pipeline.decode_to_execute_imm_data[9] ;
 wire \core_pipeline.decode_to_execute_jump ;
 wire \core_pipeline.decode_to_execute_load ;
 wire \core_pipeline.decode_to_execute_load_signed ;
 wire \core_pipeline.decode_to_execute_mret ;
 wire \core_pipeline.decode_to_execute_next_pc[0] ;
 wire \core_pipeline.decode_to_execute_next_pc[10] ;
 wire \core_pipeline.decode_to_execute_next_pc[11] ;
 wire \core_pipeline.decode_to_execute_next_pc[12] ;
 wire \core_pipeline.decode_to_execute_next_pc[13] ;
 wire \core_pipeline.decode_to_execute_next_pc[14] ;
 wire \core_pipeline.decode_to_execute_next_pc[15] ;
 wire \core_pipeline.decode_to_execute_next_pc[16] ;
 wire \core_pipeline.decode_to_execute_next_pc[17] ;
 wire \core_pipeline.decode_to_execute_next_pc[18] ;
 wire \core_pipeline.decode_to_execute_next_pc[19] ;
 wire \core_pipeline.decode_to_execute_next_pc[1] ;
 wire \core_pipeline.decode_to_execute_next_pc[20] ;
 wire \core_pipeline.decode_to_execute_next_pc[21] ;
 wire \core_pipeline.decode_to_execute_next_pc[22] ;
 wire \core_pipeline.decode_to_execute_next_pc[23] ;
 wire \core_pipeline.decode_to_execute_next_pc[24] ;
 wire \core_pipeline.decode_to_execute_next_pc[25] ;
 wire \core_pipeline.decode_to_execute_next_pc[26] ;
 wire \core_pipeline.decode_to_execute_next_pc[27] ;
 wire \core_pipeline.decode_to_execute_next_pc[28] ;
 wire \core_pipeline.decode_to_execute_next_pc[29] ;
 wire \core_pipeline.decode_to_execute_next_pc[2] ;
 wire \core_pipeline.decode_to_execute_next_pc[30] ;
 wire \core_pipeline.decode_to_execute_next_pc[31] ;
 wire \core_pipeline.decode_to_execute_next_pc[3] ;
 wire \core_pipeline.decode_to_execute_next_pc[4] ;
 wire \core_pipeline.decode_to_execute_next_pc[5] ;
 wire \core_pipeline.decode_to_execute_next_pc[6] ;
 wire \core_pipeline.decode_to_execute_next_pc[7] ;
 wire \core_pipeline.decode_to_execute_next_pc[8] ;
 wire \core_pipeline.decode_to_execute_next_pc[9] ;
 wire \core_pipeline.decode_to_execute_pc[10] ;
 wire \core_pipeline.decode_to_execute_pc[11] ;
 wire \core_pipeline.decode_to_execute_pc[12] ;
 wire \core_pipeline.decode_to_execute_pc[13] ;
 wire \core_pipeline.decode_to_execute_pc[14] ;
 wire \core_pipeline.decode_to_execute_pc[15] ;
 wire \core_pipeline.decode_to_execute_pc[16] ;
 wire \core_pipeline.decode_to_execute_pc[17] ;
 wire \core_pipeline.decode_to_execute_pc[18] ;
 wire \core_pipeline.decode_to_execute_pc[19] ;
 wire \core_pipeline.decode_to_execute_pc[20] ;
 wire \core_pipeline.decode_to_execute_pc[21] ;
 wire \core_pipeline.decode_to_execute_pc[22] ;
 wire \core_pipeline.decode_to_execute_pc[23] ;
 wire \core_pipeline.decode_to_execute_pc[24] ;
 wire \core_pipeline.decode_to_execute_pc[25] ;
 wire \core_pipeline.decode_to_execute_pc[26] ;
 wire \core_pipeline.decode_to_execute_pc[27] ;
 wire \core_pipeline.decode_to_execute_pc[28] ;
 wire \core_pipeline.decode_to_execute_pc[29] ;
 wire \core_pipeline.decode_to_execute_pc[2] ;
 wire \core_pipeline.decode_to_execute_pc[30] ;
 wire \core_pipeline.decode_to_execute_pc[31] ;
 wire \core_pipeline.decode_to_execute_pc[3] ;
 wire \core_pipeline.decode_to_execute_pc[4] ;
 wire \core_pipeline.decode_to_execute_pc[5] ;
 wire \core_pipeline.decode_to_execute_pc[6] ;
 wire \core_pipeline.decode_to_execute_pc[7] ;
 wire \core_pipeline.decode_to_execute_pc[8] ;
 wire \core_pipeline.decode_to_execute_pc[9] ;
 wire \core_pipeline.decode_to_execute_rd_address[0] ;
 wire \core_pipeline.decode_to_execute_rd_address[1] ;
 wire \core_pipeline.decode_to_execute_rd_address[2] ;
 wire \core_pipeline.decode_to_execute_rd_address[3] ;
 wire \core_pipeline.decode_to_execute_rd_address[4] ;
 wire \core_pipeline.decode_to_execute_rs1_bypass[0] ;
 wire \core_pipeline.decode_to_execute_rs1_bypass[10] ;
 wire \core_pipeline.decode_to_execute_rs1_bypass[11] ;
 wire \core_pipeline.decode_to_execute_rs1_bypass[12] ;
 wire \core_pipeline.decode_to_execute_rs1_bypass[13] ;
 wire \core_pipeline.decode_to_execute_rs1_bypass[14] ;
 wire \core_pipeline.decode_to_execute_rs1_bypass[15] ;
 wire \core_pipeline.decode_to_execute_rs1_bypass[16] ;
 wire \core_pipeline.decode_to_execute_rs1_bypass[17] ;
 wire \core_pipeline.decode_to_execute_rs1_bypass[18] ;
 wire \core_pipeline.decode_to_execute_rs1_bypass[19] ;
 wire \core_pipeline.decode_to_execute_rs1_bypass[1] ;
 wire \core_pipeline.decode_to_execute_rs1_bypass[20] ;
 wire \core_pipeline.decode_to_execute_rs1_bypass[21] ;
 wire \core_pipeline.decode_to_execute_rs1_bypass[22] ;
 wire \core_pipeline.decode_to_execute_rs1_bypass[23] ;
 wire \core_pipeline.decode_to_execute_rs1_bypass[24] ;
 wire \core_pipeline.decode_to_execute_rs1_bypass[25] ;
 wire \core_pipeline.decode_to_execute_rs1_bypass[26] ;
 wire \core_pipeline.decode_to_execute_rs1_bypass[27] ;
 wire \core_pipeline.decode_to_execute_rs1_bypass[28] ;
 wire \core_pipeline.decode_to_execute_rs1_bypass[29] ;
 wire \core_pipeline.decode_to_execute_rs1_bypass[2] ;
 wire \core_pipeline.decode_to_execute_rs1_bypass[30] ;
 wire \core_pipeline.decode_to_execute_rs1_bypass[31] ;
 wire \core_pipeline.decode_to_execute_rs1_bypass[3] ;
 wire \core_pipeline.decode_to_execute_rs1_bypass[4] ;
 wire \core_pipeline.decode_to_execute_rs1_bypass[5] ;
 wire \core_pipeline.decode_to_execute_rs1_bypass[6] ;
 wire \core_pipeline.decode_to_execute_rs1_bypass[7] ;
 wire \core_pipeline.decode_to_execute_rs1_bypass[8] ;
 wire \core_pipeline.decode_to_execute_rs1_bypass[9] ;
 wire \core_pipeline.decode_to_execute_rs1_bypassed ;
 wire \core_pipeline.decode_to_execute_rs1_data[0] ;
 wire \core_pipeline.decode_to_execute_rs1_data[10] ;
 wire \core_pipeline.decode_to_execute_rs1_data[11] ;
 wire \core_pipeline.decode_to_execute_rs1_data[12] ;
 wire \core_pipeline.decode_to_execute_rs1_data[13] ;
 wire \core_pipeline.decode_to_execute_rs1_data[14] ;
 wire \core_pipeline.decode_to_execute_rs1_data[15] ;
 wire \core_pipeline.decode_to_execute_rs1_data[16] ;
 wire \core_pipeline.decode_to_execute_rs1_data[17] ;
 wire \core_pipeline.decode_to_execute_rs1_data[18] ;
 wire \core_pipeline.decode_to_execute_rs1_data[19] ;
 wire \core_pipeline.decode_to_execute_rs1_data[1] ;
 wire \core_pipeline.decode_to_execute_rs1_data[20] ;
 wire \core_pipeline.decode_to_execute_rs1_data[21] ;
 wire \core_pipeline.decode_to_execute_rs1_data[22] ;
 wire \core_pipeline.decode_to_execute_rs1_data[23] ;
 wire \core_pipeline.decode_to_execute_rs1_data[24] ;
 wire \core_pipeline.decode_to_execute_rs1_data[25] ;
 wire \core_pipeline.decode_to_execute_rs1_data[26] ;
 wire \core_pipeline.decode_to_execute_rs1_data[27] ;
 wire \core_pipeline.decode_to_execute_rs1_data[28] ;
 wire \core_pipeline.decode_to_execute_rs1_data[29] ;
 wire \core_pipeline.decode_to_execute_rs1_data[2] ;
 wire \core_pipeline.decode_to_execute_rs1_data[30] ;
 wire \core_pipeline.decode_to_execute_rs1_data[31] ;
 wire \core_pipeline.decode_to_execute_rs1_data[3] ;
 wire \core_pipeline.decode_to_execute_rs1_data[4] ;
 wire \core_pipeline.decode_to_execute_rs1_data[5] ;
 wire \core_pipeline.decode_to_execute_rs1_data[6] ;
 wire \core_pipeline.decode_to_execute_rs1_data[7] ;
 wire \core_pipeline.decode_to_execute_rs1_data[8] ;
 wire \core_pipeline.decode_to_execute_rs1_data[9] ;
 wire \core_pipeline.decode_to_execute_rs2_bypass[0] ;
 wire \core_pipeline.decode_to_execute_rs2_bypass[10] ;
 wire \core_pipeline.decode_to_execute_rs2_bypass[11] ;
 wire \core_pipeline.decode_to_execute_rs2_bypass[12] ;
 wire \core_pipeline.decode_to_execute_rs2_bypass[13] ;
 wire \core_pipeline.decode_to_execute_rs2_bypass[14] ;
 wire \core_pipeline.decode_to_execute_rs2_bypass[15] ;
 wire \core_pipeline.decode_to_execute_rs2_bypass[16] ;
 wire \core_pipeline.decode_to_execute_rs2_bypass[17] ;
 wire \core_pipeline.decode_to_execute_rs2_bypass[18] ;
 wire \core_pipeline.decode_to_execute_rs2_bypass[19] ;
 wire \core_pipeline.decode_to_execute_rs2_bypass[1] ;
 wire \core_pipeline.decode_to_execute_rs2_bypass[20] ;
 wire \core_pipeline.decode_to_execute_rs2_bypass[21] ;
 wire \core_pipeline.decode_to_execute_rs2_bypass[22] ;
 wire \core_pipeline.decode_to_execute_rs2_bypass[23] ;
 wire \core_pipeline.decode_to_execute_rs2_bypass[24] ;
 wire \core_pipeline.decode_to_execute_rs2_bypass[25] ;
 wire \core_pipeline.decode_to_execute_rs2_bypass[26] ;
 wire \core_pipeline.decode_to_execute_rs2_bypass[27] ;
 wire \core_pipeline.decode_to_execute_rs2_bypass[28] ;
 wire \core_pipeline.decode_to_execute_rs2_bypass[29] ;
 wire \core_pipeline.decode_to_execute_rs2_bypass[2] ;
 wire \core_pipeline.decode_to_execute_rs2_bypass[30] ;
 wire \core_pipeline.decode_to_execute_rs2_bypass[31] ;
 wire \core_pipeline.decode_to_execute_rs2_bypass[3] ;
 wire \core_pipeline.decode_to_execute_rs2_bypass[4] ;
 wire \core_pipeline.decode_to_execute_rs2_bypass[5] ;
 wire \core_pipeline.decode_to_execute_rs2_bypass[6] ;
 wire \core_pipeline.decode_to_execute_rs2_bypass[7] ;
 wire \core_pipeline.decode_to_execute_rs2_bypass[8] ;
 wire \core_pipeline.decode_to_execute_rs2_bypass[9] ;
 wire \core_pipeline.decode_to_execute_rs2_bypassed ;
 wire \core_pipeline.decode_to_execute_rs2_data[0] ;
 wire \core_pipeline.decode_to_execute_rs2_data[10] ;
 wire \core_pipeline.decode_to_execute_rs2_data[11] ;
 wire \core_pipeline.decode_to_execute_rs2_data[12] ;
 wire \core_pipeline.decode_to_execute_rs2_data[13] ;
 wire \core_pipeline.decode_to_execute_rs2_data[14] ;
 wire \core_pipeline.decode_to_execute_rs2_data[15] ;
 wire \core_pipeline.decode_to_execute_rs2_data[16] ;
 wire \core_pipeline.decode_to_execute_rs2_data[17] ;
 wire \core_pipeline.decode_to_execute_rs2_data[18] ;
 wire \core_pipeline.decode_to_execute_rs2_data[19] ;
 wire \core_pipeline.decode_to_execute_rs2_data[1] ;
 wire \core_pipeline.decode_to_execute_rs2_data[20] ;
 wire \core_pipeline.decode_to_execute_rs2_data[21] ;
 wire \core_pipeline.decode_to_execute_rs2_data[22] ;
 wire \core_pipeline.decode_to_execute_rs2_data[23] ;
 wire \core_pipeline.decode_to_execute_rs2_data[24] ;
 wire \core_pipeline.decode_to_execute_rs2_data[25] ;
 wire \core_pipeline.decode_to_execute_rs2_data[26] ;
 wire \core_pipeline.decode_to_execute_rs2_data[27] ;
 wire \core_pipeline.decode_to_execute_rs2_data[28] ;
 wire \core_pipeline.decode_to_execute_rs2_data[29] ;
 wire \core_pipeline.decode_to_execute_rs2_data[2] ;
 wire \core_pipeline.decode_to_execute_rs2_data[30] ;
 wire \core_pipeline.decode_to_execute_rs2_data[31] ;
 wire \core_pipeline.decode_to_execute_rs2_data[3] ;
 wire \core_pipeline.decode_to_execute_rs2_data[4] ;
 wire \core_pipeline.decode_to_execute_rs2_data[5] ;
 wire \core_pipeline.decode_to_execute_rs2_data[6] ;
 wire \core_pipeline.decode_to_execute_rs2_data[7] ;
 wire \core_pipeline.decode_to_execute_rs2_data[8] ;
 wire \core_pipeline.decode_to_execute_rs2_data[9] ;
 wire \core_pipeline.decode_to_execute_store ;
 wire \core_pipeline.decode_to_execute_valid ;
 wire \core_pipeline.decode_to_execute_wfi ;
 wire \core_pipeline.decode_to_execute_write_select[0] ;
 wire \core_pipeline.decode_to_execute_write_select[1] ;
 wire \core_pipeline.decode_to_regfile_rs1_address[0] ;
 wire \core_pipeline.decode_to_regfile_rs1_address[1] ;
 wire \core_pipeline.decode_to_regfile_rs1_address[2] ;
 wire \core_pipeline.decode_to_regfile_rs1_address[3] ;
 wire \core_pipeline.decode_to_regfile_rs1_address[4] ;
 wire \core_pipeline.execute_to_memory_branch ;
 wire \core_pipeline.execute_to_memory_bypass_memory ;
 wire \core_pipeline.execute_to_memory_csr_address[0] ;
 wire \core_pipeline.execute_to_memory_csr_address[10] ;
 wire \core_pipeline.execute_to_memory_csr_address[11] ;
 wire \core_pipeline.execute_to_memory_csr_address[1] ;
 wire \core_pipeline.execute_to_memory_csr_address[2] ;
 wire \core_pipeline.execute_to_memory_csr_address[3] ;
 wire \core_pipeline.execute_to_memory_csr_address[4] ;
 wire \core_pipeline.execute_to_memory_csr_address[5] ;
 wire \core_pipeline.execute_to_memory_csr_address[6] ;
 wire \core_pipeline.execute_to_memory_csr_address[7] ;
 wire \core_pipeline.execute_to_memory_csr_address[8] ;
 wire \core_pipeline.execute_to_memory_csr_address[9] ;
 wire \core_pipeline.execute_to_memory_csr_data[0] ;
 wire \core_pipeline.execute_to_memory_csr_data[10] ;
 wire \core_pipeline.execute_to_memory_csr_data[11] ;
 wire \core_pipeline.execute_to_memory_csr_data[12] ;
 wire \core_pipeline.execute_to_memory_csr_data[13] ;
 wire \core_pipeline.execute_to_memory_csr_data[14] ;
 wire \core_pipeline.execute_to_memory_csr_data[15] ;
 wire \core_pipeline.execute_to_memory_csr_data[16] ;
 wire \core_pipeline.execute_to_memory_csr_data[17] ;
 wire \core_pipeline.execute_to_memory_csr_data[18] ;
 wire \core_pipeline.execute_to_memory_csr_data[19] ;
 wire \core_pipeline.execute_to_memory_csr_data[1] ;
 wire \core_pipeline.execute_to_memory_csr_data[20] ;
 wire \core_pipeline.execute_to_memory_csr_data[21] ;
 wire \core_pipeline.execute_to_memory_csr_data[22] ;
 wire \core_pipeline.execute_to_memory_csr_data[23] ;
 wire \core_pipeline.execute_to_memory_csr_data[24] ;
 wire \core_pipeline.execute_to_memory_csr_data[25] ;
 wire \core_pipeline.execute_to_memory_csr_data[26] ;
 wire \core_pipeline.execute_to_memory_csr_data[27] ;
 wire \core_pipeline.execute_to_memory_csr_data[28] ;
 wire \core_pipeline.execute_to_memory_csr_data[29] ;
 wire \core_pipeline.execute_to_memory_csr_data[2] ;
 wire \core_pipeline.execute_to_memory_csr_data[30] ;
 wire \core_pipeline.execute_to_memory_csr_data[31] ;
 wire \core_pipeline.execute_to_memory_csr_data[3] ;
 wire \core_pipeline.execute_to_memory_csr_data[4] ;
 wire \core_pipeline.execute_to_memory_csr_data[5] ;
 wire \core_pipeline.execute_to_memory_csr_data[6] ;
 wire \core_pipeline.execute_to_memory_csr_data[7] ;
 wire \core_pipeline.execute_to_memory_csr_data[8] ;
 wire \core_pipeline.execute_to_memory_csr_data[9] ;
 wire \core_pipeline.execute_to_memory_csr_write ;
 wire \core_pipeline.execute_to_memory_ecause[0] ;
 wire \core_pipeline.execute_to_memory_ecause[1] ;
 wire \core_pipeline.execute_to_memory_ecause[3] ;
 wire \core_pipeline.execute_to_memory_exception ;
 wire \core_pipeline.execute_to_memory_jump ;
 wire \core_pipeline.execute_to_memory_load ;
 wire \core_pipeline.execute_to_memory_mret ;
 wire \core_pipeline.execute_to_memory_next_pc[0] ;
 wire \core_pipeline.execute_to_memory_next_pc[10] ;
 wire \core_pipeline.execute_to_memory_next_pc[11] ;
 wire \core_pipeline.execute_to_memory_next_pc[12] ;
 wire \core_pipeline.execute_to_memory_next_pc[13] ;
 wire \core_pipeline.execute_to_memory_next_pc[14] ;
 wire \core_pipeline.execute_to_memory_next_pc[15] ;
 wire \core_pipeline.execute_to_memory_next_pc[16] ;
 wire \core_pipeline.execute_to_memory_next_pc[17] ;
 wire \core_pipeline.execute_to_memory_next_pc[18] ;
 wire \core_pipeline.execute_to_memory_next_pc[19] ;
 wire \core_pipeline.execute_to_memory_next_pc[1] ;
 wire \core_pipeline.execute_to_memory_next_pc[20] ;
 wire \core_pipeline.execute_to_memory_next_pc[21] ;
 wire \core_pipeline.execute_to_memory_next_pc[22] ;
 wire \core_pipeline.execute_to_memory_next_pc[23] ;
 wire \core_pipeline.execute_to_memory_next_pc[24] ;
 wire \core_pipeline.execute_to_memory_next_pc[25] ;
 wire \core_pipeline.execute_to_memory_next_pc[26] ;
 wire \core_pipeline.execute_to_memory_next_pc[27] ;
 wire \core_pipeline.execute_to_memory_next_pc[28] ;
 wire \core_pipeline.execute_to_memory_next_pc[29] ;
 wire \core_pipeline.execute_to_memory_next_pc[2] ;
 wire \core_pipeline.execute_to_memory_next_pc[30] ;
 wire \core_pipeline.execute_to_memory_next_pc[31] ;
 wire \core_pipeline.execute_to_memory_next_pc[3] ;
 wire \core_pipeline.execute_to_memory_next_pc[4] ;
 wire \core_pipeline.execute_to_memory_next_pc[5] ;
 wire \core_pipeline.execute_to_memory_next_pc[6] ;
 wire \core_pipeline.execute_to_memory_next_pc[7] ;
 wire \core_pipeline.execute_to_memory_next_pc[8] ;
 wire \core_pipeline.execute_to_memory_next_pc[9] ;
 wire \core_pipeline.execute_to_memory_pc[10] ;
 wire \core_pipeline.execute_to_memory_pc[11] ;
 wire \core_pipeline.execute_to_memory_pc[12] ;
 wire \core_pipeline.execute_to_memory_pc[13] ;
 wire \core_pipeline.execute_to_memory_pc[14] ;
 wire \core_pipeline.execute_to_memory_pc[15] ;
 wire \core_pipeline.execute_to_memory_pc[16] ;
 wire \core_pipeline.execute_to_memory_pc[17] ;
 wire \core_pipeline.execute_to_memory_pc[18] ;
 wire \core_pipeline.execute_to_memory_pc[19] ;
 wire \core_pipeline.execute_to_memory_pc[20] ;
 wire \core_pipeline.execute_to_memory_pc[21] ;
 wire \core_pipeline.execute_to_memory_pc[22] ;
 wire \core_pipeline.execute_to_memory_pc[23] ;
 wire \core_pipeline.execute_to_memory_pc[24] ;
 wire \core_pipeline.execute_to_memory_pc[25] ;
 wire \core_pipeline.execute_to_memory_pc[26] ;
 wire \core_pipeline.execute_to_memory_pc[27] ;
 wire \core_pipeline.execute_to_memory_pc[28] ;
 wire \core_pipeline.execute_to_memory_pc[29] ;
 wire \core_pipeline.execute_to_memory_pc[2] ;
 wire \core_pipeline.execute_to_memory_pc[30] ;
 wire \core_pipeline.execute_to_memory_pc[31] ;
 wire \core_pipeline.execute_to_memory_pc[3] ;
 wire \core_pipeline.execute_to_memory_pc[4] ;
 wire \core_pipeline.execute_to_memory_pc[5] ;
 wire \core_pipeline.execute_to_memory_pc[6] ;
 wire \core_pipeline.execute_to_memory_pc[7] ;
 wire \core_pipeline.execute_to_memory_pc[8] ;
 wire \core_pipeline.execute_to_memory_pc[9] ;
 wire \core_pipeline.execute_to_memory_rd_address[0] ;
 wire \core_pipeline.execute_to_memory_rd_address[1] ;
 wire \core_pipeline.execute_to_memory_rd_address[2] ;
 wire \core_pipeline.execute_to_memory_rd_address[3] ;
 wire \core_pipeline.execute_to_memory_rd_address[4] ;
 wire \core_pipeline.execute_to_memory_store ;
 wire \core_pipeline.execute_to_memory_valid ;
 wire \core_pipeline.execute_to_memory_wfi ;
 wire \core_pipeline.execute_to_memory_write_select[0] ;
 wire \core_pipeline.execute_to_memory_write_select[1] ;
 wire \core_pipeline.fetch_to_decode_instruction[0] ;
 wire \core_pipeline.fetch_to_decode_instruction[10] ;
 wire \core_pipeline.fetch_to_decode_instruction[11] ;
 wire \core_pipeline.fetch_to_decode_instruction[12] ;
 wire \core_pipeline.fetch_to_decode_instruction[13] ;
 wire \core_pipeline.fetch_to_decode_instruction[14] ;
 wire \core_pipeline.fetch_to_decode_instruction[1] ;
 wire \core_pipeline.fetch_to_decode_instruction[2] ;
 wire \core_pipeline.fetch_to_decode_instruction[3] ;
 wire \core_pipeline.fetch_to_decode_instruction[4] ;
 wire \core_pipeline.fetch_to_decode_instruction[5] ;
 wire \core_pipeline.fetch_to_decode_instruction[6] ;
 wire \core_pipeline.fetch_to_decode_instruction[7] ;
 wire \core_pipeline.fetch_to_decode_instruction[8] ;
 wire \core_pipeline.fetch_to_decode_instruction[9] ;
 wire \core_pipeline.fetch_to_decode_next_pc[0] ;
 wire \core_pipeline.fetch_to_decode_next_pc[10] ;
 wire \core_pipeline.fetch_to_decode_next_pc[11] ;
 wire \core_pipeline.fetch_to_decode_next_pc[12] ;
 wire \core_pipeline.fetch_to_decode_next_pc[13] ;
 wire \core_pipeline.fetch_to_decode_next_pc[14] ;
 wire \core_pipeline.fetch_to_decode_next_pc[15] ;
 wire \core_pipeline.fetch_to_decode_next_pc[16] ;
 wire \core_pipeline.fetch_to_decode_next_pc[17] ;
 wire \core_pipeline.fetch_to_decode_next_pc[18] ;
 wire \core_pipeline.fetch_to_decode_next_pc[19] ;
 wire \core_pipeline.fetch_to_decode_next_pc[1] ;
 wire \core_pipeline.fetch_to_decode_next_pc[20] ;
 wire \core_pipeline.fetch_to_decode_next_pc[21] ;
 wire \core_pipeline.fetch_to_decode_next_pc[22] ;
 wire \core_pipeline.fetch_to_decode_next_pc[23] ;
 wire \core_pipeline.fetch_to_decode_next_pc[24] ;
 wire \core_pipeline.fetch_to_decode_next_pc[25] ;
 wire \core_pipeline.fetch_to_decode_next_pc[26] ;
 wire \core_pipeline.fetch_to_decode_next_pc[27] ;
 wire \core_pipeline.fetch_to_decode_next_pc[28] ;
 wire \core_pipeline.fetch_to_decode_next_pc[29] ;
 wire \core_pipeline.fetch_to_decode_next_pc[2] ;
 wire \core_pipeline.fetch_to_decode_next_pc[30] ;
 wire \core_pipeline.fetch_to_decode_next_pc[31] ;
 wire \core_pipeline.fetch_to_decode_next_pc[3] ;
 wire \core_pipeline.fetch_to_decode_next_pc[4] ;
 wire \core_pipeline.fetch_to_decode_next_pc[5] ;
 wire \core_pipeline.fetch_to_decode_next_pc[6] ;
 wire \core_pipeline.fetch_to_decode_next_pc[7] ;
 wire \core_pipeline.fetch_to_decode_next_pc[8] ;
 wire \core_pipeline.fetch_to_decode_next_pc[9] ;
 wire \core_pipeline.fetch_to_decode_pc[10] ;
 wire \core_pipeline.fetch_to_decode_pc[11] ;
 wire \core_pipeline.fetch_to_decode_pc[12] ;
 wire \core_pipeline.fetch_to_decode_pc[13] ;
 wire \core_pipeline.fetch_to_decode_pc[14] ;
 wire \core_pipeline.fetch_to_decode_pc[15] ;
 wire \core_pipeline.fetch_to_decode_pc[16] ;
 wire \core_pipeline.fetch_to_decode_pc[17] ;
 wire \core_pipeline.fetch_to_decode_pc[18] ;
 wire \core_pipeline.fetch_to_decode_pc[19] ;
 wire \core_pipeline.fetch_to_decode_pc[20] ;
 wire \core_pipeline.fetch_to_decode_pc[21] ;
 wire \core_pipeline.fetch_to_decode_pc[22] ;
 wire \core_pipeline.fetch_to_decode_pc[23] ;
 wire \core_pipeline.fetch_to_decode_pc[24] ;
 wire \core_pipeline.fetch_to_decode_pc[25] ;
 wire \core_pipeline.fetch_to_decode_pc[26] ;
 wire \core_pipeline.fetch_to_decode_pc[27] ;
 wire \core_pipeline.fetch_to_decode_pc[28] ;
 wire \core_pipeline.fetch_to_decode_pc[29] ;
 wire \core_pipeline.fetch_to_decode_pc[2] ;
 wire \core_pipeline.fetch_to_decode_pc[30] ;
 wire \core_pipeline.fetch_to_decode_pc[31] ;
 wire \core_pipeline.fetch_to_decode_pc[3] ;
 wire \core_pipeline.fetch_to_decode_pc[4] ;
 wire \core_pipeline.fetch_to_decode_pc[5] ;
 wire \core_pipeline.fetch_to_decode_pc[6] ;
 wire \core_pipeline.fetch_to_decode_pc[7] ;
 wire \core_pipeline.fetch_to_decode_pc[8] ;
 wire \core_pipeline.fetch_to_decode_pc[9] ;
 wire \core_pipeline.fetch_to_decode_valid ;
 wire \core_pipeline.memory_to_writeback_alu_data[0] ;
 wire \core_pipeline.memory_to_writeback_alu_data[10] ;
 wire \core_pipeline.memory_to_writeback_alu_data[11] ;
 wire \core_pipeline.memory_to_writeback_alu_data[12] ;
 wire \core_pipeline.memory_to_writeback_alu_data[13] ;
 wire \core_pipeline.memory_to_writeback_alu_data[14] ;
 wire \core_pipeline.memory_to_writeback_alu_data[15] ;
 wire \core_pipeline.memory_to_writeback_alu_data[16] ;
 wire \core_pipeline.memory_to_writeback_alu_data[17] ;
 wire \core_pipeline.memory_to_writeback_alu_data[18] ;
 wire \core_pipeline.memory_to_writeback_alu_data[19] ;
 wire \core_pipeline.memory_to_writeback_alu_data[1] ;
 wire \core_pipeline.memory_to_writeback_alu_data[20] ;
 wire \core_pipeline.memory_to_writeback_alu_data[21] ;
 wire \core_pipeline.memory_to_writeback_alu_data[22] ;
 wire \core_pipeline.memory_to_writeback_alu_data[23] ;
 wire \core_pipeline.memory_to_writeback_alu_data[24] ;
 wire \core_pipeline.memory_to_writeback_alu_data[25] ;
 wire \core_pipeline.memory_to_writeback_alu_data[26] ;
 wire \core_pipeline.memory_to_writeback_alu_data[27] ;
 wire \core_pipeline.memory_to_writeback_alu_data[28] ;
 wire \core_pipeline.memory_to_writeback_alu_data[29] ;
 wire \core_pipeline.memory_to_writeback_alu_data[2] ;
 wire \core_pipeline.memory_to_writeback_alu_data[30] ;
 wire \core_pipeline.memory_to_writeback_alu_data[31] ;
 wire \core_pipeline.memory_to_writeback_alu_data[3] ;
 wire \core_pipeline.memory_to_writeback_alu_data[4] ;
 wire \core_pipeline.memory_to_writeback_alu_data[5] ;
 wire \core_pipeline.memory_to_writeback_alu_data[6] ;
 wire \core_pipeline.memory_to_writeback_alu_data[7] ;
 wire \core_pipeline.memory_to_writeback_alu_data[8] ;
 wire \core_pipeline.memory_to_writeback_alu_data[9] ;
 wire \core_pipeline.memory_to_writeback_csr_address[0] ;
 wire \core_pipeline.memory_to_writeback_csr_address[10] ;
 wire \core_pipeline.memory_to_writeback_csr_address[11] ;
 wire \core_pipeline.memory_to_writeback_csr_address[1] ;
 wire \core_pipeline.memory_to_writeback_csr_address[2] ;
 wire \core_pipeline.memory_to_writeback_csr_address[3] ;
 wire \core_pipeline.memory_to_writeback_csr_address[4] ;
 wire \core_pipeline.memory_to_writeback_csr_address[5] ;
 wire \core_pipeline.memory_to_writeback_csr_address[6] ;
 wire \core_pipeline.memory_to_writeback_csr_address[7] ;
 wire \core_pipeline.memory_to_writeback_csr_address[8] ;
 wire \core_pipeline.memory_to_writeback_csr_address[9] ;
 wire \core_pipeline.memory_to_writeback_csr_data[0] ;
 wire \core_pipeline.memory_to_writeback_csr_data[10] ;
 wire \core_pipeline.memory_to_writeback_csr_data[11] ;
 wire \core_pipeline.memory_to_writeback_csr_data[12] ;
 wire \core_pipeline.memory_to_writeback_csr_data[13] ;
 wire \core_pipeline.memory_to_writeback_csr_data[14] ;
 wire \core_pipeline.memory_to_writeback_csr_data[15] ;
 wire \core_pipeline.memory_to_writeback_csr_data[16] ;
 wire \core_pipeline.memory_to_writeback_csr_data[17] ;
 wire \core_pipeline.memory_to_writeback_csr_data[18] ;
 wire \core_pipeline.memory_to_writeback_csr_data[19] ;
 wire \core_pipeline.memory_to_writeback_csr_data[1] ;
 wire \core_pipeline.memory_to_writeback_csr_data[20] ;
 wire \core_pipeline.memory_to_writeback_csr_data[21] ;
 wire \core_pipeline.memory_to_writeback_csr_data[22] ;
 wire \core_pipeline.memory_to_writeback_csr_data[23] ;
 wire \core_pipeline.memory_to_writeback_csr_data[24] ;
 wire \core_pipeline.memory_to_writeback_csr_data[25] ;
 wire \core_pipeline.memory_to_writeback_csr_data[26] ;
 wire \core_pipeline.memory_to_writeback_csr_data[27] ;
 wire \core_pipeline.memory_to_writeback_csr_data[28] ;
 wire \core_pipeline.memory_to_writeback_csr_data[29] ;
 wire \core_pipeline.memory_to_writeback_csr_data[2] ;
 wire \core_pipeline.memory_to_writeback_csr_data[30] ;
 wire \core_pipeline.memory_to_writeback_csr_data[31] ;
 wire \core_pipeline.memory_to_writeback_csr_data[3] ;
 wire \core_pipeline.memory_to_writeback_csr_data[4] ;
 wire \core_pipeline.memory_to_writeback_csr_data[5] ;
 wire \core_pipeline.memory_to_writeback_csr_data[6] ;
 wire \core_pipeline.memory_to_writeback_csr_data[7] ;
 wire \core_pipeline.memory_to_writeback_csr_data[8] ;
 wire \core_pipeline.memory_to_writeback_csr_data[9] ;
 wire \core_pipeline.memory_to_writeback_csr_write ;
 wire \core_pipeline.memory_to_writeback_ecause[0] ;
 wire \core_pipeline.memory_to_writeback_ecause[1] ;
 wire \core_pipeline.memory_to_writeback_ecause[2] ;
 wire \core_pipeline.memory_to_writeback_ecause[3] ;
 wire \core_pipeline.memory_to_writeback_exception ;
 wire \core_pipeline.memory_to_writeback_load_data[0] ;
 wire \core_pipeline.memory_to_writeback_load_data[10] ;
 wire \core_pipeline.memory_to_writeback_load_data[11] ;
 wire \core_pipeline.memory_to_writeback_load_data[12] ;
 wire \core_pipeline.memory_to_writeback_load_data[13] ;
 wire \core_pipeline.memory_to_writeback_load_data[14] ;
 wire \core_pipeline.memory_to_writeback_load_data[15] ;
 wire \core_pipeline.memory_to_writeback_load_data[16] ;
 wire \core_pipeline.memory_to_writeback_load_data[17] ;
 wire \core_pipeline.memory_to_writeback_load_data[18] ;
 wire \core_pipeline.memory_to_writeback_load_data[19] ;
 wire \core_pipeline.memory_to_writeback_load_data[1] ;
 wire \core_pipeline.memory_to_writeback_load_data[20] ;
 wire \core_pipeline.memory_to_writeback_load_data[21] ;
 wire \core_pipeline.memory_to_writeback_load_data[22] ;
 wire \core_pipeline.memory_to_writeback_load_data[23] ;
 wire \core_pipeline.memory_to_writeback_load_data[24] ;
 wire \core_pipeline.memory_to_writeback_load_data[25] ;
 wire \core_pipeline.memory_to_writeback_load_data[26] ;
 wire \core_pipeline.memory_to_writeback_load_data[27] ;
 wire \core_pipeline.memory_to_writeback_load_data[28] ;
 wire \core_pipeline.memory_to_writeback_load_data[29] ;
 wire \core_pipeline.memory_to_writeback_load_data[2] ;
 wire \core_pipeline.memory_to_writeback_load_data[30] ;
 wire \core_pipeline.memory_to_writeback_load_data[31] ;
 wire \core_pipeline.memory_to_writeback_load_data[3] ;
 wire \core_pipeline.memory_to_writeback_load_data[4] ;
 wire \core_pipeline.memory_to_writeback_load_data[5] ;
 wire \core_pipeline.memory_to_writeback_load_data[6] ;
 wire \core_pipeline.memory_to_writeback_load_data[7] ;
 wire \core_pipeline.memory_to_writeback_load_data[8] ;
 wire \core_pipeline.memory_to_writeback_load_data[9] ;
 wire \core_pipeline.memory_to_writeback_mret ;
 wire \core_pipeline.memory_to_writeback_next_pc[0] ;
 wire \core_pipeline.memory_to_writeback_next_pc[10] ;
 wire \core_pipeline.memory_to_writeback_next_pc[11] ;
 wire \core_pipeline.memory_to_writeback_next_pc[12] ;
 wire \core_pipeline.memory_to_writeback_next_pc[13] ;
 wire \core_pipeline.memory_to_writeback_next_pc[14] ;
 wire \core_pipeline.memory_to_writeback_next_pc[15] ;
 wire \core_pipeline.memory_to_writeback_next_pc[16] ;
 wire \core_pipeline.memory_to_writeback_next_pc[17] ;
 wire \core_pipeline.memory_to_writeback_next_pc[18] ;
 wire \core_pipeline.memory_to_writeback_next_pc[19] ;
 wire \core_pipeline.memory_to_writeback_next_pc[1] ;
 wire \core_pipeline.memory_to_writeback_next_pc[20] ;
 wire \core_pipeline.memory_to_writeback_next_pc[21] ;
 wire \core_pipeline.memory_to_writeback_next_pc[22] ;
 wire \core_pipeline.memory_to_writeback_next_pc[23] ;
 wire \core_pipeline.memory_to_writeback_next_pc[24] ;
 wire \core_pipeline.memory_to_writeback_next_pc[25] ;
 wire \core_pipeline.memory_to_writeback_next_pc[26] ;
 wire \core_pipeline.memory_to_writeback_next_pc[27] ;
 wire \core_pipeline.memory_to_writeback_next_pc[28] ;
 wire \core_pipeline.memory_to_writeback_next_pc[29] ;
 wire \core_pipeline.memory_to_writeback_next_pc[2] ;
 wire \core_pipeline.memory_to_writeback_next_pc[30] ;
 wire \core_pipeline.memory_to_writeback_next_pc[31] ;
 wire \core_pipeline.memory_to_writeback_next_pc[3] ;
 wire \core_pipeline.memory_to_writeback_next_pc[4] ;
 wire \core_pipeline.memory_to_writeback_next_pc[5] ;
 wire \core_pipeline.memory_to_writeback_next_pc[6] ;
 wire \core_pipeline.memory_to_writeback_next_pc[7] ;
 wire \core_pipeline.memory_to_writeback_next_pc[8] ;
 wire \core_pipeline.memory_to_writeback_next_pc[9] ;
 wire \core_pipeline.memory_to_writeback_pc[10] ;
 wire \core_pipeline.memory_to_writeback_pc[11] ;
 wire \core_pipeline.memory_to_writeback_pc[12] ;
 wire \core_pipeline.memory_to_writeback_pc[13] ;
 wire \core_pipeline.memory_to_writeback_pc[14] ;
 wire \core_pipeline.memory_to_writeback_pc[15] ;
 wire \core_pipeline.memory_to_writeback_pc[16] ;
 wire \core_pipeline.memory_to_writeback_pc[17] ;
 wire \core_pipeline.memory_to_writeback_pc[18] ;
 wire \core_pipeline.memory_to_writeback_pc[19] ;
 wire \core_pipeline.memory_to_writeback_pc[20] ;
 wire \core_pipeline.memory_to_writeback_pc[21] ;
 wire \core_pipeline.memory_to_writeback_pc[22] ;
 wire \core_pipeline.memory_to_writeback_pc[23] ;
 wire \core_pipeline.memory_to_writeback_pc[24] ;
 wire \core_pipeline.memory_to_writeback_pc[25] ;
 wire \core_pipeline.memory_to_writeback_pc[26] ;
 wire \core_pipeline.memory_to_writeback_pc[27] ;
 wire \core_pipeline.memory_to_writeback_pc[28] ;
 wire \core_pipeline.memory_to_writeback_pc[29] ;
 wire \core_pipeline.memory_to_writeback_pc[2] ;
 wire \core_pipeline.memory_to_writeback_pc[30] ;
 wire \core_pipeline.memory_to_writeback_pc[31] ;
 wire \core_pipeline.memory_to_writeback_pc[3] ;
 wire \core_pipeline.memory_to_writeback_pc[4] ;
 wire \core_pipeline.memory_to_writeback_pc[5] ;
 wire \core_pipeline.memory_to_writeback_pc[6] ;
 wire \core_pipeline.memory_to_writeback_pc[7] ;
 wire \core_pipeline.memory_to_writeback_pc[8] ;
 wire \core_pipeline.memory_to_writeback_pc[9] ;
 wire \core_pipeline.memory_to_writeback_rd_address[0] ;
 wire \core_pipeline.memory_to_writeback_rd_address[1] ;
 wire \core_pipeline.memory_to_writeback_rd_address[2] ;
 wire \core_pipeline.memory_to_writeback_rd_address[3] ;
 wire \core_pipeline.memory_to_writeback_rd_address[4] ;
 wire \core_pipeline.memory_to_writeback_valid ;
 wire \core_pipeline.memory_to_writeback_wfi ;
 wire \core_pipeline.memory_to_writeback_write_select[0] ;
 wire \core_pipeline.memory_to_writeback_write_select[1] ;
 wire \core_pipeline.pipeline_csr.cycle[0] ;
 wire \core_pipeline.pipeline_csr.cycle[10] ;
 wire \core_pipeline.pipeline_csr.cycle[11] ;
 wire \core_pipeline.pipeline_csr.cycle[12] ;
 wire \core_pipeline.pipeline_csr.cycle[13] ;
 wire \core_pipeline.pipeline_csr.cycle[14] ;
 wire \core_pipeline.pipeline_csr.cycle[15] ;
 wire \core_pipeline.pipeline_csr.cycle[16] ;
 wire \core_pipeline.pipeline_csr.cycle[17] ;
 wire \core_pipeline.pipeline_csr.cycle[18] ;
 wire \core_pipeline.pipeline_csr.cycle[19] ;
 wire \core_pipeline.pipeline_csr.cycle[1] ;
 wire \core_pipeline.pipeline_csr.cycle[20] ;
 wire \core_pipeline.pipeline_csr.cycle[21] ;
 wire \core_pipeline.pipeline_csr.cycle[22] ;
 wire \core_pipeline.pipeline_csr.cycle[23] ;
 wire \core_pipeline.pipeline_csr.cycle[24] ;
 wire \core_pipeline.pipeline_csr.cycle[25] ;
 wire \core_pipeline.pipeline_csr.cycle[26] ;
 wire \core_pipeline.pipeline_csr.cycle[27] ;
 wire \core_pipeline.pipeline_csr.cycle[28] ;
 wire \core_pipeline.pipeline_csr.cycle[29] ;
 wire \core_pipeline.pipeline_csr.cycle[2] ;
 wire \core_pipeline.pipeline_csr.cycle[30] ;
 wire \core_pipeline.pipeline_csr.cycle[31] ;
 wire \core_pipeline.pipeline_csr.cycle[32] ;
 wire \core_pipeline.pipeline_csr.cycle[33] ;
 wire \core_pipeline.pipeline_csr.cycle[34] ;
 wire \core_pipeline.pipeline_csr.cycle[35] ;
 wire \core_pipeline.pipeline_csr.cycle[36] ;
 wire \core_pipeline.pipeline_csr.cycle[37] ;
 wire \core_pipeline.pipeline_csr.cycle[38] ;
 wire \core_pipeline.pipeline_csr.cycle[39] ;
 wire \core_pipeline.pipeline_csr.cycle[3] ;
 wire \core_pipeline.pipeline_csr.cycle[40] ;
 wire \core_pipeline.pipeline_csr.cycle[41] ;
 wire \core_pipeline.pipeline_csr.cycle[42] ;
 wire \core_pipeline.pipeline_csr.cycle[43] ;
 wire \core_pipeline.pipeline_csr.cycle[44] ;
 wire \core_pipeline.pipeline_csr.cycle[45] ;
 wire \core_pipeline.pipeline_csr.cycle[46] ;
 wire \core_pipeline.pipeline_csr.cycle[47] ;
 wire \core_pipeline.pipeline_csr.cycle[48] ;
 wire \core_pipeline.pipeline_csr.cycle[49] ;
 wire \core_pipeline.pipeline_csr.cycle[4] ;
 wire \core_pipeline.pipeline_csr.cycle[50] ;
 wire \core_pipeline.pipeline_csr.cycle[51] ;
 wire \core_pipeline.pipeline_csr.cycle[52] ;
 wire \core_pipeline.pipeline_csr.cycle[53] ;
 wire \core_pipeline.pipeline_csr.cycle[54] ;
 wire \core_pipeline.pipeline_csr.cycle[55] ;
 wire \core_pipeline.pipeline_csr.cycle[56] ;
 wire \core_pipeline.pipeline_csr.cycle[57] ;
 wire \core_pipeline.pipeline_csr.cycle[58] ;
 wire \core_pipeline.pipeline_csr.cycle[59] ;
 wire \core_pipeline.pipeline_csr.cycle[5] ;
 wire \core_pipeline.pipeline_csr.cycle[60] ;
 wire \core_pipeline.pipeline_csr.cycle[61] ;
 wire \core_pipeline.pipeline_csr.cycle[62] ;
 wire \core_pipeline.pipeline_csr.cycle[63] ;
 wire \core_pipeline.pipeline_csr.cycle[6] ;
 wire \core_pipeline.pipeline_csr.cycle[7] ;
 wire \core_pipeline.pipeline_csr.cycle[8] ;
 wire \core_pipeline.pipeline_csr.cycle[9] ;
 wire \core_pipeline.pipeline_csr.ie ;
 wire \core_pipeline.pipeline_csr.instret[0] ;
 wire \core_pipeline.pipeline_csr.instret[10] ;
 wire \core_pipeline.pipeline_csr.instret[11] ;
 wire \core_pipeline.pipeline_csr.instret[12] ;
 wire \core_pipeline.pipeline_csr.instret[13] ;
 wire \core_pipeline.pipeline_csr.instret[14] ;
 wire \core_pipeline.pipeline_csr.instret[15] ;
 wire \core_pipeline.pipeline_csr.instret[16] ;
 wire \core_pipeline.pipeline_csr.instret[17] ;
 wire \core_pipeline.pipeline_csr.instret[18] ;
 wire \core_pipeline.pipeline_csr.instret[19] ;
 wire \core_pipeline.pipeline_csr.instret[1] ;
 wire \core_pipeline.pipeline_csr.instret[20] ;
 wire \core_pipeline.pipeline_csr.instret[21] ;
 wire \core_pipeline.pipeline_csr.instret[22] ;
 wire \core_pipeline.pipeline_csr.instret[23] ;
 wire \core_pipeline.pipeline_csr.instret[24] ;
 wire \core_pipeline.pipeline_csr.instret[25] ;
 wire \core_pipeline.pipeline_csr.instret[26] ;
 wire \core_pipeline.pipeline_csr.instret[27] ;
 wire \core_pipeline.pipeline_csr.instret[28] ;
 wire \core_pipeline.pipeline_csr.instret[29] ;
 wire \core_pipeline.pipeline_csr.instret[2] ;
 wire \core_pipeline.pipeline_csr.instret[30] ;
 wire \core_pipeline.pipeline_csr.instret[31] ;
 wire \core_pipeline.pipeline_csr.instret[32] ;
 wire \core_pipeline.pipeline_csr.instret[33] ;
 wire \core_pipeline.pipeline_csr.instret[34] ;
 wire \core_pipeline.pipeline_csr.instret[35] ;
 wire \core_pipeline.pipeline_csr.instret[36] ;
 wire \core_pipeline.pipeline_csr.instret[37] ;
 wire \core_pipeline.pipeline_csr.instret[38] ;
 wire \core_pipeline.pipeline_csr.instret[39] ;
 wire \core_pipeline.pipeline_csr.instret[3] ;
 wire \core_pipeline.pipeline_csr.instret[40] ;
 wire \core_pipeline.pipeline_csr.instret[41] ;
 wire \core_pipeline.pipeline_csr.instret[42] ;
 wire \core_pipeline.pipeline_csr.instret[43] ;
 wire \core_pipeline.pipeline_csr.instret[44] ;
 wire \core_pipeline.pipeline_csr.instret[45] ;
 wire \core_pipeline.pipeline_csr.instret[46] ;
 wire \core_pipeline.pipeline_csr.instret[47] ;
 wire \core_pipeline.pipeline_csr.instret[48] ;
 wire \core_pipeline.pipeline_csr.instret[49] ;
 wire \core_pipeline.pipeline_csr.instret[4] ;
 wire \core_pipeline.pipeline_csr.instret[50] ;
 wire \core_pipeline.pipeline_csr.instret[51] ;
 wire \core_pipeline.pipeline_csr.instret[52] ;
 wire \core_pipeline.pipeline_csr.instret[53] ;
 wire \core_pipeline.pipeline_csr.instret[54] ;
 wire \core_pipeline.pipeline_csr.instret[55] ;
 wire \core_pipeline.pipeline_csr.instret[56] ;
 wire \core_pipeline.pipeline_csr.instret[57] ;
 wire \core_pipeline.pipeline_csr.instret[58] ;
 wire \core_pipeline.pipeline_csr.instret[59] ;
 wire \core_pipeline.pipeline_csr.instret[5] ;
 wire \core_pipeline.pipeline_csr.instret[60] ;
 wire \core_pipeline.pipeline_csr.instret[61] ;
 wire \core_pipeline.pipeline_csr.instret[62] ;
 wire \core_pipeline.pipeline_csr.instret[63] ;
 wire \core_pipeline.pipeline_csr.instret[6] ;
 wire \core_pipeline.pipeline_csr.instret[7] ;
 wire \core_pipeline.pipeline_csr.instret[8] ;
 wire \core_pipeline.pipeline_csr.instret[9] ;
 wire \core_pipeline.pipeline_csr.mcause[0] ;
 wire \core_pipeline.pipeline_csr.mcause[1] ;
 wire \core_pipeline.pipeline_csr.mcause[2] ;
 wire \core_pipeline.pipeline_csr.mcause[3] ;
 wire \core_pipeline.pipeline_csr.meie ;
 wire \core_pipeline.pipeline_csr.minterupt ;
 wire \core_pipeline.pipeline_csr.mscratch[0] ;
 wire \core_pipeline.pipeline_csr.mscratch[10] ;
 wire \core_pipeline.pipeline_csr.mscratch[11] ;
 wire \core_pipeline.pipeline_csr.mscratch[12] ;
 wire \core_pipeline.pipeline_csr.mscratch[13] ;
 wire \core_pipeline.pipeline_csr.mscratch[14] ;
 wire \core_pipeline.pipeline_csr.mscratch[15] ;
 wire \core_pipeline.pipeline_csr.mscratch[16] ;
 wire \core_pipeline.pipeline_csr.mscratch[17] ;
 wire \core_pipeline.pipeline_csr.mscratch[18] ;
 wire \core_pipeline.pipeline_csr.mscratch[19] ;
 wire \core_pipeline.pipeline_csr.mscratch[1] ;
 wire \core_pipeline.pipeline_csr.mscratch[20] ;
 wire \core_pipeline.pipeline_csr.mscratch[21] ;
 wire \core_pipeline.pipeline_csr.mscratch[22] ;
 wire \core_pipeline.pipeline_csr.mscratch[23] ;
 wire \core_pipeline.pipeline_csr.mscratch[24] ;
 wire \core_pipeline.pipeline_csr.mscratch[25] ;
 wire \core_pipeline.pipeline_csr.mscratch[26] ;
 wire \core_pipeline.pipeline_csr.mscratch[27] ;
 wire \core_pipeline.pipeline_csr.mscratch[28] ;
 wire \core_pipeline.pipeline_csr.mscratch[29] ;
 wire \core_pipeline.pipeline_csr.mscratch[2] ;
 wire \core_pipeline.pipeline_csr.mscratch[30] ;
 wire \core_pipeline.pipeline_csr.mscratch[31] ;
 wire \core_pipeline.pipeline_csr.mscratch[3] ;
 wire \core_pipeline.pipeline_csr.mscratch[4] ;
 wire \core_pipeline.pipeline_csr.mscratch[5] ;
 wire \core_pipeline.pipeline_csr.mscratch[6] ;
 wire \core_pipeline.pipeline_csr.mscratch[7] ;
 wire \core_pipeline.pipeline_csr.mscratch[8] ;
 wire \core_pipeline.pipeline_csr.mscratch[9] ;
 wire \core_pipeline.pipeline_csr.msie ;
 wire \core_pipeline.pipeline_csr.msip ;
 wire \core_pipeline.pipeline_csr.mtie ;
 wire \core_pipeline.pipeline_csr.mtimecmp[0] ;
 wire \core_pipeline.pipeline_csr.mtimecmp[10] ;
 wire \core_pipeline.pipeline_csr.mtimecmp[11] ;
 wire \core_pipeline.pipeline_csr.mtimecmp[12] ;
 wire \core_pipeline.pipeline_csr.mtimecmp[13] ;
 wire \core_pipeline.pipeline_csr.mtimecmp[14] ;
 wire \core_pipeline.pipeline_csr.mtimecmp[15] ;
 wire \core_pipeline.pipeline_csr.mtimecmp[16] ;
 wire \core_pipeline.pipeline_csr.mtimecmp[17] ;
 wire \core_pipeline.pipeline_csr.mtimecmp[18] ;
 wire \core_pipeline.pipeline_csr.mtimecmp[19] ;
 wire \core_pipeline.pipeline_csr.mtimecmp[1] ;
 wire \core_pipeline.pipeline_csr.mtimecmp[20] ;
 wire \core_pipeline.pipeline_csr.mtimecmp[21] ;
 wire \core_pipeline.pipeline_csr.mtimecmp[22] ;
 wire \core_pipeline.pipeline_csr.mtimecmp[23] ;
 wire \core_pipeline.pipeline_csr.mtimecmp[24] ;
 wire \core_pipeline.pipeline_csr.mtimecmp[25] ;
 wire \core_pipeline.pipeline_csr.mtimecmp[26] ;
 wire \core_pipeline.pipeline_csr.mtimecmp[27] ;
 wire \core_pipeline.pipeline_csr.mtimecmp[28] ;
 wire \core_pipeline.pipeline_csr.mtimecmp[29] ;
 wire \core_pipeline.pipeline_csr.mtimecmp[2] ;
 wire \core_pipeline.pipeline_csr.mtimecmp[30] ;
 wire \core_pipeline.pipeline_csr.mtimecmp[31] ;
 wire \core_pipeline.pipeline_csr.mtimecmp[32] ;
 wire \core_pipeline.pipeline_csr.mtimecmp[33] ;
 wire \core_pipeline.pipeline_csr.mtimecmp[34] ;
 wire \core_pipeline.pipeline_csr.mtimecmp[35] ;
 wire \core_pipeline.pipeline_csr.mtimecmp[36] ;
 wire \core_pipeline.pipeline_csr.mtimecmp[37] ;
 wire \core_pipeline.pipeline_csr.mtimecmp[38] ;
 wire \core_pipeline.pipeline_csr.mtimecmp[39] ;
 wire \core_pipeline.pipeline_csr.mtimecmp[3] ;
 wire \core_pipeline.pipeline_csr.mtimecmp[40] ;
 wire \core_pipeline.pipeline_csr.mtimecmp[41] ;
 wire \core_pipeline.pipeline_csr.mtimecmp[42] ;
 wire \core_pipeline.pipeline_csr.mtimecmp[43] ;
 wire \core_pipeline.pipeline_csr.mtimecmp[44] ;
 wire \core_pipeline.pipeline_csr.mtimecmp[45] ;
 wire \core_pipeline.pipeline_csr.mtimecmp[46] ;
 wire \core_pipeline.pipeline_csr.mtimecmp[47] ;
 wire \core_pipeline.pipeline_csr.mtimecmp[48] ;
 wire \core_pipeline.pipeline_csr.mtimecmp[49] ;
 wire \core_pipeline.pipeline_csr.mtimecmp[4] ;
 wire \core_pipeline.pipeline_csr.mtimecmp[50] ;
 wire \core_pipeline.pipeline_csr.mtimecmp[51] ;
 wire \core_pipeline.pipeline_csr.mtimecmp[52] ;
 wire \core_pipeline.pipeline_csr.mtimecmp[53] ;
 wire \core_pipeline.pipeline_csr.mtimecmp[54] ;
 wire \core_pipeline.pipeline_csr.mtimecmp[55] ;
 wire \core_pipeline.pipeline_csr.mtimecmp[56] ;
 wire \core_pipeline.pipeline_csr.mtimecmp[57] ;
 wire \core_pipeline.pipeline_csr.mtimecmp[58] ;
 wire \core_pipeline.pipeline_csr.mtimecmp[59] ;
 wire \core_pipeline.pipeline_csr.mtimecmp[5] ;
 wire \core_pipeline.pipeline_csr.mtimecmp[60] ;
 wire \core_pipeline.pipeline_csr.mtimecmp[61] ;
 wire \core_pipeline.pipeline_csr.mtimecmp[62] ;
 wire \core_pipeline.pipeline_csr.mtimecmp[63] ;
 wire \core_pipeline.pipeline_csr.mtimecmp[6] ;
 wire \core_pipeline.pipeline_csr.mtimecmp[7] ;
 wire \core_pipeline.pipeline_csr.mtimecmp[8] ;
 wire \core_pipeline.pipeline_csr.mtimecmp[9] ;
 wire \core_pipeline.pipeline_csr.mtip ;
 wire \core_pipeline.pipeline_csr.pie ;
 wire \core_pipeline.pipeline_decode.alu_select_a_out[1] ;
 wire \core_pipeline.pipeline_decode.alu_select_a_out[2] ;
 wire \core_pipeline.pipeline_decode.alu_select_b_out[1] ;
 wire \core_pipeline.pipeline_decode.alu_select_b_out[2] ;
 wire \core_pipeline.pipeline_execute.ex_alu.old_function[0] ;
 wire \core_pipeline.pipeline_execute.ex_alu.old_function[1] ;
 wire \core_pipeline.pipeline_execute.ex_alu.old_function[2] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_and_clr[0] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_and_clr[10] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_and_clr[11] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_and_clr[12] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_and_clr[13] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_and_clr[14] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_and_clr[15] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_and_clr[16] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_and_clr[17] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_and_clr[18] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_and_clr[19] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_and_clr[1] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_and_clr[20] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_and_clr[21] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_and_clr[22] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_and_clr[23] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_and_clr[24] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_and_clr[25] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_and_clr[26] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_and_clr[27] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_and_clr[28] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_and_clr[29] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_and_clr[2] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_and_clr[30] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_and_clr[31] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_and_clr[3] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_and_clr[4] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_and_clr[5] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_and_clr[6] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_and_clr[7] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_and_clr[8] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_and_clr[9] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_or[0] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_or[10] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_or[11] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_or[12] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_or[13] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_or[14] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_or[15] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_or[16] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_or[17] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_or[18] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_or[19] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_or[1] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_or[20] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_or[21] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_or[22] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_or[23] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_or[24] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_or[25] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_or[26] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_or[27] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_or[28] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_or[29] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_or[2] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_or[30] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_or[31] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_or[3] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_or[4] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_or[5] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_or[6] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_or[7] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_or[8] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_or[9] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_sll[0] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_sll[10] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_sll[11] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_sll[12] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_sll[13] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_sll[14] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_sll[15] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_sll[16] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_sll[17] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_sll[18] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_sll[19] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_sll[1] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_sll[20] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_sll[21] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_sll[22] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_sll[23] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_sll[24] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_sll[25] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_sll[26] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_sll[27] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_sll[28] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_sll[29] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_sll[2] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_sll[30] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_sll[31] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_sll[3] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_sll[4] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_sll[5] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_sll[6] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_sll[7] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_sll[8] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_sll[9] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_slt[0] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_sltu[0] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_srl_sra[0] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_srl_sra[10] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_srl_sra[11] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_srl_sra[12] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_srl_sra[13] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_srl_sra[14] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_srl_sra[15] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_srl_sra[16] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_srl_sra[17] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_srl_sra[18] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_srl_sra[19] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_srl_sra[1] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_srl_sra[20] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_srl_sra[21] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_srl_sra[22] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_srl_sra[23] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_srl_sra[24] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_srl_sra[25] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_srl_sra[26] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_srl_sra[27] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_srl_sra[28] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_srl_sra[29] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_srl_sra[2] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_srl_sra[30] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_srl_sra[31] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_srl_sra[3] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_srl_sra[4] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_srl_sra[5] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_srl_sra[6] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_srl_sra[7] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_srl_sra[8] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_srl_sra[9] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_xor[0] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_xor[10] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_xor[11] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_xor[12] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_xor[13] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_xor[14] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_xor[15] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_xor[16] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_xor[17] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_xor[18] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_xor[19] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_xor[1] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_xor[20] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_xor[21] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_xor[22] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_xor[23] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_xor[24] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_xor[25] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_xor[26] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_xor[27] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_xor[28] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_xor[29] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_xor[2] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_xor[30] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_xor[31] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_xor[3] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_xor[4] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_xor[5] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_xor[6] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_xor[7] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_xor[8] ;
 wire \core_pipeline.pipeline_execute.ex_alu.result_xor[9] ;
 wire \core_pipeline.pipeline_execute.ex_cmp.negate ;
 wire \core_pipeline.pipeline_execute.ex_cmp.quasi_result ;
 wire \core_pipeline.pipeline_fetch.pc[0] ;
 wire \core_pipeline.pipeline_fetch.pc[10] ;
 wire \core_pipeline.pipeline_fetch.pc[11] ;
 wire \core_pipeline.pipeline_fetch.pc[12] ;
 wire \core_pipeline.pipeline_fetch.pc[13] ;
 wire \core_pipeline.pipeline_fetch.pc[14] ;
 wire \core_pipeline.pipeline_fetch.pc[15] ;
 wire \core_pipeline.pipeline_fetch.pc[16] ;
 wire \core_pipeline.pipeline_fetch.pc[17] ;
 wire \core_pipeline.pipeline_fetch.pc[18] ;
 wire \core_pipeline.pipeline_fetch.pc[19] ;
 wire \core_pipeline.pipeline_fetch.pc[1] ;
 wire \core_pipeline.pipeline_fetch.pc[20] ;
 wire \core_pipeline.pipeline_fetch.pc[21] ;
 wire \core_pipeline.pipeline_fetch.pc[22] ;
 wire \core_pipeline.pipeline_fetch.pc[23] ;
 wire \core_pipeline.pipeline_fetch.pc[24] ;
 wire \core_pipeline.pipeline_fetch.pc[25] ;
 wire \core_pipeline.pipeline_fetch.pc[26] ;
 wire \core_pipeline.pipeline_fetch.pc[27] ;
 wire \core_pipeline.pipeline_fetch.pc[28] ;
 wire \core_pipeline.pipeline_fetch.pc[29] ;
 wire \core_pipeline.pipeline_fetch.pc[2] ;
 wire \core_pipeline.pipeline_fetch.pc[30] ;
 wire \core_pipeline.pipeline_fetch.pc[31] ;
 wire \core_pipeline.pipeline_fetch.pc[3] ;
 wire \core_pipeline.pipeline_fetch.pc[4] ;
 wire \core_pipeline.pipeline_fetch.pc[5] ;
 wire \core_pipeline.pipeline_fetch.pc[6] ;
 wire \core_pipeline.pipeline_fetch.pc[7] ;
 wire \core_pipeline.pipeline_fetch.pc[8] ;
 wire \core_pipeline.pipeline_fetch.pc[9] ;
 wire \core_pipeline.pipeline_registers.registers[0][0] ;
 wire \core_pipeline.pipeline_registers.registers[0][10] ;
 wire \core_pipeline.pipeline_registers.registers[0][11] ;
 wire \core_pipeline.pipeline_registers.registers[0][12] ;
 wire \core_pipeline.pipeline_registers.registers[0][13] ;
 wire \core_pipeline.pipeline_registers.registers[0][14] ;
 wire \core_pipeline.pipeline_registers.registers[0][15] ;
 wire \core_pipeline.pipeline_registers.registers[0][16] ;
 wire \core_pipeline.pipeline_registers.registers[0][17] ;
 wire \core_pipeline.pipeline_registers.registers[0][18] ;
 wire \core_pipeline.pipeline_registers.registers[0][19] ;
 wire \core_pipeline.pipeline_registers.registers[0][1] ;
 wire \core_pipeline.pipeline_registers.registers[0][20] ;
 wire \core_pipeline.pipeline_registers.registers[0][21] ;
 wire \core_pipeline.pipeline_registers.registers[0][22] ;
 wire \core_pipeline.pipeline_registers.registers[0][23] ;
 wire \core_pipeline.pipeline_registers.registers[0][24] ;
 wire \core_pipeline.pipeline_registers.registers[0][25] ;
 wire \core_pipeline.pipeline_registers.registers[0][26] ;
 wire \core_pipeline.pipeline_registers.registers[0][27] ;
 wire \core_pipeline.pipeline_registers.registers[0][28] ;
 wire \core_pipeline.pipeline_registers.registers[0][29] ;
 wire \core_pipeline.pipeline_registers.registers[0][2] ;
 wire \core_pipeline.pipeline_registers.registers[0][30] ;
 wire \core_pipeline.pipeline_registers.registers[0][31] ;
 wire \core_pipeline.pipeline_registers.registers[0][3] ;
 wire \core_pipeline.pipeline_registers.registers[0][4] ;
 wire \core_pipeline.pipeline_registers.registers[0][5] ;
 wire \core_pipeline.pipeline_registers.registers[0][6] ;
 wire \core_pipeline.pipeline_registers.registers[0][7] ;
 wire \core_pipeline.pipeline_registers.registers[0][8] ;
 wire \core_pipeline.pipeline_registers.registers[0][9] ;
 wire \core_pipeline.pipeline_registers.registers[10][0] ;
 wire \core_pipeline.pipeline_registers.registers[10][10] ;
 wire \core_pipeline.pipeline_registers.registers[10][11] ;
 wire \core_pipeline.pipeline_registers.registers[10][12] ;
 wire \core_pipeline.pipeline_registers.registers[10][13] ;
 wire \core_pipeline.pipeline_registers.registers[10][14] ;
 wire \core_pipeline.pipeline_registers.registers[10][15] ;
 wire \core_pipeline.pipeline_registers.registers[10][16] ;
 wire \core_pipeline.pipeline_registers.registers[10][17] ;
 wire \core_pipeline.pipeline_registers.registers[10][18] ;
 wire \core_pipeline.pipeline_registers.registers[10][19] ;
 wire \core_pipeline.pipeline_registers.registers[10][1] ;
 wire \core_pipeline.pipeline_registers.registers[10][20] ;
 wire \core_pipeline.pipeline_registers.registers[10][21] ;
 wire \core_pipeline.pipeline_registers.registers[10][22] ;
 wire \core_pipeline.pipeline_registers.registers[10][23] ;
 wire \core_pipeline.pipeline_registers.registers[10][24] ;
 wire \core_pipeline.pipeline_registers.registers[10][25] ;
 wire \core_pipeline.pipeline_registers.registers[10][26] ;
 wire \core_pipeline.pipeline_registers.registers[10][27] ;
 wire \core_pipeline.pipeline_registers.registers[10][28] ;
 wire \core_pipeline.pipeline_registers.registers[10][29] ;
 wire \core_pipeline.pipeline_registers.registers[10][2] ;
 wire \core_pipeline.pipeline_registers.registers[10][30] ;
 wire \core_pipeline.pipeline_registers.registers[10][31] ;
 wire \core_pipeline.pipeline_registers.registers[10][3] ;
 wire \core_pipeline.pipeline_registers.registers[10][4] ;
 wire \core_pipeline.pipeline_registers.registers[10][5] ;
 wire \core_pipeline.pipeline_registers.registers[10][6] ;
 wire \core_pipeline.pipeline_registers.registers[10][7] ;
 wire \core_pipeline.pipeline_registers.registers[10][8] ;
 wire \core_pipeline.pipeline_registers.registers[10][9] ;
 wire \core_pipeline.pipeline_registers.registers[11][0] ;
 wire \core_pipeline.pipeline_registers.registers[11][10] ;
 wire \core_pipeline.pipeline_registers.registers[11][11] ;
 wire \core_pipeline.pipeline_registers.registers[11][12] ;
 wire \core_pipeline.pipeline_registers.registers[11][13] ;
 wire \core_pipeline.pipeline_registers.registers[11][14] ;
 wire \core_pipeline.pipeline_registers.registers[11][15] ;
 wire \core_pipeline.pipeline_registers.registers[11][16] ;
 wire \core_pipeline.pipeline_registers.registers[11][17] ;
 wire \core_pipeline.pipeline_registers.registers[11][18] ;
 wire \core_pipeline.pipeline_registers.registers[11][19] ;
 wire \core_pipeline.pipeline_registers.registers[11][1] ;
 wire \core_pipeline.pipeline_registers.registers[11][20] ;
 wire \core_pipeline.pipeline_registers.registers[11][21] ;
 wire \core_pipeline.pipeline_registers.registers[11][22] ;
 wire \core_pipeline.pipeline_registers.registers[11][23] ;
 wire \core_pipeline.pipeline_registers.registers[11][24] ;
 wire \core_pipeline.pipeline_registers.registers[11][25] ;
 wire \core_pipeline.pipeline_registers.registers[11][26] ;
 wire \core_pipeline.pipeline_registers.registers[11][27] ;
 wire \core_pipeline.pipeline_registers.registers[11][28] ;
 wire \core_pipeline.pipeline_registers.registers[11][29] ;
 wire \core_pipeline.pipeline_registers.registers[11][2] ;
 wire \core_pipeline.pipeline_registers.registers[11][30] ;
 wire \core_pipeline.pipeline_registers.registers[11][31] ;
 wire \core_pipeline.pipeline_registers.registers[11][3] ;
 wire \core_pipeline.pipeline_registers.registers[11][4] ;
 wire \core_pipeline.pipeline_registers.registers[11][5] ;
 wire \core_pipeline.pipeline_registers.registers[11][6] ;
 wire \core_pipeline.pipeline_registers.registers[11][7] ;
 wire \core_pipeline.pipeline_registers.registers[11][8] ;
 wire \core_pipeline.pipeline_registers.registers[11][9] ;
 wire \core_pipeline.pipeline_registers.registers[12][0] ;
 wire \core_pipeline.pipeline_registers.registers[12][10] ;
 wire \core_pipeline.pipeline_registers.registers[12][11] ;
 wire \core_pipeline.pipeline_registers.registers[12][12] ;
 wire \core_pipeline.pipeline_registers.registers[12][13] ;
 wire \core_pipeline.pipeline_registers.registers[12][14] ;
 wire \core_pipeline.pipeline_registers.registers[12][15] ;
 wire \core_pipeline.pipeline_registers.registers[12][16] ;
 wire \core_pipeline.pipeline_registers.registers[12][17] ;
 wire \core_pipeline.pipeline_registers.registers[12][18] ;
 wire \core_pipeline.pipeline_registers.registers[12][19] ;
 wire \core_pipeline.pipeline_registers.registers[12][1] ;
 wire \core_pipeline.pipeline_registers.registers[12][20] ;
 wire \core_pipeline.pipeline_registers.registers[12][21] ;
 wire \core_pipeline.pipeline_registers.registers[12][22] ;
 wire \core_pipeline.pipeline_registers.registers[12][23] ;
 wire \core_pipeline.pipeline_registers.registers[12][24] ;
 wire \core_pipeline.pipeline_registers.registers[12][25] ;
 wire \core_pipeline.pipeline_registers.registers[12][26] ;
 wire \core_pipeline.pipeline_registers.registers[12][27] ;
 wire \core_pipeline.pipeline_registers.registers[12][28] ;
 wire \core_pipeline.pipeline_registers.registers[12][29] ;
 wire \core_pipeline.pipeline_registers.registers[12][2] ;
 wire \core_pipeline.pipeline_registers.registers[12][30] ;
 wire \core_pipeline.pipeline_registers.registers[12][31] ;
 wire \core_pipeline.pipeline_registers.registers[12][3] ;
 wire \core_pipeline.pipeline_registers.registers[12][4] ;
 wire \core_pipeline.pipeline_registers.registers[12][5] ;
 wire \core_pipeline.pipeline_registers.registers[12][6] ;
 wire \core_pipeline.pipeline_registers.registers[12][7] ;
 wire \core_pipeline.pipeline_registers.registers[12][8] ;
 wire \core_pipeline.pipeline_registers.registers[12][9] ;
 wire \core_pipeline.pipeline_registers.registers[13][0] ;
 wire \core_pipeline.pipeline_registers.registers[13][10] ;
 wire \core_pipeline.pipeline_registers.registers[13][11] ;
 wire \core_pipeline.pipeline_registers.registers[13][12] ;
 wire \core_pipeline.pipeline_registers.registers[13][13] ;
 wire \core_pipeline.pipeline_registers.registers[13][14] ;
 wire \core_pipeline.pipeline_registers.registers[13][15] ;
 wire \core_pipeline.pipeline_registers.registers[13][16] ;
 wire \core_pipeline.pipeline_registers.registers[13][17] ;
 wire \core_pipeline.pipeline_registers.registers[13][18] ;
 wire \core_pipeline.pipeline_registers.registers[13][19] ;
 wire \core_pipeline.pipeline_registers.registers[13][1] ;
 wire \core_pipeline.pipeline_registers.registers[13][20] ;
 wire \core_pipeline.pipeline_registers.registers[13][21] ;
 wire \core_pipeline.pipeline_registers.registers[13][22] ;
 wire \core_pipeline.pipeline_registers.registers[13][23] ;
 wire \core_pipeline.pipeline_registers.registers[13][24] ;
 wire \core_pipeline.pipeline_registers.registers[13][25] ;
 wire \core_pipeline.pipeline_registers.registers[13][26] ;
 wire \core_pipeline.pipeline_registers.registers[13][27] ;
 wire \core_pipeline.pipeline_registers.registers[13][28] ;
 wire \core_pipeline.pipeline_registers.registers[13][29] ;
 wire \core_pipeline.pipeline_registers.registers[13][2] ;
 wire \core_pipeline.pipeline_registers.registers[13][30] ;
 wire \core_pipeline.pipeline_registers.registers[13][31] ;
 wire \core_pipeline.pipeline_registers.registers[13][3] ;
 wire \core_pipeline.pipeline_registers.registers[13][4] ;
 wire \core_pipeline.pipeline_registers.registers[13][5] ;
 wire \core_pipeline.pipeline_registers.registers[13][6] ;
 wire \core_pipeline.pipeline_registers.registers[13][7] ;
 wire \core_pipeline.pipeline_registers.registers[13][8] ;
 wire \core_pipeline.pipeline_registers.registers[13][9] ;
 wire \core_pipeline.pipeline_registers.registers[14][0] ;
 wire \core_pipeline.pipeline_registers.registers[14][10] ;
 wire \core_pipeline.pipeline_registers.registers[14][11] ;
 wire \core_pipeline.pipeline_registers.registers[14][12] ;
 wire \core_pipeline.pipeline_registers.registers[14][13] ;
 wire \core_pipeline.pipeline_registers.registers[14][14] ;
 wire \core_pipeline.pipeline_registers.registers[14][15] ;
 wire \core_pipeline.pipeline_registers.registers[14][16] ;
 wire \core_pipeline.pipeline_registers.registers[14][17] ;
 wire \core_pipeline.pipeline_registers.registers[14][18] ;
 wire \core_pipeline.pipeline_registers.registers[14][19] ;
 wire \core_pipeline.pipeline_registers.registers[14][1] ;
 wire \core_pipeline.pipeline_registers.registers[14][20] ;
 wire \core_pipeline.pipeline_registers.registers[14][21] ;
 wire \core_pipeline.pipeline_registers.registers[14][22] ;
 wire \core_pipeline.pipeline_registers.registers[14][23] ;
 wire \core_pipeline.pipeline_registers.registers[14][24] ;
 wire \core_pipeline.pipeline_registers.registers[14][25] ;
 wire \core_pipeline.pipeline_registers.registers[14][26] ;
 wire \core_pipeline.pipeline_registers.registers[14][27] ;
 wire \core_pipeline.pipeline_registers.registers[14][28] ;
 wire \core_pipeline.pipeline_registers.registers[14][29] ;
 wire \core_pipeline.pipeline_registers.registers[14][2] ;
 wire \core_pipeline.pipeline_registers.registers[14][30] ;
 wire \core_pipeline.pipeline_registers.registers[14][31] ;
 wire \core_pipeline.pipeline_registers.registers[14][3] ;
 wire \core_pipeline.pipeline_registers.registers[14][4] ;
 wire \core_pipeline.pipeline_registers.registers[14][5] ;
 wire \core_pipeline.pipeline_registers.registers[14][6] ;
 wire \core_pipeline.pipeline_registers.registers[14][7] ;
 wire \core_pipeline.pipeline_registers.registers[14][8] ;
 wire \core_pipeline.pipeline_registers.registers[14][9] ;
 wire \core_pipeline.pipeline_registers.registers[15][0] ;
 wire \core_pipeline.pipeline_registers.registers[15][10] ;
 wire \core_pipeline.pipeline_registers.registers[15][11] ;
 wire \core_pipeline.pipeline_registers.registers[15][12] ;
 wire \core_pipeline.pipeline_registers.registers[15][13] ;
 wire \core_pipeline.pipeline_registers.registers[15][14] ;
 wire \core_pipeline.pipeline_registers.registers[15][15] ;
 wire \core_pipeline.pipeline_registers.registers[15][16] ;
 wire \core_pipeline.pipeline_registers.registers[15][17] ;
 wire \core_pipeline.pipeline_registers.registers[15][18] ;
 wire \core_pipeline.pipeline_registers.registers[15][19] ;
 wire \core_pipeline.pipeline_registers.registers[15][1] ;
 wire \core_pipeline.pipeline_registers.registers[15][20] ;
 wire \core_pipeline.pipeline_registers.registers[15][21] ;
 wire \core_pipeline.pipeline_registers.registers[15][22] ;
 wire \core_pipeline.pipeline_registers.registers[15][23] ;
 wire \core_pipeline.pipeline_registers.registers[15][24] ;
 wire \core_pipeline.pipeline_registers.registers[15][25] ;
 wire \core_pipeline.pipeline_registers.registers[15][26] ;
 wire \core_pipeline.pipeline_registers.registers[15][27] ;
 wire \core_pipeline.pipeline_registers.registers[15][28] ;
 wire \core_pipeline.pipeline_registers.registers[15][29] ;
 wire \core_pipeline.pipeline_registers.registers[15][2] ;
 wire \core_pipeline.pipeline_registers.registers[15][30] ;
 wire \core_pipeline.pipeline_registers.registers[15][31] ;
 wire \core_pipeline.pipeline_registers.registers[15][3] ;
 wire \core_pipeline.pipeline_registers.registers[15][4] ;
 wire \core_pipeline.pipeline_registers.registers[15][5] ;
 wire \core_pipeline.pipeline_registers.registers[15][6] ;
 wire \core_pipeline.pipeline_registers.registers[15][7] ;
 wire \core_pipeline.pipeline_registers.registers[15][8] ;
 wire \core_pipeline.pipeline_registers.registers[15][9] ;
 wire \core_pipeline.pipeline_registers.registers[16][0] ;
 wire \core_pipeline.pipeline_registers.registers[16][10] ;
 wire \core_pipeline.pipeline_registers.registers[16][11] ;
 wire \core_pipeline.pipeline_registers.registers[16][12] ;
 wire \core_pipeline.pipeline_registers.registers[16][13] ;
 wire \core_pipeline.pipeline_registers.registers[16][14] ;
 wire \core_pipeline.pipeline_registers.registers[16][15] ;
 wire \core_pipeline.pipeline_registers.registers[16][16] ;
 wire \core_pipeline.pipeline_registers.registers[16][17] ;
 wire \core_pipeline.pipeline_registers.registers[16][18] ;
 wire \core_pipeline.pipeline_registers.registers[16][19] ;
 wire \core_pipeline.pipeline_registers.registers[16][1] ;
 wire \core_pipeline.pipeline_registers.registers[16][20] ;
 wire \core_pipeline.pipeline_registers.registers[16][21] ;
 wire \core_pipeline.pipeline_registers.registers[16][22] ;
 wire \core_pipeline.pipeline_registers.registers[16][23] ;
 wire \core_pipeline.pipeline_registers.registers[16][24] ;
 wire \core_pipeline.pipeline_registers.registers[16][25] ;
 wire \core_pipeline.pipeline_registers.registers[16][26] ;
 wire \core_pipeline.pipeline_registers.registers[16][27] ;
 wire \core_pipeline.pipeline_registers.registers[16][28] ;
 wire \core_pipeline.pipeline_registers.registers[16][29] ;
 wire \core_pipeline.pipeline_registers.registers[16][2] ;
 wire \core_pipeline.pipeline_registers.registers[16][30] ;
 wire \core_pipeline.pipeline_registers.registers[16][31] ;
 wire \core_pipeline.pipeline_registers.registers[16][3] ;
 wire \core_pipeline.pipeline_registers.registers[16][4] ;
 wire \core_pipeline.pipeline_registers.registers[16][5] ;
 wire \core_pipeline.pipeline_registers.registers[16][6] ;
 wire \core_pipeline.pipeline_registers.registers[16][7] ;
 wire \core_pipeline.pipeline_registers.registers[16][8] ;
 wire \core_pipeline.pipeline_registers.registers[16][9] ;
 wire \core_pipeline.pipeline_registers.registers[17][0] ;
 wire \core_pipeline.pipeline_registers.registers[17][10] ;
 wire \core_pipeline.pipeline_registers.registers[17][11] ;
 wire \core_pipeline.pipeline_registers.registers[17][12] ;
 wire \core_pipeline.pipeline_registers.registers[17][13] ;
 wire \core_pipeline.pipeline_registers.registers[17][14] ;
 wire \core_pipeline.pipeline_registers.registers[17][15] ;
 wire \core_pipeline.pipeline_registers.registers[17][16] ;
 wire \core_pipeline.pipeline_registers.registers[17][17] ;
 wire \core_pipeline.pipeline_registers.registers[17][18] ;
 wire \core_pipeline.pipeline_registers.registers[17][19] ;
 wire \core_pipeline.pipeline_registers.registers[17][1] ;
 wire \core_pipeline.pipeline_registers.registers[17][20] ;
 wire \core_pipeline.pipeline_registers.registers[17][21] ;
 wire \core_pipeline.pipeline_registers.registers[17][22] ;
 wire \core_pipeline.pipeline_registers.registers[17][23] ;
 wire \core_pipeline.pipeline_registers.registers[17][24] ;
 wire \core_pipeline.pipeline_registers.registers[17][25] ;
 wire \core_pipeline.pipeline_registers.registers[17][26] ;
 wire \core_pipeline.pipeline_registers.registers[17][27] ;
 wire \core_pipeline.pipeline_registers.registers[17][28] ;
 wire \core_pipeline.pipeline_registers.registers[17][29] ;
 wire \core_pipeline.pipeline_registers.registers[17][2] ;
 wire \core_pipeline.pipeline_registers.registers[17][30] ;
 wire \core_pipeline.pipeline_registers.registers[17][31] ;
 wire \core_pipeline.pipeline_registers.registers[17][3] ;
 wire \core_pipeline.pipeline_registers.registers[17][4] ;
 wire \core_pipeline.pipeline_registers.registers[17][5] ;
 wire \core_pipeline.pipeline_registers.registers[17][6] ;
 wire \core_pipeline.pipeline_registers.registers[17][7] ;
 wire \core_pipeline.pipeline_registers.registers[17][8] ;
 wire \core_pipeline.pipeline_registers.registers[17][9] ;
 wire \core_pipeline.pipeline_registers.registers[18][0] ;
 wire \core_pipeline.pipeline_registers.registers[18][10] ;
 wire \core_pipeline.pipeline_registers.registers[18][11] ;
 wire \core_pipeline.pipeline_registers.registers[18][12] ;
 wire \core_pipeline.pipeline_registers.registers[18][13] ;
 wire \core_pipeline.pipeline_registers.registers[18][14] ;
 wire \core_pipeline.pipeline_registers.registers[18][15] ;
 wire \core_pipeline.pipeline_registers.registers[18][16] ;
 wire \core_pipeline.pipeline_registers.registers[18][17] ;
 wire \core_pipeline.pipeline_registers.registers[18][18] ;
 wire \core_pipeline.pipeline_registers.registers[18][19] ;
 wire \core_pipeline.pipeline_registers.registers[18][1] ;
 wire \core_pipeline.pipeline_registers.registers[18][20] ;
 wire \core_pipeline.pipeline_registers.registers[18][21] ;
 wire \core_pipeline.pipeline_registers.registers[18][22] ;
 wire \core_pipeline.pipeline_registers.registers[18][23] ;
 wire \core_pipeline.pipeline_registers.registers[18][24] ;
 wire \core_pipeline.pipeline_registers.registers[18][25] ;
 wire \core_pipeline.pipeline_registers.registers[18][26] ;
 wire \core_pipeline.pipeline_registers.registers[18][27] ;
 wire \core_pipeline.pipeline_registers.registers[18][28] ;
 wire \core_pipeline.pipeline_registers.registers[18][29] ;
 wire \core_pipeline.pipeline_registers.registers[18][2] ;
 wire \core_pipeline.pipeline_registers.registers[18][30] ;
 wire \core_pipeline.pipeline_registers.registers[18][31] ;
 wire \core_pipeline.pipeline_registers.registers[18][3] ;
 wire \core_pipeline.pipeline_registers.registers[18][4] ;
 wire \core_pipeline.pipeline_registers.registers[18][5] ;
 wire \core_pipeline.pipeline_registers.registers[18][6] ;
 wire \core_pipeline.pipeline_registers.registers[18][7] ;
 wire \core_pipeline.pipeline_registers.registers[18][8] ;
 wire \core_pipeline.pipeline_registers.registers[18][9] ;
 wire \core_pipeline.pipeline_registers.registers[19][0] ;
 wire \core_pipeline.pipeline_registers.registers[19][10] ;
 wire \core_pipeline.pipeline_registers.registers[19][11] ;
 wire \core_pipeline.pipeline_registers.registers[19][12] ;
 wire \core_pipeline.pipeline_registers.registers[19][13] ;
 wire \core_pipeline.pipeline_registers.registers[19][14] ;
 wire \core_pipeline.pipeline_registers.registers[19][15] ;
 wire \core_pipeline.pipeline_registers.registers[19][16] ;
 wire \core_pipeline.pipeline_registers.registers[19][17] ;
 wire \core_pipeline.pipeline_registers.registers[19][18] ;
 wire \core_pipeline.pipeline_registers.registers[19][19] ;
 wire \core_pipeline.pipeline_registers.registers[19][1] ;
 wire \core_pipeline.pipeline_registers.registers[19][20] ;
 wire \core_pipeline.pipeline_registers.registers[19][21] ;
 wire \core_pipeline.pipeline_registers.registers[19][22] ;
 wire \core_pipeline.pipeline_registers.registers[19][23] ;
 wire \core_pipeline.pipeline_registers.registers[19][24] ;
 wire \core_pipeline.pipeline_registers.registers[19][25] ;
 wire \core_pipeline.pipeline_registers.registers[19][26] ;
 wire \core_pipeline.pipeline_registers.registers[19][27] ;
 wire \core_pipeline.pipeline_registers.registers[19][28] ;
 wire \core_pipeline.pipeline_registers.registers[19][29] ;
 wire \core_pipeline.pipeline_registers.registers[19][2] ;
 wire \core_pipeline.pipeline_registers.registers[19][30] ;
 wire \core_pipeline.pipeline_registers.registers[19][31] ;
 wire \core_pipeline.pipeline_registers.registers[19][3] ;
 wire \core_pipeline.pipeline_registers.registers[19][4] ;
 wire \core_pipeline.pipeline_registers.registers[19][5] ;
 wire \core_pipeline.pipeline_registers.registers[19][6] ;
 wire \core_pipeline.pipeline_registers.registers[19][7] ;
 wire \core_pipeline.pipeline_registers.registers[19][8] ;
 wire \core_pipeline.pipeline_registers.registers[19][9] ;
 wire \core_pipeline.pipeline_registers.registers[1][0] ;
 wire \core_pipeline.pipeline_registers.registers[1][10] ;
 wire \core_pipeline.pipeline_registers.registers[1][11] ;
 wire \core_pipeline.pipeline_registers.registers[1][12] ;
 wire \core_pipeline.pipeline_registers.registers[1][13] ;
 wire \core_pipeline.pipeline_registers.registers[1][14] ;
 wire \core_pipeline.pipeline_registers.registers[1][15] ;
 wire \core_pipeline.pipeline_registers.registers[1][16] ;
 wire \core_pipeline.pipeline_registers.registers[1][17] ;
 wire \core_pipeline.pipeline_registers.registers[1][18] ;
 wire \core_pipeline.pipeline_registers.registers[1][19] ;
 wire \core_pipeline.pipeline_registers.registers[1][1] ;
 wire \core_pipeline.pipeline_registers.registers[1][20] ;
 wire \core_pipeline.pipeline_registers.registers[1][21] ;
 wire \core_pipeline.pipeline_registers.registers[1][22] ;
 wire \core_pipeline.pipeline_registers.registers[1][23] ;
 wire \core_pipeline.pipeline_registers.registers[1][24] ;
 wire \core_pipeline.pipeline_registers.registers[1][25] ;
 wire \core_pipeline.pipeline_registers.registers[1][26] ;
 wire \core_pipeline.pipeline_registers.registers[1][27] ;
 wire \core_pipeline.pipeline_registers.registers[1][28] ;
 wire \core_pipeline.pipeline_registers.registers[1][29] ;
 wire \core_pipeline.pipeline_registers.registers[1][2] ;
 wire \core_pipeline.pipeline_registers.registers[1][30] ;
 wire \core_pipeline.pipeline_registers.registers[1][31] ;
 wire \core_pipeline.pipeline_registers.registers[1][3] ;
 wire \core_pipeline.pipeline_registers.registers[1][4] ;
 wire \core_pipeline.pipeline_registers.registers[1][5] ;
 wire \core_pipeline.pipeline_registers.registers[1][6] ;
 wire \core_pipeline.pipeline_registers.registers[1][7] ;
 wire \core_pipeline.pipeline_registers.registers[1][8] ;
 wire \core_pipeline.pipeline_registers.registers[1][9] ;
 wire \core_pipeline.pipeline_registers.registers[20][0] ;
 wire \core_pipeline.pipeline_registers.registers[20][10] ;
 wire \core_pipeline.pipeline_registers.registers[20][11] ;
 wire \core_pipeline.pipeline_registers.registers[20][12] ;
 wire \core_pipeline.pipeline_registers.registers[20][13] ;
 wire \core_pipeline.pipeline_registers.registers[20][14] ;
 wire \core_pipeline.pipeline_registers.registers[20][15] ;
 wire \core_pipeline.pipeline_registers.registers[20][16] ;
 wire \core_pipeline.pipeline_registers.registers[20][17] ;
 wire \core_pipeline.pipeline_registers.registers[20][18] ;
 wire \core_pipeline.pipeline_registers.registers[20][19] ;
 wire \core_pipeline.pipeline_registers.registers[20][1] ;
 wire \core_pipeline.pipeline_registers.registers[20][20] ;
 wire \core_pipeline.pipeline_registers.registers[20][21] ;
 wire \core_pipeline.pipeline_registers.registers[20][22] ;
 wire \core_pipeline.pipeline_registers.registers[20][23] ;
 wire \core_pipeline.pipeline_registers.registers[20][24] ;
 wire \core_pipeline.pipeline_registers.registers[20][25] ;
 wire \core_pipeline.pipeline_registers.registers[20][26] ;
 wire \core_pipeline.pipeline_registers.registers[20][27] ;
 wire \core_pipeline.pipeline_registers.registers[20][28] ;
 wire \core_pipeline.pipeline_registers.registers[20][29] ;
 wire \core_pipeline.pipeline_registers.registers[20][2] ;
 wire \core_pipeline.pipeline_registers.registers[20][30] ;
 wire \core_pipeline.pipeline_registers.registers[20][31] ;
 wire \core_pipeline.pipeline_registers.registers[20][3] ;
 wire \core_pipeline.pipeline_registers.registers[20][4] ;
 wire \core_pipeline.pipeline_registers.registers[20][5] ;
 wire \core_pipeline.pipeline_registers.registers[20][6] ;
 wire \core_pipeline.pipeline_registers.registers[20][7] ;
 wire \core_pipeline.pipeline_registers.registers[20][8] ;
 wire \core_pipeline.pipeline_registers.registers[20][9] ;
 wire \core_pipeline.pipeline_registers.registers[21][0] ;
 wire \core_pipeline.pipeline_registers.registers[21][10] ;
 wire \core_pipeline.pipeline_registers.registers[21][11] ;
 wire \core_pipeline.pipeline_registers.registers[21][12] ;
 wire \core_pipeline.pipeline_registers.registers[21][13] ;
 wire \core_pipeline.pipeline_registers.registers[21][14] ;
 wire \core_pipeline.pipeline_registers.registers[21][15] ;
 wire \core_pipeline.pipeline_registers.registers[21][16] ;
 wire \core_pipeline.pipeline_registers.registers[21][17] ;
 wire \core_pipeline.pipeline_registers.registers[21][18] ;
 wire \core_pipeline.pipeline_registers.registers[21][19] ;
 wire \core_pipeline.pipeline_registers.registers[21][1] ;
 wire \core_pipeline.pipeline_registers.registers[21][20] ;
 wire \core_pipeline.pipeline_registers.registers[21][21] ;
 wire \core_pipeline.pipeline_registers.registers[21][22] ;
 wire \core_pipeline.pipeline_registers.registers[21][23] ;
 wire \core_pipeline.pipeline_registers.registers[21][24] ;
 wire \core_pipeline.pipeline_registers.registers[21][25] ;
 wire \core_pipeline.pipeline_registers.registers[21][26] ;
 wire \core_pipeline.pipeline_registers.registers[21][27] ;
 wire \core_pipeline.pipeline_registers.registers[21][28] ;
 wire \core_pipeline.pipeline_registers.registers[21][29] ;
 wire \core_pipeline.pipeline_registers.registers[21][2] ;
 wire \core_pipeline.pipeline_registers.registers[21][30] ;
 wire \core_pipeline.pipeline_registers.registers[21][31] ;
 wire \core_pipeline.pipeline_registers.registers[21][3] ;
 wire \core_pipeline.pipeline_registers.registers[21][4] ;
 wire \core_pipeline.pipeline_registers.registers[21][5] ;
 wire \core_pipeline.pipeline_registers.registers[21][6] ;
 wire \core_pipeline.pipeline_registers.registers[21][7] ;
 wire \core_pipeline.pipeline_registers.registers[21][8] ;
 wire \core_pipeline.pipeline_registers.registers[21][9] ;
 wire \core_pipeline.pipeline_registers.registers[22][0] ;
 wire \core_pipeline.pipeline_registers.registers[22][10] ;
 wire \core_pipeline.pipeline_registers.registers[22][11] ;
 wire \core_pipeline.pipeline_registers.registers[22][12] ;
 wire \core_pipeline.pipeline_registers.registers[22][13] ;
 wire \core_pipeline.pipeline_registers.registers[22][14] ;
 wire \core_pipeline.pipeline_registers.registers[22][15] ;
 wire \core_pipeline.pipeline_registers.registers[22][16] ;
 wire \core_pipeline.pipeline_registers.registers[22][17] ;
 wire \core_pipeline.pipeline_registers.registers[22][18] ;
 wire \core_pipeline.pipeline_registers.registers[22][19] ;
 wire \core_pipeline.pipeline_registers.registers[22][1] ;
 wire \core_pipeline.pipeline_registers.registers[22][20] ;
 wire \core_pipeline.pipeline_registers.registers[22][21] ;
 wire \core_pipeline.pipeline_registers.registers[22][22] ;
 wire \core_pipeline.pipeline_registers.registers[22][23] ;
 wire \core_pipeline.pipeline_registers.registers[22][24] ;
 wire \core_pipeline.pipeline_registers.registers[22][25] ;
 wire \core_pipeline.pipeline_registers.registers[22][26] ;
 wire \core_pipeline.pipeline_registers.registers[22][27] ;
 wire \core_pipeline.pipeline_registers.registers[22][28] ;
 wire \core_pipeline.pipeline_registers.registers[22][29] ;
 wire \core_pipeline.pipeline_registers.registers[22][2] ;
 wire \core_pipeline.pipeline_registers.registers[22][30] ;
 wire \core_pipeline.pipeline_registers.registers[22][31] ;
 wire \core_pipeline.pipeline_registers.registers[22][3] ;
 wire \core_pipeline.pipeline_registers.registers[22][4] ;
 wire \core_pipeline.pipeline_registers.registers[22][5] ;
 wire \core_pipeline.pipeline_registers.registers[22][6] ;
 wire \core_pipeline.pipeline_registers.registers[22][7] ;
 wire \core_pipeline.pipeline_registers.registers[22][8] ;
 wire \core_pipeline.pipeline_registers.registers[22][9] ;
 wire \core_pipeline.pipeline_registers.registers[23][0] ;
 wire \core_pipeline.pipeline_registers.registers[23][10] ;
 wire \core_pipeline.pipeline_registers.registers[23][11] ;
 wire \core_pipeline.pipeline_registers.registers[23][12] ;
 wire \core_pipeline.pipeline_registers.registers[23][13] ;
 wire \core_pipeline.pipeline_registers.registers[23][14] ;
 wire \core_pipeline.pipeline_registers.registers[23][15] ;
 wire \core_pipeline.pipeline_registers.registers[23][16] ;
 wire \core_pipeline.pipeline_registers.registers[23][17] ;
 wire \core_pipeline.pipeline_registers.registers[23][18] ;
 wire \core_pipeline.pipeline_registers.registers[23][19] ;
 wire \core_pipeline.pipeline_registers.registers[23][1] ;
 wire \core_pipeline.pipeline_registers.registers[23][20] ;
 wire \core_pipeline.pipeline_registers.registers[23][21] ;
 wire \core_pipeline.pipeline_registers.registers[23][22] ;
 wire \core_pipeline.pipeline_registers.registers[23][23] ;
 wire \core_pipeline.pipeline_registers.registers[23][24] ;
 wire \core_pipeline.pipeline_registers.registers[23][25] ;
 wire \core_pipeline.pipeline_registers.registers[23][26] ;
 wire \core_pipeline.pipeline_registers.registers[23][27] ;
 wire \core_pipeline.pipeline_registers.registers[23][28] ;
 wire \core_pipeline.pipeline_registers.registers[23][29] ;
 wire \core_pipeline.pipeline_registers.registers[23][2] ;
 wire \core_pipeline.pipeline_registers.registers[23][30] ;
 wire \core_pipeline.pipeline_registers.registers[23][31] ;
 wire \core_pipeline.pipeline_registers.registers[23][3] ;
 wire \core_pipeline.pipeline_registers.registers[23][4] ;
 wire \core_pipeline.pipeline_registers.registers[23][5] ;
 wire \core_pipeline.pipeline_registers.registers[23][6] ;
 wire \core_pipeline.pipeline_registers.registers[23][7] ;
 wire \core_pipeline.pipeline_registers.registers[23][8] ;
 wire \core_pipeline.pipeline_registers.registers[23][9] ;
 wire \core_pipeline.pipeline_registers.registers[24][0] ;
 wire \core_pipeline.pipeline_registers.registers[24][10] ;
 wire \core_pipeline.pipeline_registers.registers[24][11] ;
 wire \core_pipeline.pipeline_registers.registers[24][12] ;
 wire \core_pipeline.pipeline_registers.registers[24][13] ;
 wire \core_pipeline.pipeline_registers.registers[24][14] ;
 wire \core_pipeline.pipeline_registers.registers[24][15] ;
 wire \core_pipeline.pipeline_registers.registers[24][16] ;
 wire \core_pipeline.pipeline_registers.registers[24][17] ;
 wire \core_pipeline.pipeline_registers.registers[24][18] ;
 wire \core_pipeline.pipeline_registers.registers[24][19] ;
 wire \core_pipeline.pipeline_registers.registers[24][1] ;
 wire \core_pipeline.pipeline_registers.registers[24][20] ;
 wire \core_pipeline.pipeline_registers.registers[24][21] ;
 wire \core_pipeline.pipeline_registers.registers[24][22] ;
 wire \core_pipeline.pipeline_registers.registers[24][23] ;
 wire \core_pipeline.pipeline_registers.registers[24][24] ;
 wire \core_pipeline.pipeline_registers.registers[24][25] ;
 wire \core_pipeline.pipeline_registers.registers[24][26] ;
 wire \core_pipeline.pipeline_registers.registers[24][27] ;
 wire \core_pipeline.pipeline_registers.registers[24][28] ;
 wire \core_pipeline.pipeline_registers.registers[24][29] ;
 wire \core_pipeline.pipeline_registers.registers[24][2] ;
 wire \core_pipeline.pipeline_registers.registers[24][30] ;
 wire \core_pipeline.pipeline_registers.registers[24][31] ;
 wire \core_pipeline.pipeline_registers.registers[24][3] ;
 wire \core_pipeline.pipeline_registers.registers[24][4] ;
 wire \core_pipeline.pipeline_registers.registers[24][5] ;
 wire \core_pipeline.pipeline_registers.registers[24][6] ;
 wire \core_pipeline.pipeline_registers.registers[24][7] ;
 wire \core_pipeline.pipeline_registers.registers[24][8] ;
 wire \core_pipeline.pipeline_registers.registers[24][9] ;
 wire \core_pipeline.pipeline_registers.registers[25][0] ;
 wire \core_pipeline.pipeline_registers.registers[25][10] ;
 wire \core_pipeline.pipeline_registers.registers[25][11] ;
 wire \core_pipeline.pipeline_registers.registers[25][12] ;
 wire \core_pipeline.pipeline_registers.registers[25][13] ;
 wire \core_pipeline.pipeline_registers.registers[25][14] ;
 wire \core_pipeline.pipeline_registers.registers[25][15] ;
 wire \core_pipeline.pipeline_registers.registers[25][16] ;
 wire \core_pipeline.pipeline_registers.registers[25][17] ;
 wire \core_pipeline.pipeline_registers.registers[25][18] ;
 wire \core_pipeline.pipeline_registers.registers[25][19] ;
 wire \core_pipeline.pipeline_registers.registers[25][1] ;
 wire \core_pipeline.pipeline_registers.registers[25][20] ;
 wire \core_pipeline.pipeline_registers.registers[25][21] ;
 wire \core_pipeline.pipeline_registers.registers[25][22] ;
 wire \core_pipeline.pipeline_registers.registers[25][23] ;
 wire \core_pipeline.pipeline_registers.registers[25][24] ;
 wire \core_pipeline.pipeline_registers.registers[25][25] ;
 wire \core_pipeline.pipeline_registers.registers[25][26] ;
 wire \core_pipeline.pipeline_registers.registers[25][27] ;
 wire \core_pipeline.pipeline_registers.registers[25][28] ;
 wire \core_pipeline.pipeline_registers.registers[25][29] ;
 wire \core_pipeline.pipeline_registers.registers[25][2] ;
 wire \core_pipeline.pipeline_registers.registers[25][30] ;
 wire \core_pipeline.pipeline_registers.registers[25][31] ;
 wire \core_pipeline.pipeline_registers.registers[25][3] ;
 wire \core_pipeline.pipeline_registers.registers[25][4] ;
 wire \core_pipeline.pipeline_registers.registers[25][5] ;
 wire \core_pipeline.pipeline_registers.registers[25][6] ;
 wire \core_pipeline.pipeline_registers.registers[25][7] ;
 wire \core_pipeline.pipeline_registers.registers[25][8] ;
 wire \core_pipeline.pipeline_registers.registers[25][9] ;
 wire \core_pipeline.pipeline_registers.registers[26][0] ;
 wire \core_pipeline.pipeline_registers.registers[26][10] ;
 wire \core_pipeline.pipeline_registers.registers[26][11] ;
 wire \core_pipeline.pipeline_registers.registers[26][12] ;
 wire \core_pipeline.pipeline_registers.registers[26][13] ;
 wire \core_pipeline.pipeline_registers.registers[26][14] ;
 wire \core_pipeline.pipeline_registers.registers[26][15] ;
 wire \core_pipeline.pipeline_registers.registers[26][16] ;
 wire \core_pipeline.pipeline_registers.registers[26][17] ;
 wire \core_pipeline.pipeline_registers.registers[26][18] ;
 wire \core_pipeline.pipeline_registers.registers[26][19] ;
 wire \core_pipeline.pipeline_registers.registers[26][1] ;
 wire \core_pipeline.pipeline_registers.registers[26][20] ;
 wire \core_pipeline.pipeline_registers.registers[26][21] ;
 wire \core_pipeline.pipeline_registers.registers[26][22] ;
 wire \core_pipeline.pipeline_registers.registers[26][23] ;
 wire \core_pipeline.pipeline_registers.registers[26][24] ;
 wire \core_pipeline.pipeline_registers.registers[26][25] ;
 wire \core_pipeline.pipeline_registers.registers[26][26] ;
 wire \core_pipeline.pipeline_registers.registers[26][27] ;
 wire \core_pipeline.pipeline_registers.registers[26][28] ;
 wire \core_pipeline.pipeline_registers.registers[26][29] ;
 wire \core_pipeline.pipeline_registers.registers[26][2] ;
 wire \core_pipeline.pipeline_registers.registers[26][30] ;
 wire \core_pipeline.pipeline_registers.registers[26][31] ;
 wire \core_pipeline.pipeline_registers.registers[26][3] ;
 wire \core_pipeline.pipeline_registers.registers[26][4] ;
 wire \core_pipeline.pipeline_registers.registers[26][5] ;
 wire \core_pipeline.pipeline_registers.registers[26][6] ;
 wire \core_pipeline.pipeline_registers.registers[26][7] ;
 wire \core_pipeline.pipeline_registers.registers[26][8] ;
 wire \core_pipeline.pipeline_registers.registers[26][9] ;
 wire \core_pipeline.pipeline_registers.registers[27][0] ;
 wire \core_pipeline.pipeline_registers.registers[27][10] ;
 wire \core_pipeline.pipeline_registers.registers[27][11] ;
 wire \core_pipeline.pipeline_registers.registers[27][12] ;
 wire \core_pipeline.pipeline_registers.registers[27][13] ;
 wire \core_pipeline.pipeline_registers.registers[27][14] ;
 wire \core_pipeline.pipeline_registers.registers[27][15] ;
 wire \core_pipeline.pipeline_registers.registers[27][16] ;
 wire \core_pipeline.pipeline_registers.registers[27][17] ;
 wire \core_pipeline.pipeline_registers.registers[27][18] ;
 wire \core_pipeline.pipeline_registers.registers[27][19] ;
 wire \core_pipeline.pipeline_registers.registers[27][1] ;
 wire \core_pipeline.pipeline_registers.registers[27][20] ;
 wire \core_pipeline.pipeline_registers.registers[27][21] ;
 wire \core_pipeline.pipeline_registers.registers[27][22] ;
 wire \core_pipeline.pipeline_registers.registers[27][23] ;
 wire \core_pipeline.pipeline_registers.registers[27][24] ;
 wire \core_pipeline.pipeline_registers.registers[27][25] ;
 wire \core_pipeline.pipeline_registers.registers[27][26] ;
 wire \core_pipeline.pipeline_registers.registers[27][27] ;
 wire \core_pipeline.pipeline_registers.registers[27][28] ;
 wire \core_pipeline.pipeline_registers.registers[27][29] ;
 wire \core_pipeline.pipeline_registers.registers[27][2] ;
 wire \core_pipeline.pipeline_registers.registers[27][30] ;
 wire \core_pipeline.pipeline_registers.registers[27][31] ;
 wire \core_pipeline.pipeline_registers.registers[27][3] ;
 wire \core_pipeline.pipeline_registers.registers[27][4] ;
 wire \core_pipeline.pipeline_registers.registers[27][5] ;
 wire \core_pipeline.pipeline_registers.registers[27][6] ;
 wire \core_pipeline.pipeline_registers.registers[27][7] ;
 wire \core_pipeline.pipeline_registers.registers[27][8] ;
 wire \core_pipeline.pipeline_registers.registers[27][9] ;
 wire \core_pipeline.pipeline_registers.registers[28][0] ;
 wire \core_pipeline.pipeline_registers.registers[28][10] ;
 wire \core_pipeline.pipeline_registers.registers[28][11] ;
 wire \core_pipeline.pipeline_registers.registers[28][12] ;
 wire \core_pipeline.pipeline_registers.registers[28][13] ;
 wire \core_pipeline.pipeline_registers.registers[28][14] ;
 wire \core_pipeline.pipeline_registers.registers[28][15] ;
 wire \core_pipeline.pipeline_registers.registers[28][16] ;
 wire \core_pipeline.pipeline_registers.registers[28][17] ;
 wire \core_pipeline.pipeline_registers.registers[28][18] ;
 wire \core_pipeline.pipeline_registers.registers[28][19] ;
 wire \core_pipeline.pipeline_registers.registers[28][1] ;
 wire \core_pipeline.pipeline_registers.registers[28][20] ;
 wire \core_pipeline.pipeline_registers.registers[28][21] ;
 wire \core_pipeline.pipeline_registers.registers[28][22] ;
 wire \core_pipeline.pipeline_registers.registers[28][23] ;
 wire \core_pipeline.pipeline_registers.registers[28][24] ;
 wire \core_pipeline.pipeline_registers.registers[28][25] ;
 wire \core_pipeline.pipeline_registers.registers[28][26] ;
 wire \core_pipeline.pipeline_registers.registers[28][27] ;
 wire \core_pipeline.pipeline_registers.registers[28][28] ;
 wire \core_pipeline.pipeline_registers.registers[28][29] ;
 wire \core_pipeline.pipeline_registers.registers[28][2] ;
 wire \core_pipeline.pipeline_registers.registers[28][30] ;
 wire \core_pipeline.pipeline_registers.registers[28][31] ;
 wire \core_pipeline.pipeline_registers.registers[28][3] ;
 wire \core_pipeline.pipeline_registers.registers[28][4] ;
 wire \core_pipeline.pipeline_registers.registers[28][5] ;
 wire \core_pipeline.pipeline_registers.registers[28][6] ;
 wire \core_pipeline.pipeline_registers.registers[28][7] ;
 wire \core_pipeline.pipeline_registers.registers[28][8] ;
 wire \core_pipeline.pipeline_registers.registers[28][9] ;
 wire \core_pipeline.pipeline_registers.registers[29][0] ;
 wire \core_pipeline.pipeline_registers.registers[29][10] ;
 wire \core_pipeline.pipeline_registers.registers[29][11] ;
 wire \core_pipeline.pipeline_registers.registers[29][12] ;
 wire \core_pipeline.pipeline_registers.registers[29][13] ;
 wire \core_pipeline.pipeline_registers.registers[29][14] ;
 wire \core_pipeline.pipeline_registers.registers[29][15] ;
 wire \core_pipeline.pipeline_registers.registers[29][16] ;
 wire \core_pipeline.pipeline_registers.registers[29][17] ;
 wire \core_pipeline.pipeline_registers.registers[29][18] ;
 wire \core_pipeline.pipeline_registers.registers[29][19] ;
 wire \core_pipeline.pipeline_registers.registers[29][1] ;
 wire \core_pipeline.pipeline_registers.registers[29][20] ;
 wire \core_pipeline.pipeline_registers.registers[29][21] ;
 wire \core_pipeline.pipeline_registers.registers[29][22] ;
 wire \core_pipeline.pipeline_registers.registers[29][23] ;
 wire \core_pipeline.pipeline_registers.registers[29][24] ;
 wire \core_pipeline.pipeline_registers.registers[29][25] ;
 wire \core_pipeline.pipeline_registers.registers[29][26] ;
 wire \core_pipeline.pipeline_registers.registers[29][27] ;
 wire \core_pipeline.pipeline_registers.registers[29][28] ;
 wire \core_pipeline.pipeline_registers.registers[29][29] ;
 wire \core_pipeline.pipeline_registers.registers[29][2] ;
 wire \core_pipeline.pipeline_registers.registers[29][30] ;
 wire \core_pipeline.pipeline_registers.registers[29][31] ;
 wire \core_pipeline.pipeline_registers.registers[29][3] ;
 wire \core_pipeline.pipeline_registers.registers[29][4] ;
 wire \core_pipeline.pipeline_registers.registers[29][5] ;
 wire \core_pipeline.pipeline_registers.registers[29][6] ;
 wire \core_pipeline.pipeline_registers.registers[29][7] ;
 wire \core_pipeline.pipeline_registers.registers[29][8] ;
 wire \core_pipeline.pipeline_registers.registers[29][9] ;
 wire \core_pipeline.pipeline_registers.registers[2][0] ;
 wire \core_pipeline.pipeline_registers.registers[2][10] ;
 wire \core_pipeline.pipeline_registers.registers[2][11] ;
 wire \core_pipeline.pipeline_registers.registers[2][12] ;
 wire \core_pipeline.pipeline_registers.registers[2][13] ;
 wire \core_pipeline.pipeline_registers.registers[2][14] ;
 wire \core_pipeline.pipeline_registers.registers[2][15] ;
 wire \core_pipeline.pipeline_registers.registers[2][16] ;
 wire \core_pipeline.pipeline_registers.registers[2][17] ;
 wire \core_pipeline.pipeline_registers.registers[2][18] ;
 wire \core_pipeline.pipeline_registers.registers[2][19] ;
 wire \core_pipeline.pipeline_registers.registers[2][1] ;
 wire \core_pipeline.pipeline_registers.registers[2][20] ;
 wire \core_pipeline.pipeline_registers.registers[2][21] ;
 wire \core_pipeline.pipeline_registers.registers[2][22] ;
 wire \core_pipeline.pipeline_registers.registers[2][23] ;
 wire \core_pipeline.pipeline_registers.registers[2][24] ;
 wire \core_pipeline.pipeline_registers.registers[2][25] ;
 wire \core_pipeline.pipeline_registers.registers[2][26] ;
 wire \core_pipeline.pipeline_registers.registers[2][27] ;
 wire \core_pipeline.pipeline_registers.registers[2][28] ;
 wire \core_pipeline.pipeline_registers.registers[2][29] ;
 wire \core_pipeline.pipeline_registers.registers[2][2] ;
 wire \core_pipeline.pipeline_registers.registers[2][30] ;
 wire \core_pipeline.pipeline_registers.registers[2][31] ;
 wire \core_pipeline.pipeline_registers.registers[2][3] ;
 wire \core_pipeline.pipeline_registers.registers[2][4] ;
 wire \core_pipeline.pipeline_registers.registers[2][5] ;
 wire \core_pipeline.pipeline_registers.registers[2][6] ;
 wire \core_pipeline.pipeline_registers.registers[2][7] ;
 wire \core_pipeline.pipeline_registers.registers[2][8] ;
 wire \core_pipeline.pipeline_registers.registers[2][9] ;
 wire \core_pipeline.pipeline_registers.registers[30][0] ;
 wire \core_pipeline.pipeline_registers.registers[30][10] ;
 wire \core_pipeline.pipeline_registers.registers[30][11] ;
 wire \core_pipeline.pipeline_registers.registers[30][12] ;
 wire \core_pipeline.pipeline_registers.registers[30][13] ;
 wire \core_pipeline.pipeline_registers.registers[30][14] ;
 wire \core_pipeline.pipeline_registers.registers[30][15] ;
 wire \core_pipeline.pipeline_registers.registers[30][16] ;
 wire \core_pipeline.pipeline_registers.registers[30][17] ;
 wire \core_pipeline.pipeline_registers.registers[30][18] ;
 wire \core_pipeline.pipeline_registers.registers[30][19] ;
 wire \core_pipeline.pipeline_registers.registers[30][1] ;
 wire \core_pipeline.pipeline_registers.registers[30][20] ;
 wire \core_pipeline.pipeline_registers.registers[30][21] ;
 wire \core_pipeline.pipeline_registers.registers[30][22] ;
 wire \core_pipeline.pipeline_registers.registers[30][23] ;
 wire \core_pipeline.pipeline_registers.registers[30][24] ;
 wire \core_pipeline.pipeline_registers.registers[30][25] ;
 wire \core_pipeline.pipeline_registers.registers[30][26] ;
 wire \core_pipeline.pipeline_registers.registers[30][27] ;
 wire \core_pipeline.pipeline_registers.registers[30][28] ;
 wire \core_pipeline.pipeline_registers.registers[30][29] ;
 wire \core_pipeline.pipeline_registers.registers[30][2] ;
 wire \core_pipeline.pipeline_registers.registers[30][30] ;
 wire \core_pipeline.pipeline_registers.registers[30][31] ;
 wire \core_pipeline.pipeline_registers.registers[30][3] ;
 wire \core_pipeline.pipeline_registers.registers[30][4] ;
 wire \core_pipeline.pipeline_registers.registers[30][5] ;
 wire \core_pipeline.pipeline_registers.registers[30][6] ;
 wire \core_pipeline.pipeline_registers.registers[30][7] ;
 wire \core_pipeline.pipeline_registers.registers[30][8] ;
 wire \core_pipeline.pipeline_registers.registers[30][9] ;
 wire \core_pipeline.pipeline_registers.registers[31][0] ;
 wire \core_pipeline.pipeline_registers.registers[31][10] ;
 wire \core_pipeline.pipeline_registers.registers[31][11] ;
 wire \core_pipeline.pipeline_registers.registers[31][12] ;
 wire \core_pipeline.pipeline_registers.registers[31][13] ;
 wire \core_pipeline.pipeline_registers.registers[31][14] ;
 wire \core_pipeline.pipeline_registers.registers[31][15] ;
 wire \core_pipeline.pipeline_registers.registers[31][16] ;
 wire \core_pipeline.pipeline_registers.registers[31][17] ;
 wire \core_pipeline.pipeline_registers.registers[31][18] ;
 wire \core_pipeline.pipeline_registers.registers[31][19] ;
 wire \core_pipeline.pipeline_registers.registers[31][1] ;
 wire \core_pipeline.pipeline_registers.registers[31][20] ;
 wire \core_pipeline.pipeline_registers.registers[31][21] ;
 wire \core_pipeline.pipeline_registers.registers[31][22] ;
 wire \core_pipeline.pipeline_registers.registers[31][23] ;
 wire \core_pipeline.pipeline_registers.registers[31][24] ;
 wire \core_pipeline.pipeline_registers.registers[31][25] ;
 wire \core_pipeline.pipeline_registers.registers[31][26] ;
 wire \core_pipeline.pipeline_registers.registers[31][27] ;
 wire \core_pipeline.pipeline_registers.registers[31][28] ;
 wire \core_pipeline.pipeline_registers.registers[31][29] ;
 wire \core_pipeline.pipeline_registers.registers[31][2] ;
 wire \core_pipeline.pipeline_registers.registers[31][30] ;
 wire \core_pipeline.pipeline_registers.registers[31][31] ;
 wire \core_pipeline.pipeline_registers.registers[31][3] ;
 wire \core_pipeline.pipeline_registers.registers[31][4] ;
 wire \core_pipeline.pipeline_registers.registers[31][5] ;
 wire \core_pipeline.pipeline_registers.registers[31][6] ;
 wire \core_pipeline.pipeline_registers.registers[31][7] ;
 wire \core_pipeline.pipeline_registers.registers[31][8] ;
 wire \core_pipeline.pipeline_registers.registers[31][9] ;
 wire \core_pipeline.pipeline_registers.registers[3][0] ;
 wire \core_pipeline.pipeline_registers.registers[3][10] ;
 wire \core_pipeline.pipeline_registers.registers[3][11] ;
 wire \core_pipeline.pipeline_registers.registers[3][12] ;
 wire \core_pipeline.pipeline_registers.registers[3][13] ;
 wire \core_pipeline.pipeline_registers.registers[3][14] ;
 wire \core_pipeline.pipeline_registers.registers[3][15] ;
 wire \core_pipeline.pipeline_registers.registers[3][16] ;
 wire \core_pipeline.pipeline_registers.registers[3][17] ;
 wire \core_pipeline.pipeline_registers.registers[3][18] ;
 wire \core_pipeline.pipeline_registers.registers[3][19] ;
 wire \core_pipeline.pipeline_registers.registers[3][1] ;
 wire \core_pipeline.pipeline_registers.registers[3][20] ;
 wire \core_pipeline.pipeline_registers.registers[3][21] ;
 wire \core_pipeline.pipeline_registers.registers[3][22] ;
 wire \core_pipeline.pipeline_registers.registers[3][23] ;
 wire \core_pipeline.pipeline_registers.registers[3][24] ;
 wire \core_pipeline.pipeline_registers.registers[3][25] ;
 wire \core_pipeline.pipeline_registers.registers[3][26] ;
 wire \core_pipeline.pipeline_registers.registers[3][27] ;
 wire \core_pipeline.pipeline_registers.registers[3][28] ;
 wire \core_pipeline.pipeline_registers.registers[3][29] ;
 wire \core_pipeline.pipeline_registers.registers[3][2] ;
 wire \core_pipeline.pipeline_registers.registers[3][30] ;
 wire \core_pipeline.pipeline_registers.registers[3][31] ;
 wire \core_pipeline.pipeline_registers.registers[3][3] ;
 wire \core_pipeline.pipeline_registers.registers[3][4] ;
 wire \core_pipeline.pipeline_registers.registers[3][5] ;
 wire \core_pipeline.pipeline_registers.registers[3][6] ;
 wire \core_pipeline.pipeline_registers.registers[3][7] ;
 wire \core_pipeline.pipeline_registers.registers[3][8] ;
 wire \core_pipeline.pipeline_registers.registers[3][9] ;
 wire \core_pipeline.pipeline_registers.registers[4][0] ;
 wire \core_pipeline.pipeline_registers.registers[4][10] ;
 wire \core_pipeline.pipeline_registers.registers[4][11] ;
 wire \core_pipeline.pipeline_registers.registers[4][12] ;
 wire \core_pipeline.pipeline_registers.registers[4][13] ;
 wire \core_pipeline.pipeline_registers.registers[4][14] ;
 wire \core_pipeline.pipeline_registers.registers[4][15] ;
 wire \core_pipeline.pipeline_registers.registers[4][16] ;
 wire \core_pipeline.pipeline_registers.registers[4][17] ;
 wire \core_pipeline.pipeline_registers.registers[4][18] ;
 wire \core_pipeline.pipeline_registers.registers[4][19] ;
 wire \core_pipeline.pipeline_registers.registers[4][1] ;
 wire \core_pipeline.pipeline_registers.registers[4][20] ;
 wire \core_pipeline.pipeline_registers.registers[4][21] ;
 wire \core_pipeline.pipeline_registers.registers[4][22] ;
 wire \core_pipeline.pipeline_registers.registers[4][23] ;
 wire \core_pipeline.pipeline_registers.registers[4][24] ;
 wire \core_pipeline.pipeline_registers.registers[4][25] ;
 wire \core_pipeline.pipeline_registers.registers[4][26] ;
 wire \core_pipeline.pipeline_registers.registers[4][27] ;
 wire \core_pipeline.pipeline_registers.registers[4][28] ;
 wire \core_pipeline.pipeline_registers.registers[4][29] ;
 wire \core_pipeline.pipeline_registers.registers[4][2] ;
 wire \core_pipeline.pipeline_registers.registers[4][30] ;
 wire \core_pipeline.pipeline_registers.registers[4][31] ;
 wire \core_pipeline.pipeline_registers.registers[4][3] ;
 wire \core_pipeline.pipeline_registers.registers[4][4] ;
 wire \core_pipeline.pipeline_registers.registers[4][5] ;
 wire \core_pipeline.pipeline_registers.registers[4][6] ;
 wire \core_pipeline.pipeline_registers.registers[4][7] ;
 wire \core_pipeline.pipeline_registers.registers[4][8] ;
 wire \core_pipeline.pipeline_registers.registers[4][9] ;
 wire \core_pipeline.pipeline_registers.registers[5][0] ;
 wire \core_pipeline.pipeline_registers.registers[5][10] ;
 wire \core_pipeline.pipeline_registers.registers[5][11] ;
 wire \core_pipeline.pipeline_registers.registers[5][12] ;
 wire \core_pipeline.pipeline_registers.registers[5][13] ;
 wire \core_pipeline.pipeline_registers.registers[5][14] ;
 wire \core_pipeline.pipeline_registers.registers[5][15] ;
 wire \core_pipeline.pipeline_registers.registers[5][16] ;
 wire \core_pipeline.pipeline_registers.registers[5][17] ;
 wire \core_pipeline.pipeline_registers.registers[5][18] ;
 wire \core_pipeline.pipeline_registers.registers[5][19] ;
 wire \core_pipeline.pipeline_registers.registers[5][1] ;
 wire \core_pipeline.pipeline_registers.registers[5][20] ;
 wire \core_pipeline.pipeline_registers.registers[5][21] ;
 wire \core_pipeline.pipeline_registers.registers[5][22] ;
 wire \core_pipeline.pipeline_registers.registers[5][23] ;
 wire \core_pipeline.pipeline_registers.registers[5][24] ;
 wire \core_pipeline.pipeline_registers.registers[5][25] ;
 wire \core_pipeline.pipeline_registers.registers[5][26] ;
 wire \core_pipeline.pipeline_registers.registers[5][27] ;
 wire \core_pipeline.pipeline_registers.registers[5][28] ;
 wire \core_pipeline.pipeline_registers.registers[5][29] ;
 wire \core_pipeline.pipeline_registers.registers[5][2] ;
 wire \core_pipeline.pipeline_registers.registers[5][30] ;
 wire \core_pipeline.pipeline_registers.registers[5][31] ;
 wire \core_pipeline.pipeline_registers.registers[5][3] ;
 wire \core_pipeline.pipeline_registers.registers[5][4] ;
 wire \core_pipeline.pipeline_registers.registers[5][5] ;
 wire \core_pipeline.pipeline_registers.registers[5][6] ;
 wire \core_pipeline.pipeline_registers.registers[5][7] ;
 wire \core_pipeline.pipeline_registers.registers[5][8] ;
 wire \core_pipeline.pipeline_registers.registers[5][9] ;
 wire \core_pipeline.pipeline_registers.registers[6][0] ;
 wire \core_pipeline.pipeline_registers.registers[6][10] ;
 wire \core_pipeline.pipeline_registers.registers[6][11] ;
 wire \core_pipeline.pipeline_registers.registers[6][12] ;
 wire \core_pipeline.pipeline_registers.registers[6][13] ;
 wire \core_pipeline.pipeline_registers.registers[6][14] ;
 wire \core_pipeline.pipeline_registers.registers[6][15] ;
 wire \core_pipeline.pipeline_registers.registers[6][16] ;
 wire \core_pipeline.pipeline_registers.registers[6][17] ;
 wire \core_pipeline.pipeline_registers.registers[6][18] ;
 wire \core_pipeline.pipeline_registers.registers[6][19] ;
 wire \core_pipeline.pipeline_registers.registers[6][1] ;
 wire \core_pipeline.pipeline_registers.registers[6][20] ;
 wire \core_pipeline.pipeline_registers.registers[6][21] ;
 wire \core_pipeline.pipeline_registers.registers[6][22] ;
 wire \core_pipeline.pipeline_registers.registers[6][23] ;
 wire \core_pipeline.pipeline_registers.registers[6][24] ;
 wire \core_pipeline.pipeline_registers.registers[6][25] ;
 wire \core_pipeline.pipeline_registers.registers[6][26] ;
 wire \core_pipeline.pipeline_registers.registers[6][27] ;
 wire \core_pipeline.pipeline_registers.registers[6][28] ;
 wire \core_pipeline.pipeline_registers.registers[6][29] ;
 wire \core_pipeline.pipeline_registers.registers[6][2] ;
 wire \core_pipeline.pipeline_registers.registers[6][30] ;
 wire \core_pipeline.pipeline_registers.registers[6][31] ;
 wire \core_pipeline.pipeline_registers.registers[6][3] ;
 wire \core_pipeline.pipeline_registers.registers[6][4] ;
 wire \core_pipeline.pipeline_registers.registers[6][5] ;
 wire \core_pipeline.pipeline_registers.registers[6][6] ;
 wire \core_pipeline.pipeline_registers.registers[6][7] ;
 wire \core_pipeline.pipeline_registers.registers[6][8] ;
 wire \core_pipeline.pipeline_registers.registers[6][9] ;
 wire \core_pipeline.pipeline_registers.registers[7][0] ;
 wire \core_pipeline.pipeline_registers.registers[7][10] ;
 wire \core_pipeline.pipeline_registers.registers[7][11] ;
 wire \core_pipeline.pipeline_registers.registers[7][12] ;
 wire \core_pipeline.pipeline_registers.registers[7][13] ;
 wire \core_pipeline.pipeline_registers.registers[7][14] ;
 wire \core_pipeline.pipeline_registers.registers[7][15] ;
 wire \core_pipeline.pipeline_registers.registers[7][16] ;
 wire \core_pipeline.pipeline_registers.registers[7][17] ;
 wire \core_pipeline.pipeline_registers.registers[7][18] ;
 wire \core_pipeline.pipeline_registers.registers[7][19] ;
 wire \core_pipeline.pipeline_registers.registers[7][1] ;
 wire \core_pipeline.pipeline_registers.registers[7][20] ;
 wire \core_pipeline.pipeline_registers.registers[7][21] ;
 wire \core_pipeline.pipeline_registers.registers[7][22] ;
 wire \core_pipeline.pipeline_registers.registers[7][23] ;
 wire \core_pipeline.pipeline_registers.registers[7][24] ;
 wire \core_pipeline.pipeline_registers.registers[7][25] ;
 wire \core_pipeline.pipeline_registers.registers[7][26] ;
 wire \core_pipeline.pipeline_registers.registers[7][27] ;
 wire \core_pipeline.pipeline_registers.registers[7][28] ;
 wire \core_pipeline.pipeline_registers.registers[7][29] ;
 wire \core_pipeline.pipeline_registers.registers[7][2] ;
 wire \core_pipeline.pipeline_registers.registers[7][30] ;
 wire \core_pipeline.pipeline_registers.registers[7][31] ;
 wire \core_pipeline.pipeline_registers.registers[7][3] ;
 wire \core_pipeline.pipeline_registers.registers[7][4] ;
 wire \core_pipeline.pipeline_registers.registers[7][5] ;
 wire \core_pipeline.pipeline_registers.registers[7][6] ;
 wire \core_pipeline.pipeline_registers.registers[7][7] ;
 wire \core_pipeline.pipeline_registers.registers[7][8] ;
 wire \core_pipeline.pipeline_registers.registers[7][9] ;
 wire \core_pipeline.pipeline_registers.registers[8][0] ;
 wire \core_pipeline.pipeline_registers.registers[8][10] ;
 wire \core_pipeline.pipeline_registers.registers[8][11] ;
 wire \core_pipeline.pipeline_registers.registers[8][12] ;
 wire \core_pipeline.pipeline_registers.registers[8][13] ;
 wire \core_pipeline.pipeline_registers.registers[8][14] ;
 wire \core_pipeline.pipeline_registers.registers[8][15] ;
 wire \core_pipeline.pipeline_registers.registers[8][16] ;
 wire \core_pipeline.pipeline_registers.registers[8][17] ;
 wire \core_pipeline.pipeline_registers.registers[8][18] ;
 wire \core_pipeline.pipeline_registers.registers[8][19] ;
 wire \core_pipeline.pipeline_registers.registers[8][1] ;
 wire \core_pipeline.pipeline_registers.registers[8][20] ;
 wire \core_pipeline.pipeline_registers.registers[8][21] ;
 wire \core_pipeline.pipeline_registers.registers[8][22] ;
 wire \core_pipeline.pipeline_registers.registers[8][23] ;
 wire \core_pipeline.pipeline_registers.registers[8][24] ;
 wire \core_pipeline.pipeline_registers.registers[8][25] ;
 wire \core_pipeline.pipeline_registers.registers[8][26] ;
 wire \core_pipeline.pipeline_registers.registers[8][27] ;
 wire \core_pipeline.pipeline_registers.registers[8][28] ;
 wire \core_pipeline.pipeline_registers.registers[8][29] ;
 wire \core_pipeline.pipeline_registers.registers[8][2] ;
 wire \core_pipeline.pipeline_registers.registers[8][30] ;
 wire \core_pipeline.pipeline_registers.registers[8][31] ;
 wire \core_pipeline.pipeline_registers.registers[8][3] ;
 wire \core_pipeline.pipeline_registers.registers[8][4] ;
 wire \core_pipeline.pipeline_registers.registers[8][5] ;
 wire \core_pipeline.pipeline_registers.registers[8][6] ;
 wire \core_pipeline.pipeline_registers.registers[8][7] ;
 wire \core_pipeline.pipeline_registers.registers[8][8] ;
 wire \core_pipeline.pipeline_registers.registers[8][9] ;
 wire \core_pipeline.pipeline_registers.registers[9][0] ;
 wire \core_pipeline.pipeline_registers.registers[9][10] ;
 wire \core_pipeline.pipeline_registers.registers[9][11] ;
 wire \core_pipeline.pipeline_registers.registers[9][12] ;
 wire \core_pipeline.pipeline_registers.registers[9][13] ;
 wire \core_pipeline.pipeline_registers.registers[9][14] ;
 wire \core_pipeline.pipeline_registers.registers[9][15] ;
 wire \core_pipeline.pipeline_registers.registers[9][16] ;
 wire \core_pipeline.pipeline_registers.registers[9][17] ;
 wire \core_pipeline.pipeline_registers.registers[9][18] ;
 wire \core_pipeline.pipeline_registers.registers[9][19] ;
 wire \core_pipeline.pipeline_registers.registers[9][1] ;
 wire \core_pipeline.pipeline_registers.registers[9][20] ;
 wire \core_pipeline.pipeline_registers.registers[9][21] ;
 wire \core_pipeline.pipeline_registers.registers[9][22] ;
 wire \core_pipeline.pipeline_registers.registers[9][23] ;
 wire \core_pipeline.pipeline_registers.registers[9][24] ;
 wire \core_pipeline.pipeline_registers.registers[9][25] ;
 wire \core_pipeline.pipeline_registers.registers[9][26] ;
 wire \core_pipeline.pipeline_registers.registers[9][27] ;
 wire \core_pipeline.pipeline_registers.registers[9][28] ;
 wire \core_pipeline.pipeline_registers.registers[9][29] ;
 wire \core_pipeline.pipeline_registers.registers[9][2] ;
 wire \core_pipeline.pipeline_registers.registers[9][30] ;
 wire \core_pipeline.pipeline_registers.registers[9][31] ;
 wire \core_pipeline.pipeline_registers.registers[9][3] ;
 wire \core_pipeline.pipeline_registers.registers[9][4] ;
 wire \core_pipeline.pipeline_registers.registers[9][5] ;
 wire \core_pipeline.pipeline_registers.registers[9][6] ;
 wire \core_pipeline.pipeline_registers.registers[9][7] ;
 wire \core_pipeline.pipeline_registers.registers[9][8] ;
 wire \core_pipeline.pipeline_registers.registers[9][9] ;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net31;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net32;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net33;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net34;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net35;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net36;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net37;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net38;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net39;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net4;
 wire net40;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net41;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net42;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net43;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net44;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net45;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net46;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net47;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net48;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net49;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net5;
 wire net50;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net51;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net52;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net53;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net54;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net55;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net56;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net57;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net58;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net59;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net6;
 wire net60;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net61;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net62;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net63;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net64;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net65;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;

 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(_03749_));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(_05877_));
 sky130_fd_sc_hd__diode_2 ANTENNA_100 (.DIODE(\core_busio.mem_address[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_101 (.DIODE(\core_busio.mem_address[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_102 (.DIODE(\core_pipeline.csr_to_fetch_trap_vector[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_103 (.DIODE(\core_pipeline.decode_to_execute_csr_data[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_104 (.DIODE(\core_pipeline.decode_to_execute_csr_data[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_105 (.DIODE(\core_pipeline.memory_to_writeback_alu_data[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_106 (.DIODE(\core_pipeline.memory_to_writeback_alu_data[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_107 (.DIODE(\core_pipeline.pipeline_execute.ex_alu.result_sll[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_108 (.DIODE(\core_pipeline.pipeline_fetch.pc[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_109 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(_05885_));
 sky130_fd_sc_hd__diode_2 ANTENNA_110 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_111 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_112 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_113 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA_114 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_115 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA_116 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA_117 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA_118 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_119 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(_05925_));
 sky130_fd_sc_hd__diode_2 ANTENNA_120 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA_121 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA_122 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_123 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA_124 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA_125 (.DIODE(net521));
 sky130_fd_sc_hd__diode_2 ANTENNA_126 (.DIODE(net569));
 sky130_fd_sc_hd__diode_2 ANTENNA_127 (.DIODE(net578));
 sky130_fd_sc_hd__diode_2 ANTENNA_128 (.DIODE(net578));
 sky130_fd_sc_hd__diode_2 ANTENNA_129 (.DIODE(net581));
 sky130_fd_sc_hd__diode_2 ANTENNA_13 (.DIODE(_05965_));
 sky130_fd_sc_hd__diode_2 ANTENNA_130 (.DIODE(\core_pipeline.memory_to_writeback_alu_data[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_131 (.DIODE(\core_pipeline.memory_to_writeback_alu_data[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_132 (.DIODE(\core_pipeline.pipeline_fetch.pc[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_133 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_134 (.DIODE(\core_pipeline.pipeline_fetch.pc[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_14 (.DIODE(_05965_));
 sky130_fd_sc_hd__diode_2 ANTENNA_15 (.DIODE(_06626_));
 sky130_fd_sc_hd__diode_2 ANTENNA_16 (.DIODE(\core_busio.mem_address[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_17 (.DIODE(\core_busio.mem_address[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_18 (.DIODE(\core_busio.mem_address[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_19 (.DIODE(\core_busio.mem_address[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(_03866_));
 sky130_fd_sc_hd__diode_2 ANTENNA_20 (.DIODE(\core_pipeline.decode_to_csr_read_address[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_21 (.DIODE(\core_pipeline.decode_to_execute_csr_data[19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_22 (.DIODE(\core_pipeline.decode_to_execute_csr_data[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_23 (.DIODE(\core_pipeline.decode_to_execute_csr_data[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_24 (.DIODE(\core_pipeline.decode_to_execute_pc[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_25 (.DIODE(\core_pipeline.execute_to_memory_csr_data[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_26 (.DIODE(\core_pipeline.memory_to_writeback_alu_data[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_27 (.DIODE(\core_pipeline.memory_to_writeback_alu_data[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_28 (.DIODE(\core_pipeline.memory_to_writeback_alu_data[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_29 (.DIODE(\core_pipeline.memory_to_writeback_alu_data[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(_04828_));
 sky130_fd_sc_hd__diode_2 ANTENNA_30 (.DIODE(\core_pipeline.memory_to_writeback_alu_data[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_31 (.DIODE(\core_pipeline.memory_to_writeback_alu_data[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_32 (.DIODE(\core_pipeline.memory_to_writeback_alu_data[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_33 (.DIODE(\core_pipeline.memory_to_writeback_alu_data[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_34 (.DIODE(\core_pipeline.memory_to_writeback_alu_data[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_35 (.DIODE(\core_pipeline.memory_to_writeback_alu_data[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_36 (.DIODE(\core_pipeline.pipeline_execute.ex_alu.result_sll[19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_37 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA_38 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA_39 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(_04853_));
 sky130_fd_sc_hd__diode_2 ANTENNA_40 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA_41 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_42 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_43 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA_44 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_45 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA_46 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_47 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_48 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_49 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(_04901_));
 sky130_fd_sc_hd__diode_2 ANTENNA_50 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA_51 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_52 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA_53 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA_54 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA_55 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA_56 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA_57 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA_58 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA_59 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(_04901_));
 sky130_fd_sc_hd__diode_2 ANTENNA_60 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA_61 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA_62 (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA_63 (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA_64 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA_65 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA_66 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA_67 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_68 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_69 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(_04958_));
 sky130_fd_sc_hd__diode_2 ANTENNA_70 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_71 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA_72 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_73 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA_74 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_75 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_76 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA_77 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_78 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_79 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(_05022_));
 sky130_fd_sc_hd__diode_2 ANTENNA_80 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA_81 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA_82 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_83 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA_84 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_85 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA_86 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA_87 (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA_88 (.DIODE(net569));
 sky130_fd_sc_hd__diode_2 ANTENNA_89 (.DIODE(_03674_));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(_05102_));
 sky130_fd_sc_hd__diode_2 ANTENNA_90 (.DIODE(_03786_));
 sky130_fd_sc_hd__diode_2 ANTENNA_91 (.DIODE(_04618_));
 sky130_fd_sc_hd__diode_2 ANTENNA_92 (.DIODE(_04694_));
 sky130_fd_sc_hd__diode_2 ANTENNA_93 (.DIODE(_04694_));
 sky130_fd_sc_hd__diode_2 ANTENNA_94 (.DIODE(_04810_));
 sky130_fd_sc_hd__diode_2 ANTENNA_95 (.DIODE(_04810_));
 sky130_fd_sc_hd__diode_2 ANTENNA_96 (.DIODE(_05042_));
 sky130_fd_sc_hd__diode_2 ANTENNA_97 (.DIODE(_05753_));
 sky130_fd_sc_hd__diode_2 ANTENNA_98 (.DIODE(_05885_));
 sky130_fd_sc_hd__diode_2 ANTENNA_99 (.DIODE(\core_busio.mem_address[22] ));
 sky130_fd_sc_hd__decap_3 FILLER_0_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1014 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1034 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1058 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1089 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1115 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_628 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_790 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_880 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_908 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_931 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_966 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1019 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_1059 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1072 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_210 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_286 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_487 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_543 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_578 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_850 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_890 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_911 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_938 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1006 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_1113 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_255 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_33 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_366 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_583 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_685 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_774 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_798 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_807 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_822 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_855 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_912 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_938 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_964 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_976 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_984 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1018 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1055 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1067 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_1115 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_226 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_48 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_762 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_843 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_936 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_948 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_960 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_992 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1020 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1032 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1044 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_1056 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_1113 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_378 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_600 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_684 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_704 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_740 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_859 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_883 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_908 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_942 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_973 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_986 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_994 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1019 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_1028 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1105 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_275 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_302 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_384 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_404 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_443 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_512 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_616 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_674 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_719 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_836 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_888 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_92 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_944 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_952 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_990 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_1039 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1046 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_1058 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_1113 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_187 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_272 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_356 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_527 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_603 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_668 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_747 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_812 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_878 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_931 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_944 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_984 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_1010 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_1023 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1048 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1072 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_484 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_504 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_674 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_743 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_775 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_788 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_843 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_855 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_889 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_944 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_955 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_978 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_989 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_1113 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_202 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_572 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_666 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_761 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_873 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_882 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_907 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_915 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_928 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_964 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_986 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_994 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1000 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_1012 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_1024 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1042 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1054 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1066 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1078 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_438 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_544 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_604 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_836 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_844 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_889 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_909 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_934 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_956 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_988 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_1025 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1046 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_1058 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_1113 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_308 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_408 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_590 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_636 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_684 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_705 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_759 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_782 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_801 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_836 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_906 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_914 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_961 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_978 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_986 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_996 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1011 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1055 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1067 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1079 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_190 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_212 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_329 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_624 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_788 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_886 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_943 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_956 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_993 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_1010 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1018 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_1115 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_112 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_324 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_437 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_64 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_728 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_776 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_786 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_874 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_889 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_910 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_930 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_938 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_958 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_979 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_991 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_999 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_1005 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_1016 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1036 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1048 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_1113 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_415 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_572 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_600 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_803 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_823 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_838 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_874 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_90 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_907 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_934 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_938 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_967 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_1008 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1012 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_1032 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1073 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1105 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_120 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_427 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_494 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_728 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_848 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_854 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_932 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_957 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_970 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_977 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_988 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1019 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1031 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1043 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1063 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1071 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1075 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1087 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1099 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_1111 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_231 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_439 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_593 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_700 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_760 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_855 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_871 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_917 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_937 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_974 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_98 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_986 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1000 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1012 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1024 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_171 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_270 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_383 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_556 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_60 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_627 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_684 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_719 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_744 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_787 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_798 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_809 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_860 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_891 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_903 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_911 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_986 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1027 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1089 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_1113 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_124 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_144 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_252 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_420 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_815 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_822 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_859 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_877 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_906 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_930 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_975 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_991 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_999 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_1005 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_1027 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1055 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1067 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_136 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_282 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_380 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_551 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_572 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_616 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_675 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_730 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_788 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_810 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_834 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_843 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_883 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_907 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_916 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_956 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_976 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_985 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1007 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_1046 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1079 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1091 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_1103 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_1109 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_1115 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_140 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_200 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_238 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_352 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_423 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_570 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_684 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_762 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_838 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_848 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_86 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_872 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_915 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_926 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_930 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_934 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_978 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_990 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1002 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1008 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1055 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_1072 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_1080 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_176 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_451 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_542 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_570 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_606 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_775 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_788 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_79 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_804 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_830 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_842 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_885 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_902 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_947 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_968 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_1004 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_1032 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1036 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_1083 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1103 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_1115 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_238 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_408 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_644 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_696 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_733 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_759 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_772 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_801 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_816 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_850 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_858 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_884 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_916 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_935 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_958 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_966 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_992 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_1005 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1024 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1115 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_13 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_25 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_260 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_703 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_716 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_740 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_764 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_782 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_812 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_864 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_884 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_903 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_932 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_944 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_1002 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1006 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1014 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1020 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1024 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_1056 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1064 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_1082 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_329 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_440 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_542 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_575 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_688 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_734 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_768 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_780 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_786 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_828 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_833 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_845 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_903 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_973 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_990 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_1020 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1029 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1044 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_1075 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1083 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1103 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1115 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_143 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_407 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_42 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_455 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_500 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_552 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_604 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_762 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_796 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_808 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_828 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_832 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_859 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_874 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_906 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_918 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_928 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_936 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_958 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_966 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_975 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_990 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_1002 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1006 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1046 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_1058 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1062 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_1083 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_159 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_275 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_338 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_439 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_452 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_46 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_495 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_582 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_619 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_739 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_766 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_824 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_844 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_852 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_886 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_906 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_910 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_935 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_957 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_966 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_1027 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_1036 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_1047 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_1075 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1097 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_1109 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_42 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_440 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_46 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_594 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_647 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_668 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_807 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_884 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_927 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_978 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_997 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_1000 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1024 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1061 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_115 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_179 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_215 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_283 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_400 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_46 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_516 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_67 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_675 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_683 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_842 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_880 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_888 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_907 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_937 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_944 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_968 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1027 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_1036 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_1056 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_1081 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1092 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_1104 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_1109 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_1115 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_124 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_367 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_499 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_526 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_647 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_664 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_702 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_758 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_820 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_864 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_876 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_895 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_911 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_918 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_926 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_970 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_982 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1003 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1024 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_103 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1045 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_1070 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_219 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_231 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_380 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_434 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_454 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_560 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_635 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_651 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_72 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_731 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_768 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_804 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_858 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_866 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_886 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_898 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_907 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_918 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_939 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_954 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1006 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_1029 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1041 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_1061 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_1065 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_148 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_18 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_466 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_646 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_704 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_8 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_815 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_832 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_861 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_874 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_894 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_914 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_926 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_962 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_974 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_978 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_983 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1013 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1046 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1053 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1066 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1078 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1082 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_176 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_280 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_378 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_600 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_72 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_754 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_787 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_800 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_832 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_836 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_846 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_888 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_896 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_900 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_946 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_968 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_978 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1006 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_1030 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_1053 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1103 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1115 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_476 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_534 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_572 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_592 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_751 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_804 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_810 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_850 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_882 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_915 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_922 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_964 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_972 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_980 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_988 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1001 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_1025 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_1033 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1059 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1071 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_336 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_493 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_510 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_624 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_656 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_697 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_810 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_850 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_882 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_906 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_916 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_937 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_947 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_955 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_964 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_993 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_1011 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1019 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_1027 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_1034 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1067 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_1075 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_387 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_659 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_667 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_712 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_754 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_795 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_850 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_879 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_891 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_899 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_943 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_970 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_977 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_992 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_1020 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_1028 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1039 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_107 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_1073 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1096 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_1108 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1116 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_316 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_372 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_544 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_654 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_685 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_750 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_76 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_762 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_816 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_837 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_850 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_863 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_874 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_88 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_894 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_911 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_972 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1005 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1109 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1115 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_176 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_244 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_437 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_450 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_620 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_712 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_724 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_807 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_844 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_848 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_932 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_938 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_946 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_954 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_958 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_985 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_1000 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_1027 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1039 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1075 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1087 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_17 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_196 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_556 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_578 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_632 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_650 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_740 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_859 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_878 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_907 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_928 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_950 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_967 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1000 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_1012 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_104 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_1042 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_1050 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_1077 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1086 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_1115 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_159 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_537 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_675 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_688 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_719 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_822 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_834 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_844 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_856 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_894 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_915 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_960 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_964 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_974 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_986 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_992 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_1005 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_1040 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1055 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1062 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1071 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1089 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_1113 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_118 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_132 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_32 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_515 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_570 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_598 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_628 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_637 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_664 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_739 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_747 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_817 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_850 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_871 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_880 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_903 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_923 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_968 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_975 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_985 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_997 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_1004 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1010 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_1018 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_1056 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_1064 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_1088 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_235 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_269 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_331 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_385 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_452 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_48 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_518 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_676 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_768 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_808 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_937 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_1006 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_1029 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_1071 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_1079 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1098 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1110 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1116 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_124 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_358 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_422 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_459 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_496 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_527 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_668 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_806 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_851 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_859 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_866 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_874 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_881 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_890 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_918 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_929 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_962 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_1008 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1013 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1026 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1046 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_1061 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1070 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1074 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1083 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_116 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_219 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_339 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_380 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_453 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_470 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_544 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_619 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_675 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_766 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_781 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_852 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_892 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_904 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_943 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_956 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_973 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_991 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_1002 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_1018 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_1047 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_1055 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_1072 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_1085 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_1095 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_1103 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_1109 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_1115 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_124 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_160 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_30 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_594 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_740 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_751 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_759 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_806 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_838 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_851 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_870 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_930 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_971 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1006 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_1032 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1058 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_1113 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_266 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_532 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_598 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_634 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_644 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_740 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_758 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_766 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_820 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_832 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_849 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_860 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_884 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_918 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_926 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_100 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_1012 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_1061 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_1078 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1111 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_544 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_618 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_659 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_672 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_681 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_775 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_808 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_836 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_856 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_888 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_902 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_938 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_990 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_994 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_1002 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_102 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_1023 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_1055 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_1084 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_1109 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_188 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_212 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_216 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_254 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_40 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_528 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_536 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_630 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_687 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_703 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_763 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_778 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_812 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_832 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_851 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_878 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_906 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_912 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_929 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_94 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_963 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_970 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_990 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1019 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_1048 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_1060 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1064 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_1102 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_1110 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1116 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_271 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_448 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_498 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_544 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_550 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_600 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_636 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_722 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_754 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_810 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_827 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_901 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_952 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_963 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_978 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_995 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1027 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_1047 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_1074 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_1081 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_120 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_144 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_236 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_243 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_588 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_650 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_663 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_748 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_822 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_834 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_84 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_892 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_950 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_971 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_980 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_1018 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_1044 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_1068 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_1080 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_263 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_38 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_607 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_768 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_780 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_786 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_796 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_846 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_883 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_896 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_962 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_987 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_999 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_1020 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_1031 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_1047 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_1071 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_1094 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_1110 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1116 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_183 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_347 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_375 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_471 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_576 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_596 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_656 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_684 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_704 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_836 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_868 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_872 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_939 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_950 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_992 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_1015 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_1023 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_1055 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_1070 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_154 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_176 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_268 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_290 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_495 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_506 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_548 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_565 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_635 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_688 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_787 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_830 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_898 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_944 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_952 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_956 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_968 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_992 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_998 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_1032 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_1103 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_1115 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_140 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_231 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_325 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_420 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_691 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_848 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_854 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_915 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_946 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_971 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_990 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_1002 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1024 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1067 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_1088 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1105 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_268 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_379 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_450 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_551 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_672 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_724 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_830 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_843 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_902 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_922 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_962 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_1020 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1028 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_1036 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_1048 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1111 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_22 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_243 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_354 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_471 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_540 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_588 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_628 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_708 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_747 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_884 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_973 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_999 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1011 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1024 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1073 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_324 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_380 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_63 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_665 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_712 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_723 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_747 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_775 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_808 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_819 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_831 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_848 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_882 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_907 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_943 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_956 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_991 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_1002 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1049 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_1061 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_146 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_339 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_375 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_508 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_564 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_595 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_72 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_844 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_856 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_864 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_891 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_898 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_904 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_934 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_947 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1027 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1039 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1059 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1075 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1092 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1104 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1116 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_267 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_372 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_498 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_578 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_588 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_648 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_706 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_758 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_852 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_927 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_962 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_984 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_995 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_1002 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_1013 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_1046 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_1071 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_1081 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1098 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1110 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1116 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_275 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_292 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_38 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_450 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_552 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_599 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_619 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_778 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_786 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_831 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_843 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_851 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_896 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_904 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_922 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_944 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_956 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_965 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_994 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_1027 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_1039 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_1062 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1087 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1099 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_243 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_420 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_578 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_595 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_610 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_706 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_754 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_846 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_873 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_930 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_975 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_985 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1019 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1055 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_1067 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_1077 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_1088 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_116 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_271 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_339 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_407 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_448 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_540 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_596 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_60 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_696 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_723 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_761 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_774 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_810 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_830 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_847 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_866 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_884 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_918 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_935 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_950 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_956 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_964 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_1006 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_1057 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1063 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1071 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1092 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_1104 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_1115 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_263 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_274 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_303 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_357 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_364 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_646 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_742 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_796 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_814 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_854 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_862 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_871 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_895 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_912 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_924 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_960 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_967 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_1018 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1048 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_1066 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_1086 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_528 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_59 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_626 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_636 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_676 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_684 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_694 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_730 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_742 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_788 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_834 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_838 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_842 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_885 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_902 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_943 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_955 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1033 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1043 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_1071 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1079 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1103 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_1115 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_254 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_263 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_579 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_608 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_704 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_846 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_850 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_863 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_87 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_902 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_908 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_928 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_962 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_969 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_973 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_990 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1006 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_1018 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_1055 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1071 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_184 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_320 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_338 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_519 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_555 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_602 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_658 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_675 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_731 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_744 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_781 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_847 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_904 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_943 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_963 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_986 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_998 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_1027 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_1039 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_1050 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1096 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_1108 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1116 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_243 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_257 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_762 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_798 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_871 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_880 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_916 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_931 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_944 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_968 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_988 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1040 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1044 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1113 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_500 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_744 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_756 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_760 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_794 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_864 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_868 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_908 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_919 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_927 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_939 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_949 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_986 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_1006 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_1059 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_1070 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1105 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_273 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_280 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_288 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_496 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_508 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_620 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_675 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_712 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_754 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_789 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_800 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_823 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_851 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_883 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_892 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_902 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_943 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_957 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_965 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_992 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_1018 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_1026 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1044 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1071 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1083 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1095 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_1107 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_1115 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_179 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_376 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_411 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_486 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_710 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_720 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_778 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_799 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_810 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_816 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_861 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_874 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_920 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_932 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_963 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_967 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_975 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_987 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_995 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_1003 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_1027 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1053 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_1062 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_1115 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_112 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_147 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_327 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_504 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_552 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_658 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_692 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_740 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_768 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_788 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_792 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_822 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_850 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_862 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_904 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_992 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_101 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_1018 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1024 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1034 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_1046 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1052 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_1060 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1081 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_319 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_354 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_375 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_484 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_660 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_747 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_759 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_905 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_930 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_963 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_973 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_995 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_1007 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_1015 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_1046 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1050 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_1059 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1080 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_158 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_288 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_370 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_487 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_528 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_676 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_712 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_802 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_875 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_883 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_894 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_902 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_921 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_937 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_948 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_956 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_990 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1024 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1044 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_1062 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1113 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_124 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_247 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_413 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_523 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_544 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_760 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_794 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_806 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_814 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_872 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_876 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_902 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_906 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_916 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_926 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_930 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_936 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_942 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_964 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_976 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_988 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_995 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_1006 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_1016 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_1024 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_1043 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1051 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1080 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_435 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_455 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_744 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_768 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_793 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_804 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_828 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_840 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_854 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_903 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_978 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_1018 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_1026 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_1039 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1071 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1083 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1095 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_1107 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_1115 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_123 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_134 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_247 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_352 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_378 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_412 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_781 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_791 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_832 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_874 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_878 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_883 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_902 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_926 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_948 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_968 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_982 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_994 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1075 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_224 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_244 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_438 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_487 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_542 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_563 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_730 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_754 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_782 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_786 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_826 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_878 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_956 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1007 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1022 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_1034 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1038 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1071 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1083 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1095 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_1107 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_1115 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_199 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_357 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_422 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_656 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_752 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_776 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_834 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_854 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_861 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_868 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_880 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_90 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_903 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_926 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_932 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_940 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_962 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_970 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1004 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1062 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1086 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1105 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_264 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_284 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_430 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_607 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_676 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_730 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_750 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_773 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_786 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_798 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_847 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_860 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_881 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_891 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_899 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_911 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_956 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_968 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_978 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_990 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_994 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_1004 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_1012 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1018 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_1027 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1034 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_1067 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_1088 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1115 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_156 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_213 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_238 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_451 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_470 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_496 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_551 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_622 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_768 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_830 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_894 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_939 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_950 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_956 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_992 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_1002 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_1036 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1074 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1086 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1098 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_1110 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1116 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_484 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_523 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_610 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_646 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_691 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_758 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_804 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_864 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_875 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_915 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_973 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_995 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_1067 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1105 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_126 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_712 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_731 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_748 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_791 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_830 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_839 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_880 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_904 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_922 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_957 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_978 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_989 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1025 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1031 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_1043 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_1056 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_1113 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_202 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_366 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_532 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_628 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_684 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_763 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_767 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_803 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_909 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_927 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_939 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_962 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_973 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_988 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_998 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1006 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_1018 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_228 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_275 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_506 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_600 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_604 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_719 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_742 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_811 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_834 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_891 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_945 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_1018 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1026 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_1032 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_1043 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_1113 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_158 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_666 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_692 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_748 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_816 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_838 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_859 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_868 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_876 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_916 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_926 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_935 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_946 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_960 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_982 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1006 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1018 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_1027 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_1034 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1069 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_1081 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_507 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_520 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_582 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_628 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_775 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_810 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_826 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_860 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_923 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_931 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_989 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_1049 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1089 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_1109 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_1115 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_16 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_40 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_571 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_637 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_684 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_690 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_702 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_747 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_839 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_874 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_908 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_912 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_957 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_974 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_998 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1015 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1046 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1058 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1070 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_1082 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_338 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_570 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_710 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_768 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_772 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_810 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_833 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_858 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_874 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_898 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_944 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_964 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_992 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_1000 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1028 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1040 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1052 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_1113 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_476 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_522 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_684 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_715 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_807 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_856 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_876 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_906 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_914 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_935 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_962 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_970 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_978 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_990 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1083 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1095 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_1107 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1115 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_126 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_257 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_627 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_649 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_724 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_747 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_758 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_766 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_862 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_871 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_927 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_971 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_980 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_988 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_996 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_549 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_786 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_830 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_878 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_884 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_947 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_958 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1007 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1023 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1047 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_1113 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_303 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_590 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_628 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_641 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_691 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_812 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_821 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_832 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_863 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_883 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_912 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_949 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_976 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_982 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1003 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_1012 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_1032 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_352 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_791 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_892 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_904 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_943 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_1016 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1024 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1036 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1048 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_1113 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_584 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_628 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_646 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_684 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_704 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_735 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_745 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_812 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_818 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_861 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_870 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_878 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_915 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_973 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_995 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_452 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_472 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_624 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_663 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_826 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_834 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_900 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_912 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_935 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1014 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1026 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1038 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_1104 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_1115 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_482 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_648 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_783 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_807 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_878 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_884 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_919 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_939 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1011 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_464 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_494 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_607 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_632 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_684 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_712 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_781 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_864 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_873 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_914 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_939 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_956 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_968 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_999 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_1113 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_350 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_588 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_628 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_644 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_668 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_802 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_814 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_823 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_856 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_867 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_874 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_895 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_911 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_934 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_989 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_1015 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_1044 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_1085 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_1099 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_1103 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_1109 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_1115 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_239 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_628 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_763 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_767 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_792 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_876 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1007 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1019 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1070 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_180 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_460 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_49 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_62 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_712 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_736 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_829 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_848 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_903 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_954 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_978 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_996 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1004 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1027 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1039 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1109 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1115 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_13 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_426 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_608 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_712 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_810 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_820 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_870 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_961 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1089 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1115 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_415 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_646 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_703 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_760 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_873 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_894 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_919 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_931 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1016 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1048 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1052 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_455 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_510 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_551 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_568 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_631 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_763 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_792 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_820 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_906 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_943 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_992 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1071 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1083 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1095 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_1107 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1115 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_466 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_593 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_646 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_747 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_783 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_791 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_808 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_816 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_872 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_915 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_948 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_983 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1010 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_1030 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1064 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1105 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_519 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_712 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_768 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_808 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_832 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_882 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_903 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_936 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_944 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_956 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_976 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1040 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1076 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1088 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1100 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1112 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1116 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_186 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_372 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_524 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_592 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_703 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_744 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_756 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_822 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_832 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_847 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_884 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_910 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_920 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_930 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_973 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_986 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_999 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_1004 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1010 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1032 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1053 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1070 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_439 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_544 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_556 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_605 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_649 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_680 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_777 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_834 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_846 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_866 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_900 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_922 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_938 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_960 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_979 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_1020 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1040 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1052 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1074 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1086 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1098 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1110 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1116 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_351 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_46 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_511 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_639 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_759 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_834 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_857 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_931 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_984 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_997 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1055 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1067 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1079 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1109 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_114 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_264 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_283 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_680 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_790 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_832 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_844 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_899 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_936 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_960 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_968 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_999 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1020 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1058 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1113 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_255 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_471 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_482 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_523 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_711 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_752 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_771 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_796 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_815 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_864 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_868 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_910 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_914 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_931 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_964 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_970 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_997 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1034 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1045 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1062 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1074 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1086 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_115 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_172 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_454 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_488 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_606 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_656 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_718 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_731 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_739 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_766 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_807 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_817 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_834 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_842 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_883 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_896 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_907 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_947 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_960 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_968 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_994 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1044 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1113 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_366 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_424 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_703 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_716 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_748 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_852 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_880 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_915 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_932 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_970 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_982 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_992 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_565 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_808 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_865 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_888 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_908 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_943 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_955 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_967 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1001 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1059 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1071 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_112 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_160 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_25 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_33 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_495 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_640 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_664 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_733 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_826 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_844 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_852 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_860 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_904 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_916 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_942 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_954 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_989 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1043 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1113 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_30 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_467 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_525 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_579 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_638 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_704 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_831 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_852 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_864 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_923 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_99 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1050 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1074 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1086 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_627 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_740 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_775 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_788 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_824 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_850 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_904 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_943 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_956 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_999 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1016 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1041 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1113 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_579 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_691 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_745 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_859 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_86 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_915 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_939 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_965 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_982 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1019 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1023 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1066 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1078 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1115 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_244 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_272 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_641 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_787 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_800 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_832 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_849 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_936 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_942 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_976 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_994 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_998 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_1000 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1013 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_1038 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1048 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1089 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1113 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_17 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_704 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_817 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_856 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_968 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_991 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1004 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1010 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1044 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1072 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_358 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_507 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_524 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_554 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_71 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_788 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_880 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_893 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_936 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_942 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_952 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_962 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1004 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_1036 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1044 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1088 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1100 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1112 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1116 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_303 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_406 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_479 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_590 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_668 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_716 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_791 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_801 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_859 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_892 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_921 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1003 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_1048 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1056 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1078 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_382 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_632 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_665 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_724 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_764 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_772 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_803 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_823 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_833 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_854 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_864 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_920 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_959 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_976 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_1000 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1048 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1098 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1110 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1116 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_330 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_47 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_496 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_71 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_792 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_800 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_859 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_872 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_905 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_918 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_930 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_974 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_978 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_99 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1113 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_460 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_523 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_590 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_649 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_716 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_760 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_814 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_934 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_938 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1024 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1053 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_13 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_170 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_247 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_378 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_435 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_470 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_564 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_607 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_651 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_684 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_721 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_831 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_864 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_898 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_936 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_955 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_978 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1007 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1046 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1063 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1071 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1081 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1109 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1115 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_355 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_411 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_462 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_655 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_695 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_707 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_722 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_863 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_875 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_906 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_914 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_932 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_964 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_976 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_988 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1011 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1059 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1075 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1105 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_226 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_269 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_322 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_339 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_448 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_554 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_634 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_656 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_668 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_832 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_911 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_943 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1007 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1036 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1042 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1088 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1100 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1112 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1116 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_484 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_497 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_532 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_644 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_664 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_695 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_708 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_790 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_817 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_854 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_87 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_874 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_908 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_912 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_960 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_966 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_988 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1003 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1020 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_1034 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1053 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1078 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1086 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_1093 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_11 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1111 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_270 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_295 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_490 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_663 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_675 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_788 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_856 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_892 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_905 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_936 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_942 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_959 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_999 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1020 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_1032 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_1040 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1083 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1095 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_1107 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1115 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_131 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_320 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_523 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_647 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_714 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_753 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_838 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_871 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_907 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_915 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_927 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_964 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_968 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_990 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_1008 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1016 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1023 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1049 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1072 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_163 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_183 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_507 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_524 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_636 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_680 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_712 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_875 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_908 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_943 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_955 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_992 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_998 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1032 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1044 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_1056 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1113 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_136 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_476 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_644 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_693 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_705 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_722 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_782 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_812 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_816 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_836 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_864 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_906 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_918 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_926 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_964 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_976 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_995 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_1000 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_1008 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1032 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1061 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1105 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_172 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_434 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_607 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_721 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_75 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_835 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_856 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_880 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_884 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_906 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_910 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_964 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_968 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1032 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1083 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_1095 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1115 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_129 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_299 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_348 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_466 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_574 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_610 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_762 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_807 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_815 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_84 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_864 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_876 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_894 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_905 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_962 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_551 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_628 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_694 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_768 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_856 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_875 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_922 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_952 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_964 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1055 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1075 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1088 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_216 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_383 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_434 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_484 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_504 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_556 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_616 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_628 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_638 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_692 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_776 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_844 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_864 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_945 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1050 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1088 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1113 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_179 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_196 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_292 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_715 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_762 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_920 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_926 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_964 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_974 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_986 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_994 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_1005 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1020 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1070 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1081 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_182 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_383 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_798 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_836 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_848 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_880 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_906 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_993 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1027 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1046 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1059 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1083 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1103 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1115 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_668 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_754 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_821 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_856 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_878 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_915 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_971 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_988 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1014 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1070 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_215 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_324 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_378 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_444 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_608 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_626 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_634 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_663 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_728 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_775 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_788 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_796 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_806 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_839 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_907 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_932 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_956 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_993 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1027 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1047 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1083 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1095 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_1107 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1115 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_348 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_514 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_534 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_554 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_636 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_759 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_809 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_851 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_855 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_876 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_915 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_928 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_964 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_970 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1005 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1018 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1068 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1088 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_1115 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_45 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_486 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_62 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_656 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_712 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_787 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_836 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_842 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_867 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_902 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_936 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_940 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_992 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_1020 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1028 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1076 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1088 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1100 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1112 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1116 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_142 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_422 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_574 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_635 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_648 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_702 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_756 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_794 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_859 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_880 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_928 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_961 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_999 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1018 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1048 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1072 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_284 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_327 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_544 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_675 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_796 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_880 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_902 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_952 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_962 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_988 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_997 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1020 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_1032 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_1040 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1052 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1089 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1113 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_299 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_355 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_471 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_479 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_554 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_75 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_758 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_794 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_894 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_912 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_935 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_951 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_968 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_1113 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_579 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_684 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_760 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_864 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_884 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_934 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_965 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1019 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1032 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1041 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1058 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1070 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1080 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_112 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_159 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_416 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_674 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_707 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_724 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_796 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_900 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_957 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_999 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1002 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1029 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1083 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1095 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1115 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_187 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_28 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_290 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_311 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_348 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_366 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_621 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_747 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_780 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_859 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_916 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_928 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_976 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_99 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1011 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_1060 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1068 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1079 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_330 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_339 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_386 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_448 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_575 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_663 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_710 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_767 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_787 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_880 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_899 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1018 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_1031 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_1042 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1063 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1069 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1086 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1098 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_1110 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1116 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_367 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_603 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_697 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_708 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_760 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_803 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_859 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_883 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_935 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_964 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_970 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1003 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1016 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_1028 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1049 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_1061 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1069 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_1086 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_1093 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1115 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_319 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_544 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_566 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_674 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_864 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_962 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_992 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_1020 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1028 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1038 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1050 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1087 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_1111 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_308 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_431 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_735 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_859 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_915 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_966 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1003 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1058 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1062 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_226 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_439 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_454 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_495 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_607 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_728 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_831 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_880 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_884 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_902 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_936 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_940 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_957 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_992 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_1002 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1039 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1043 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1060 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1088 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1100 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1112 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1116 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_515 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_579 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_682 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_726 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_756 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_839 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_935 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_964 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_972 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_990 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1044 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1048 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1080 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1093 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_112 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_339 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_356 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_571 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_60 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_723 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_733 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_798 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_920 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_944 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_964 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_999 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1042 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1075 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1087 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1099 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_1111 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_183 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_242 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_300 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_372 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_590 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_610 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_718 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_759 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_859 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_892 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_919 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_973 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_986 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_990 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_1000 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1013 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1105 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_163 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_394 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_784 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_832 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_864 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_900 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_912 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_952 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_964 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_968 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_978 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1004 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_1030 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1074 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_1086 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1105 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_440 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_495 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_640 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_672 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_720 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_763 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_780 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_786 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_943 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_955 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_992 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_1016 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1022 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1088 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_1100 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_1108 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1115 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_130 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_308 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_351 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_49 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_516 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_540 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_588 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_682 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_758 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_851 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_872 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_908 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_916 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_946 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_100 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_1008 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1016 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1034 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1059 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_1084 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1099 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_1111 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_327 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_378 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_456 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_495 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_506 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_512 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_544 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_621 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_67 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_752 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_836 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_846 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_866 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_988 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1006 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1038 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1083 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1103 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1115 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_126 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_412 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_492 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_52 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_583 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_690 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_707 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_742 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_859 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_872 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_908 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_951 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_976 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_986 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_1005 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1020 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1055 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1072 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1104 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1116 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_213 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_270 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_295 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_56 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_675 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_799 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_831 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_864 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_907 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_943 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_957 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_995 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1039 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1052 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1083 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1095 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_1107 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1115 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_294 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_532 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_682 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_707 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_760 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_880 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_934 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_971 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_988 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_994 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1012 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1024 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1048 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_1060 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1088 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_13 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_23 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_515 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_526 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_676 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_728 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_748 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_75 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_779 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_843 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_876 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_896 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_934 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_944 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_954 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_991 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_1041 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1083 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1095 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_1107 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1115 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_467 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_47 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_556 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_637 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_648 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_702 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_836 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_84 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_870 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_890 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_935 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_960 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_964 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_985 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_1014 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_1081 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_380 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_516 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_787 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_899 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_92 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_936 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_940 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_978 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1042 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1076 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1088 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1102 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1115 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_47 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_480 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_526 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_596 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_744 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_754 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_834 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_866 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_870 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_905 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_950 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_983 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_1113 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_486 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_496 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_522 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_571 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_647 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_660 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_683 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_880 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_893 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_908 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_912 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_974 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_994 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1004 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_1017 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1088 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_154 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_210 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_230 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_280 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_298 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_443 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_460 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_616 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_831 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_906 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_941 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_964 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_968 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_992 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_1040 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_1088 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1096 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_1108 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1116 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_299 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_600 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_762 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_782 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_800 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_832 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_940 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_985 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_996 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_1015 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_1028 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_1048 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_1060 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_1068 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_107 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_1086 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_499 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_656 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_676 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_684 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_710 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_778 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_856 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_896 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_900 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_936 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_960 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_990 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_1006 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_1038 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_1058 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1078 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1102 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_1114 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_431 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_575 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_599 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_627 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_871 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_927 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_964 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_968 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_974 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_987 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_1044 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1052 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1071 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_428 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_490 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_64 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_675 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_739 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_768 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_788 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_936 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_940 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1004 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1027 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1062 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1071 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1088 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1100 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1112 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1116 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_243 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_411 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_588 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_650 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_692 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_751 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_766 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_814 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_859 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_892 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_92 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_921 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_934 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_950 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_984 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_1004 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1012 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_106 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1090 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1115 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_22 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_326 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_575 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_634 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_656 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_666 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_721 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_732 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_738 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_754 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_792 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_840 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_880 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_900 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_1027 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_1040 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_1088 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_1113 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_266 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_424 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_478 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_575 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_612 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_640 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_750 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_806 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_816 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_878 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_931 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_964 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_970 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_991 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_1066 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_1086 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_120 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_275 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_387 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_443 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_504 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_544 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_658 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_681 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_710 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_782 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_786 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_803 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_843 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_880 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_884 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_967 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_999 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_1004 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1087 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1099 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_1111 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_296 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_319 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_648 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_724 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_818 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_838 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_857 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_88 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_907 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_913 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_951 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_959 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_977 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1024 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_163 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_618 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_712 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_730 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_856 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_865 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_947 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_1004 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1048 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_1060 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1068 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1078 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1105 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_275 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_496 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_504 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_52 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_624 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_675 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_732 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_843 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_891 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_979 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_987 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1002 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_1030 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1042 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1074 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1096 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_1108 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1116 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_244 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_456 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_482 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_516 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_805 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_826 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_880 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_911 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_930 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1003 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1015 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1027 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1059 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1070 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_378 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_426 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_600 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_631 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_744 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_798 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_836 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_860 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_949 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_1032 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_1042 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1083 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1095 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_1107 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1115 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_351 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_431 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_480 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_655 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_702 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_79 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_810 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_814 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_846 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_866 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_886 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_927 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_978 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_998 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_1058 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_106 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_273 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_506 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_565 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_666 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_730 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_768 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_844 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_848 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_880 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_888 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_907 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_954 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_966 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_1076 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1115 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_410 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_426 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_500 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_666 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_691 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_708 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_722 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_735 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_752 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_783 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_821 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_846 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_850 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_878 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_915 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_936 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_940 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_964 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_976 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_988 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_1018 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1024 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1055 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_114 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_172 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_271 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_296 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_437 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_674 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_711 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_719 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_748 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_79 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_790 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_833 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_850 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_890 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_898 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_936 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_942 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_959 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1020 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_1032 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_1113 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_140 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_260 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_440 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_480 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_552 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_740 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_758 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_859 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_912 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_930 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_994 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1072 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_271 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_386 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_518 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_59 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_912 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_943 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_952 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_960 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_992 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_1030 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1083 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1095 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_1107 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_1115 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_245 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_487 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_494 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_532 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_636 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_740 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_760 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_796 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_852 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_876 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_884 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_908 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_974 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_982 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_999 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1002 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1027 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1113 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_599 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_647 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_684 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_749 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_803 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_815 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_871 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_920 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_950 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_977 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_194 ();
 sky130_fd_sc_hd__decap_3 PHY_195 ();
 sky130_fd_sc_hd__decap_3 PHY_196 ();
 sky130_fd_sc_hd__decap_3 PHY_197 ();
 sky130_fd_sc_hd__decap_3 PHY_198 ();
 sky130_fd_sc_hd__decap_3 PHY_199 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_200 ();
 sky130_fd_sc_hd__decap_3 PHY_201 ();
 sky130_fd_sc_hd__decap_3 PHY_202 ();
 sky130_fd_sc_hd__decap_3 PHY_203 ();
 sky130_fd_sc_hd__decap_3 PHY_204 ();
 sky130_fd_sc_hd__decap_3 PHY_205 ();
 sky130_fd_sc_hd__decap_3 PHY_206 ();
 sky130_fd_sc_hd__decap_3 PHY_207 ();
 sky130_fd_sc_hd__decap_3 PHY_208 ();
 sky130_fd_sc_hd__decap_3 PHY_209 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_210 ();
 sky130_fd_sc_hd__decap_3 PHY_211 ();
 sky130_fd_sc_hd__decap_3 PHY_212 ();
 sky130_fd_sc_hd__decap_3 PHY_213 ();
 sky130_fd_sc_hd__decap_3 PHY_214 ();
 sky130_fd_sc_hd__decap_3 PHY_215 ();
 sky130_fd_sc_hd__decap_3 PHY_216 ();
 sky130_fd_sc_hd__decap_3 PHY_217 ();
 sky130_fd_sc_hd__decap_3 PHY_218 ();
 sky130_fd_sc_hd__decap_3 PHY_219 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_220 ();
 sky130_fd_sc_hd__decap_3 PHY_221 ();
 sky130_fd_sc_hd__decap_3 PHY_222 ();
 sky130_fd_sc_hd__decap_3 PHY_223 ();
 sky130_fd_sc_hd__decap_3 PHY_224 ();
 sky130_fd_sc_hd__decap_3 PHY_225 ();
 sky130_fd_sc_hd__decap_3 PHY_226 ();
 sky130_fd_sc_hd__decap_3 PHY_227 ();
 sky130_fd_sc_hd__decap_3 PHY_228 ();
 sky130_fd_sc_hd__decap_3 PHY_229 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_230 ();
 sky130_fd_sc_hd__decap_3 PHY_231 ();
 sky130_fd_sc_hd__decap_3 PHY_232 ();
 sky130_fd_sc_hd__decap_3 PHY_233 ();
 sky130_fd_sc_hd__decap_3 PHY_234 ();
 sky130_fd_sc_hd__decap_3 PHY_235 ();
 sky130_fd_sc_hd__decap_3 PHY_236 ();
 sky130_fd_sc_hd__decap_3 PHY_237 ();
 sky130_fd_sc_hd__decap_3 PHY_238 ();
 sky130_fd_sc_hd__decap_3 PHY_239 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_240 ();
 sky130_fd_sc_hd__decap_3 PHY_241 ();
 sky130_fd_sc_hd__decap_3 PHY_242 ();
 sky130_fd_sc_hd__decap_3 PHY_243 ();
 sky130_fd_sc_hd__decap_3 PHY_244 ();
 sky130_fd_sc_hd__decap_3 PHY_245 ();
 sky130_fd_sc_hd__decap_3 PHY_246 ();
 sky130_fd_sc_hd__decap_3 PHY_247 ();
 sky130_fd_sc_hd__decap_3 PHY_248 ();
 sky130_fd_sc_hd__decap_3 PHY_249 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_250 ();
 sky130_fd_sc_hd__decap_3 PHY_251 ();
 sky130_fd_sc_hd__decap_3 PHY_252 ();
 sky130_fd_sc_hd__decap_3 PHY_253 ();
 sky130_fd_sc_hd__decap_3 PHY_254 ();
 sky130_fd_sc_hd__decap_3 PHY_255 ();
 sky130_fd_sc_hd__decap_3 PHY_256 ();
 sky130_fd_sc_hd__decap_3 PHY_257 ();
 sky130_fd_sc_hd__decap_3 PHY_258 ();
 sky130_fd_sc_hd__decap_3 PHY_259 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_260 ();
 sky130_fd_sc_hd__decap_3 PHY_261 ();
 sky130_fd_sc_hd__decap_3 PHY_262 ();
 sky130_fd_sc_hd__decap_3 PHY_263 ();
 sky130_fd_sc_hd__decap_3 PHY_264 ();
 sky130_fd_sc_hd__decap_3 PHY_265 ();
 sky130_fd_sc_hd__decap_3 PHY_266 ();
 sky130_fd_sc_hd__decap_3 PHY_267 ();
 sky130_fd_sc_hd__decap_3 PHY_268 ();
 sky130_fd_sc_hd__decap_3 PHY_269 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_270 ();
 sky130_fd_sc_hd__decap_3 PHY_271 ();
 sky130_fd_sc_hd__decap_3 PHY_272 ();
 sky130_fd_sc_hd__decap_3 PHY_273 ();
 sky130_fd_sc_hd__decap_3 PHY_274 ();
 sky130_fd_sc_hd__decap_3 PHY_275 ();
 sky130_fd_sc_hd__decap_3 PHY_276 ();
 sky130_fd_sc_hd__decap_3 PHY_277 ();
 sky130_fd_sc_hd__decap_3 PHY_278 ();
 sky130_fd_sc_hd__decap_3 PHY_279 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_280 ();
 sky130_fd_sc_hd__decap_3 PHY_281 ();
 sky130_fd_sc_hd__decap_3 PHY_282 ();
 sky130_fd_sc_hd__decap_3 PHY_283 ();
 sky130_fd_sc_hd__decap_3 PHY_284 ();
 sky130_fd_sc_hd__decap_3 PHY_285 ();
 sky130_fd_sc_hd__decap_3 PHY_286 ();
 sky130_fd_sc_hd__decap_3 PHY_287 ();
 sky130_fd_sc_hd__decap_3 PHY_288 ();
 sky130_fd_sc_hd__decap_3 PHY_289 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_290 ();
 sky130_fd_sc_hd__decap_3 PHY_291 ();
 sky130_fd_sc_hd__decap_3 PHY_292 ();
 sky130_fd_sc_hd__decap_3 PHY_293 ();
 sky130_fd_sc_hd__decap_3 PHY_294 ();
 sky130_fd_sc_hd__decap_3 PHY_295 ();
 sky130_fd_sc_hd__decap_3 PHY_296 ();
 sky130_fd_sc_hd__decap_3 PHY_297 ();
 sky130_fd_sc_hd__decap_3 PHY_298 ();
 sky130_fd_sc_hd__decap_3 PHY_299 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_300 ();
 sky130_fd_sc_hd__decap_3 PHY_301 ();
 sky130_fd_sc_hd__decap_3 PHY_302 ();
 sky130_fd_sc_hd__decap_3 PHY_303 ();
 sky130_fd_sc_hd__decap_3 PHY_304 ();
 sky130_fd_sc_hd__decap_3 PHY_305 ();
 sky130_fd_sc_hd__decap_3 PHY_306 ();
 sky130_fd_sc_hd__decap_3 PHY_307 ();
 sky130_fd_sc_hd__decap_3 PHY_308 ();
 sky130_fd_sc_hd__decap_3 PHY_309 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_310 ();
 sky130_fd_sc_hd__decap_3 PHY_311 ();
 sky130_fd_sc_hd__decap_3 PHY_312 ();
 sky130_fd_sc_hd__decap_3 PHY_313 ();
 sky130_fd_sc_hd__decap_3 PHY_314 ();
 sky130_fd_sc_hd__decap_3 PHY_315 ();
 sky130_fd_sc_hd__decap_3 PHY_316 ();
 sky130_fd_sc_hd__decap_3 PHY_317 ();
 sky130_fd_sc_hd__decap_3 PHY_318 ();
 sky130_fd_sc_hd__decap_3 PHY_319 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_320 ();
 sky130_fd_sc_hd__decap_3 PHY_321 ();
 sky130_fd_sc_hd__decap_3 PHY_322 ();
 sky130_fd_sc_hd__decap_3 PHY_323 ();
 sky130_fd_sc_hd__decap_3 PHY_324 ();
 sky130_fd_sc_hd__decap_3 PHY_325 ();
 sky130_fd_sc_hd__decap_3 PHY_326 ();
 sky130_fd_sc_hd__decap_3 PHY_327 ();
 sky130_fd_sc_hd__decap_3 PHY_328 ();
 sky130_fd_sc_hd__decap_3 PHY_329 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_330 ();
 sky130_fd_sc_hd__decap_3 PHY_331 ();
 sky130_fd_sc_hd__decap_3 PHY_332 ();
 sky130_fd_sc_hd__decap_3 PHY_333 ();
 sky130_fd_sc_hd__decap_3 PHY_334 ();
 sky130_fd_sc_hd__decap_3 PHY_335 ();
 sky130_fd_sc_hd__decap_3 PHY_336 ();
 sky130_fd_sc_hd__decap_3 PHY_337 ();
 sky130_fd_sc_hd__decap_3 PHY_338 ();
 sky130_fd_sc_hd__decap_3 PHY_339 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_340 ();
 sky130_fd_sc_hd__decap_3 PHY_341 ();
 sky130_fd_sc_hd__decap_3 PHY_342 ();
 sky130_fd_sc_hd__decap_3 PHY_343 ();
 sky130_fd_sc_hd__decap_3 PHY_344 ();
 sky130_fd_sc_hd__decap_3 PHY_345 ();
 sky130_fd_sc_hd__decap_3 PHY_346 ();
 sky130_fd_sc_hd__decap_3 PHY_347 ();
 sky130_fd_sc_hd__decap_3 PHY_348 ();
 sky130_fd_sc_hd__decap_3 PHY_349 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_350 ();
 sky130_fd_sc_hd__decap_3 PHY_351 ();
 sky130_fd_sc_hd__decap_3 PHY_352 ();
 sky130_fd_sc_hd__decap_3 PHY_353 ();
 sky130_fd_sc_hd__decap_3 PHY_354 ();
 sky130_fd_sc_hd__decap_3 PHY_355 ();
 sky130_fd_sc_hd__decap_3 PHY_356 ();
 sky130_fd_sc_hd__decap_3 PHY_357 ();
 sky130_fd_sc_hd__decap_3 PHY_358 ();
 sky130_fd_sc_hd__decap_3 PHY_359 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_360 ();
 sky130_fd_sc_hd__decap_3 PHY_361 ();
 sky130_fd_sc_hd__decap_3 PHY_362 ();
 sky130_fd_sc_hd__decap_3 PHY_363 ();
 sky130_fd_sc_hd__decap_3 PHY_364 ();
 sky130_fd_sc_hd__decap_3 PHY_365 ();
 sky130_fd_sc_hd__decap_3 PHY_366 ();
 sky130_fd_sc_hd__decap_3 PHY_367 ();
 sky130_fd_sc_hd__decap_3 PHY_368 ();
 sky130_fd_sc_hd__decap_3 PHY_369 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_370 ();
 sky130_fd_sc_hd__decap_3 PHY_371 ();
 sky130_fd_sc_hd__decap_3 PHY_372 ();
 sky130_fd_sc_hd__decap_3 PHY_373 ();
 sky130_fd_sc_hd__decap_3 PHY_374 ();
 sky130_fd_sc_hd__decap_3 PHY_375 ();
 sky130_fd_sc_hd__decap_3 PHY_376 ();
 sky130_fd_sc_hd__decap_3 PHY_377 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__inv_2 _06658_ (.A(\core_pipeline.pipeline_fetch.pc[2] ),
    .Y(_03312_));
 sky130_fd_sc_hd__inv_2 _06659_ (.A(\core_pipeline.fetch_to_decode_instruction[14] ),
    .Y(_03313_));
 sky130_fd_sc_hd__inv_2 _06660_ (.A(net505),
    .Y(_03314_));
 sky130_fd_sc_hd__inv_2 _06661_ (.A(\core_busio.mem_size[1] ),
    .Y(_03315_));
 sky130_fd_sc_hd__inv_2 _06662_ (.A(\core_busio.mem_size[0] ),
    .Y(_03316_));
 sky130_fd_sc_hd__inv_2 _06663_ (.A(\core_pipeline.decode_to_execute_rd_address[0] ),
    .Y(_03317_));
 sky130_fd_sc_hd__inv_2 _06664_ (.A(\core_pipeline.decode_to_execute_rd_address[3] ),
    .Y(_03318_));
 sky130_fd_sc_hd__inv_2 _06665_ (.A(\core_pipeline.decode_to_execute_rd_address[2] ),
    .Y(_03319_));
 sky130_fd_sc_hd__inv_2 _06666_ (.A(\core_pipeline.decode_to_execute_rd_address[4] ),
    .Y(_03320_));
 sky130_fd_sc_hd__inv_2 _06667_ (.A(\core_pipeline.fetch_to_decode_instruction[13] ),
    .Y(_03321_));
 sky130_fd_sc_hd__inv_2 _06668_ (.A(\core_pipeline.fetch_to_decode_instruction[5] ),
    .Y(_03322_));
 sky130_fd_sc_hd__inv_6 _06669_ (.A(net595),
    .Y(_03323_));
 sky130_fd_sc_hd__inv_2 _06670_ (.A(net579),
    .Y(_03324_));
 sky130_fd_sc_hd__inv_4 _06671_ (.A(net573),
    .Y(_03325_));
 sky130_fd_sc_hd__clkinv_4 _06672_ (.A(net567),
    .Y(_03326_));
 sky130_fd_sc_hd__inv_6 _06673_ (.A(net565),
    .Y(_03327_));
 sky130_fd_sc_hd__inv_6 _06674_ (.A(net542),
    .Y(_03328_));
 sky130_fd_sc_hd__clkinv_8 _06675_ (.A(net522),
    .Y(_03329_));
 sky130_fd_sc_hd__inv_8 _06676_ (.A(net511),
    .Y(_03330_));
 sky130_fd_sc_hd__inv_2 _06677_ (.A(\core_pipeline.execute_to_memory_rd_address[1] ),
    .Y(_03331_));
 sky130_fd_sc_hd__inv_2 _06678_ (.A(\core_pipeline.execute_to_memory_rd_address[0] ),
    .Y(_03332_));
 sky130_fd_sc_hd__inv_2 _06679_ (.A(\core_pipeline.execute_to_memory_rd_address[3] ),
    .Y(_03333_));
 sky130_fd_sc_hd__inv_2 _06680_ (.A(\core_pipeline.execute_to_memory_rd_address[2] ),
    .Y(_03334_));
 sky130_fd_sc_hd__inv_2 _06681_ (.A(\core_pipeline.execute_to_memory_rd_address[4] ),
    .Y(_03335_));
 sky130_fd_sc_hd__inv_2 _06682_ (.A(\core_pipeline.execute_to_memory_bypass_memory ),
    .Y(_03336_));
 sky130_fd_sc_hd__inv_2 _06683_ (.A(\core_pipeline.decode_to_execute_csr_write ),
    .Y(_03337_));
 sky130_fd_sc_hd__inv_2 _06684_ (.A(net35),
    .Y(_03338_));
 sky130_fd_sc_hd__inv_2 _06685_ (.A(\core_pipeline.decode_to_csr_read_address[10] ),
    .Y(_03339_));
 sky130_fd_sc_hd__inv_2 _06686_ (.A(\core_pipeline.pipeline_csr.mtimecmp[63] ),
    .Y(_03340_));
 sky130_fd_sc_hd__inv_2 _06687_ (.A(\core_pipeline.pipeline_csr.mtimecmp[31] ),
    .Y(_03341_));
 sky130_fd_sc_hd__inv_2 _06688_ (.A(\core_pipeline.pipeline_csr.cycle[31] ),
    .Y(_03342_));
 sky130_fd_sc_hd__inv_2 _06689_ (.A(\core_pipeline.pipeline_csr.mtimecmp[62] ),
    .Y(_03343_));
 sky130_fd_sc_hd__inv_2 _06690_ (.A(\core_pipeline.pipeline_csr.mtimecmp[30] ),
    .Y(_03344_));
 sky130_fd_sc_hd__inv_2 _06691_ (.A(\core_pipeline.pipeline_csr.cycle[30] ),
    .Y(_03345_));
 sky130_fd_sc_hd__inv_2 _06692_ (.A(\core_pipeline.pipeline_csr.mtimecmp[61] ),
    .Y(_03346_));
 sky130_fd_sc_hd__inv_2 _06693_ (.A(\core_pipeline.pipeline_csr.mtimecmp[29] ),
    .Y(_03347_));
 sky130_fd_sc_hd__inv_2 _06694_ (.A(\core_pipeline.pipeline_csr.cycle[29] ),
    .Y(_03348_));
 sky130_fd_sc_hd__inv_2 _06695_ (.A(\core_pipeline.pipeline_csr.cycle[60] ),
    .Y(_03349_));
 sky130_fd_sc_hd__inv_2 _06696_ (.A(\core_pipeline.pipeline_csr.cycle[28] ),
    .Y(_03350_));
 sky130_fd_sc_hd__inv_2 _06697_ (.A(\core_pipeline.pipeline_csr.mtimecmp[59] ),
    .Y(_03351_));
 sky130_fd_sc_hd__inv_2 _06698_ (.A(\core_pipeline.pipeline_csr.cycle[59] ),
    .Y(_03352_));
 sky130_fd_sc_hd__inv_2 _06699_ (.A(\core_pipeline.pipeline_csr.cycle[27] ),
    .Y(_03353_));
 sky130_fd_sc_hd__inv_2 _06700_ (.A(\core_pipeline.pipeline_csr.mtimecmp[58] ),
    .Y(_03354_));
 sky130_fd_sc_hd__inv_2 _06701_ (.A(\core_pipeline.pipeline_csr.cycle[26] ),
    .Y(_03355_));
 sky130_fd_sc_hd__inv_2 _06702_ (.A(\core_pipeline.pipeline_csr.mtimecmp[25] ),
    .Y(_03356_));
 sky130_fd_sc_hd__inv_2 _06703_ (.A(\core_pipeline.pipeline_csr.cycle[57] ),
    .Y(_03357_));
 sky130_fd_sc_hd__inv_2 _06704_ (.A(\core_pipeline.pipeline_csr.mtimecmp[24] ),
    .Y(_03358_));
 sky130_fd_sc_hd__inv_2 _06705_ (.A(\core_pipeline.pipeline_csr.cycle[56] ),
    .Y(_03359_));
 sky130_fd_sc_hd__inv_2 _06706_ (.A(\core_pipeline.pipeline_csr.mtimecmp[23] ),
    .Y(_03360_));
 sky130_fd_sc_hd__inv_2 _06707_ (.A(\core_pipeline.pipeline_csr.cycle[55] ),
    .Y(_03361_));
 sky130_fd_sc_hd__inv_2 _06708_ (.A(\core_pipeline.pipeline_csr.mtimecmp[54] ),
    .Y(_03362_));
 sky130_fd_sc_hd__inv_2 _06709_ (.A(\core_pipeline.pipeline_csr.cycle[22] ),
    .Y(_03363_));
 sky130_fd_sc_hd__inv_2 _06710_ (.A(\core_pipeline.pipeline_csr.mtimecmp[53] ),
    .Y(_03364_));
 sky130_fd_sc_hd__inv_2 _06711_ (.A(\core_pipeline.pipeline_csr.cycle[21] ),
    .Y(_03365_));
 sky130_fd_sc_hd__inv_2 _06712_ (.A(\core_pipeline.pipeline_csr.mtimecmp[20] ),
    .Y(_03366_));
 sky130_fd_sc_hd__inv_2 _06713_ (.A(\core_pipeline.pipeline_csr.cycle[52] ),
    .Y(_03367_));
 sky130_fd_sc_hd__inv_2 _06714_ (.A(\core_pipeline.pipeline_csr.mtimecmp[19] ),
    .Y(_03368_));
 sky130_fd_sc_hd__inv_2 _06715_ (.A(\core_pipeline.pipeline_csr.cycle[51] ),
    .Y(_03369_));
 sky130_fd_sc_hd__inv_2 _06716_ (.A(\core_pipeline.pipeline_csr.mtimecmp[50] ),
    .Y(_03370_));
 sky130_fd_sc_hd__inv_2 _06717_ (.A(\core_pipeline.pipeline_csr.mtimecmp[18] ),
    .Y(_03371_));
 sky130_fd_sc_hd__inv_2 _06718_ (.A(\core_pipeline.pipeline_csr.mtimecmp[49] ),
    .Y(_03372_));
 sky130_fd_sc_hd__inv_2 _06719_ (.A(\core_pipeline.pipeline_csr.mtimecmp[17] ),
    .Y(_03373_));
 sky130_fd_sc_hd__inv_2 _06720_ (.A(\core_pipeline.pipeline_csr.mtimecmp[48] ),
    .Y(_03374_));
 sky130_fd_sc_hd__inv_2 _06721_ (.A(\core_pipeline.pipeline_csr.mtimecmp[16] ),
    .Y(_03375_));
 sky130_fd_sc_hd__inv_2 _06722_ (.A(\core_pipeline.pipeline_csr.cycle[47] ),
    .Y(_03376_));
 sky130_fd_sc_hd__inv_2 _06723_ (.A(\core_pipeline.pipeline_csr.cycle[15] ),
    .Y(_03377_));
 sky130_fd_sc_hd__inv_2 _06724_ (.A(\core_pipeline.pipeline_csr.cycle[46] ),
    .Y(_03378_));
 sky130_fd_sc_hd__inv_2 _06725_ (.A(\core_pipeline.pipeline_csr.cycle[14] ),
    .Y(_03379_));
 sky130_fd_sc_hd__inv_2 _06726_ (.A(\core_pipeline.pipeline_csr.cycle[45] ),
    .Y(_03380_));
 sky130_fd_sc_hd__inv_2 _06727_ (.A(\core_pipeline.pipeline_csr.cycle[13] ),
    .Y(_03381_));
 sky130_fd_sc_hd__clkinv_2 _06728_ (.A(\core_pipeline.pipeline_csr.mtimecmp[44] ),
    .Y(_03382_));
 sky130_fd_sc_hd__inv_2 _06729_ (.A(\core_pipeline.pipeline_csr.cycle[12] ),
    .Y(_03383_));
 sky130_fd_sc_hd__clkinv_2 _06730_ (.A(\core_pipeline.pipeline_csr.mtimecmp[43] ),
    .Y(_03384_));
 sky130_fd_sc_hd__inv_2 _06731_ (.A(\core_pipeline.pipeline_csr.cycle[11] ),
    .Y(_03385_));
 sky130_fd_sc_hd__inv_2 _06732_ (.A(\core_pipeline.pipeline_csr.cycle[42] ),
    .Y(_03386_));
 sky130_fd_sc_hd__inv_2 _06733_ (.A(\core_pipeline.pipeline_csr.cycle[10] ),
    .Y(_03387_));
 sky130_fd_sc_hd__inv_2 _06734_ (.A(\core_pipeline.pipeline_csr.mtimecmp[41] ),
    .Y(_03388_));
 sky130_fd_sc_hd__inv_2 _06735_ (.A(\core_pipeline.pipeline_csr.cycle[9] ),
    .Y(_03389_));
 sky130_fd_sc_hd__inv_2 _06736_ (.A(\core_pipeline.pipeline_csr.mtimecmp[40] ),
    .Y(_03390_));
 sky130_fd_sc_hd__clkinv_2 _06737_ (.A(\core_pipeline.pipeline_csr.cycle[8] ),
    .Y(_03391_));
 sky130_fd_sc_hd__inv_2 _06738_ (.A(\core_pipeline.pipeline_csr.mtimecmp[39] ),
    .Y(_03392_));
 sky130_fd_sc_hd__inv_2 _06739_ (.A(\core_pipeline.pipeline_csr.cycle[7] ),
    .Y(_03393_));
 sky130_fd_sc_hd__inv_2 _06740_ (.A(\core_pipeline.pipeline_csr.mtimecmp[38] ),
    .Y(_03394_));
 sky130_fd_sc_hd__inv_2 _06741_ (.A(\core_pipeline.pipeline_csr.cycle[6] ),
    .Y(_03395_));
 sky130_fd_sc_hd__inv_2 _06742_ (.A(\core_pipeline.pipeline_csr.mtimecmp[37] ),
    .Y(_03396_));
 sky130_fd_sc_hd__inv_2 _06743_ (.A(\core_pipeline.pipeline_csr.cycle[37] ),
    .Y(_03397_));
 sky130_fd_sc_hd__inv_2 _06744_ (.A(\core_pipeline.pipeline_csr.cycle[5] ),
    .Y(_03398_));
 sky130_fd_sc_hd__inv_2 _06745_ (.A(\core_pipeline.pipeline_csr.mtimecmp[36] ),
    .Y(_03399_));
 sky130_fd_sc_hd__inv_2 _06746_ (.A(\core_pipeline.pipeline_csr.cycle[36] ),
    .Y(_03400_));
 sky130_fd_sc_hd__inv_2 _06747_ (.A(\core_pipeline.pipeline_csr.cycle[4] ),
    .Y(_03401_));
 sky130_fd_sc_hd__inv_2 _06748_ (.A(\core_pipeline.pipeline_csr.cycle[35] ),
    .Y(_03402_));
 sky130_fd_sc_hd__inv_2 _06749_ (.A(\core_pipeline.pipeline_csr.cycle[3] ),
    .Y(_03403_));
 sky130_fd_sc_hd__inv_2 _06750_ (.A(\core_pipeline.pipeline_csr.mtimecmp[34] ),
    .Y(_03404_));
 sky130_fd_sc_hd__inv_2 _06751_ (.A(\core_pipeline.pipeline_csr.cycle[34] ),
    .Y(_03405_));
 sky130_fd_sc_hd__inv_2 _06752_ (.A(\core_pipeline.pipeline_csr.cycle[2] ),
    .Y(_03406_));
 sky130_fd_sc_hd__inv_2 _06753_ (.A(\core_pipeline.pipeline_csr.mtimecmp[33] ),
    .Y(_03407_));
 sky130_fd_sc_hd__inv_2 _06754_ (.A(\core_pipeline.pipeline_csr.cycle[33] ),
    .Y(_03408_));
 sky130_fd_sc_hd__inv_2 _06755_ (.A(\core_pipeline.pipeline_csr.cycle[1] ),
    .Y(_03409_));
 sky130_fd_sc_hd__inv_2 _06756_ (.A(\core_pipeline.pipeline_csr.cycle[32] ),
    .Y(_03410_));
 sky130_fd_sc_hd__inv_2 _06757_ (.A(\core_pipeline.pipeline_csr.cycle[0] ),
    .Y(_03411_));
 sky130_fd_sc_hd__inv_2 _06758_ (.A(\core_pipeline.decode_to_execute_csr_read ),
    .Y(_03412_));
 sky130_fd_sc_hd__inv_2 _06759_ (.A(net17),
    .Y(_03413_));
 sky130_fd_sc_hd__inv_2 _06760_ (.A(net18),
    .Y(_03414_));
 sky130_fd_sc_hd__inv_2 _06761_ (.A(net19),
    .Y(_03415_));
 sky130_fd_sc_hd__inv_2 _06762_ (.A(net20),
    .Y(_03416_));
 sky130_fd_sc_hd__inv_2 _06763_ (.A(net21),
    .Y(_03417_));
 sky130_fd_sc_hd__inv_2 _06764_ (.A(net22),
    .Y(_03418_));
 sky130_fd_sc_hd__inv_2 _06765_ (.A(net24),
    .Y(_03419_));
 sky130_fd_sc_hd__inv_2 _06766_ (.A(\core_pipeline.pipeline_execute.ex_alu.old_function[2] ),
    .Y(_03420_));
 sky130_fd_sc_hd__inv_2 _06767_ (.A(\core_pipeline.pipeline_execute.ex_alu.old_function[1] ),
    .Y(_03421_));
 sky130_fd_sc_hd__inv_2 _06768_ (.A(\core_pipeline.decode_to_execute_cmp_function[1] ),
    .Y(_03422_));
 sky130_fd_sc_hd__clkinv_4 _06769_ (.A(net635),
    .Y(_03423_));
 sky130_fd_sc_hd__or2_2 _06770_ (.A(\core_busio.mem_size[1] ),
    .B(\core_busio.mem_size[0] ),
    .X(_03424_));
 sky130_fd_sc_hd__and3b_4 _06771_ (.A_N(net490),
    .B(\core_busio.mem_size[1] ),
    .C(_03316_),
    .X(_03425_));
 sky130_fd_sc_hd__o2bb2a_4 _06772_ (.A1_N(net495),
    .A2_N(_03424_),
    .B1(_03425_),
    .B2(_03315_),
    .X(_03426_));
 sky130_fd_sc_hd__nand2_1 _06773_ (.A(\core_pipeline.execute_to_memory_valid ),
    .B(_03426_),
    .Y(_03427_));
 sky130_fd_sc_hd__nor2_2 _06774_ (.A(\core_pipeline.execute_to_memory_load ),
    .B(\core_pipeline.execute_to_memory_store ),
    .Y(_03428_));
 sky130_fd_sc_hd__nor3_2 _06775_ (.A(\core_pipeline.execute_to_memory_exception ),
    .B(_03427_),
    .C(_03428_),
    .Y(_03429_));
 sky130_fd_sc_hd__inv_4 _06776_ (.A(net261),
    .Y(net66));
 sky130_fd_sc_hd__or2_2 _06777_ (.A(net33),
    .B(net66),
    .X(_03430_));
 sky130_fd_sc_hd__and2_4 _06778_ (.A(net505),
    .B(\core_pipeline.memory_to_writeback_valid ),
    .X(_03431_));
 sky130_fd_sc_hd__nand2_8 _06779_ (.A(net505),
    .B(\core_pipeline.memory_to_writeback_valid ),
    .Y(_03432_));
 sky130_fd_sc_hd__nand2_1 _06780_ (.A(\core_pipeline.execute_to_memory_valid ),
    .B(\core_pipeline.execute_to_memory_mret ),
    .Y(_03433_));
 sky130_fd_sc_hd__and3_4 _06781_ (.A(_03430_),
    .B(net454),
    .C(_03433_),
    .X(_03434_));
 sky130_fd_sc_hd__nand3_2 _06782_ (.A(_03430_),
    .B(net454),
    .C(_03433_),
    .Y(_03435_));
 sky130_fd_sc_hd__and3_1 _06783_ (.A(\core_pipeline.fetch_to_decode_instruction[1] ),
    .B(\core_pipeline.fetch_to_decode_instruction[0] ),
    .C(\core_pipeline.fetch_to_decode_instruction[2] ),
    .X(_03436_));
 sky130_fd_sc_hd__and4b_4 _06784_ (.A_N(\core_pipeline.fetch_to_decode_instruction[4] ),
    .B(_03436_),
    .C(\core_pipeline.fetch_to_decode_instruction[6] ),
    .D(\core_pipeline.fetch_to_decode_instruction[5] ),
    .X(_03437_));
 sky130_fd_sc_hd__nand2b_2 _06785_ (.A_N(\core_pipeline.fetch_to_decode_instruction[3] ),
    .B(_03437_),
    .Y(_03438_));
 sky130_fd_sc_hd__or4bb_2 _06786_ (.A(\core_pipeline.fetch_to_decode_instruction[2] ),
    .B(\core_pipeline.fetch_to_decode_instruction[3] ),
    .C_N(\core_pipeline.fetch_to_decode_instruction[1] ),
    .D_N(\core_pipeline.fetch_to_decode_instruction[0] ),
    .X(_03439_));
 sky130_fd_sc_hd__or2_4 _06787_ (.A(_03322_),
    .B(_03439_),
    .X(_03440_));
 sky130_fd_sc_hd__inv_2 _06788_ (.A(_03440_),
    .Y(_03441_));
 sky130_fd_sc_hd__nor2_8 _06789_ (.A(\core_pipeline.fetch_to_decode_instruction[4] ),
    .B(_03440_),
    .Y(_03442_));
 sky130_fd_sc_hd__nor2_1 _06790_ (.A(\core_pipeline.fetch_to_decode_instruction[6] ),
    .B(_03439_),
    .Y(_03443_));
 sky130_fd_sc_hd__or2_1 _06791_ (.A(\core_pipeline.fetch_to_decode_instruction[6] ),
    .B(_03439_),
    .X(_03444_));
 sky130_fd_sc_hd__and2_2 _06792_ (.A(\core_pipeline.fetch_to_decode_instruction[6] ),
    .B(_03442_),
    .X(_03445_));
 sky130_fd_sc_hd__o211ai_2 _06793_ (.A1(\core_pipeline.fetch_to_decode_instruction[4] ),
    .A2(_03440_),
    .B1(_03444_),
    .C1(_03438_),
    .Y(_03446_));
 sky130_fd_sc_hd__nor2_1 _06794_ (.A(\core_pipeline.fetch_to_decode_instruction[13] ),
    .B(\core_pipeline.fetch_to_decode_instruction[12] ),
    .Y(_03447_));
 sky130_fd_sc_hd__or2_4 _06795_ (.A(\core_pipeline.fetch_to_decode_instruction[13] ),
    .B(\core_pipeline.fetch_to_decode_instruction[12] ),
    .X(_03448_));
 sky130_fd_sc_hd__nor2_1 _06796_ (.A(\core_pipeline.fetch_to_decode_instruction[14] ),
    .B(_03447_),
    .Y(_03449_));
 sky130_fd_sc_hd__inv_2 _06797_ (.A(_03449_),
    .Y(_03450_));
 sky130_fd_sc_hd__and3_4 _06798_ (.A(\core_pipeline.fetch_to_decode_instruction[6] ),
    .B(\core_pipeline.fetch_to_decode_instruction[4] ),
    .C(_03441_),
    .X(_03451_));
 sky130_fd_sc_hd__or2_2 _06799_ (.A(_03446_),
    .B(_03451_),
    .X(_03452_));
 sky130_fd_sc_hd__o211a_2 _06800_ (.A1(_03446_),
    .A2(_03449_),
    .B1(_03452_),
    .C1(\core_pipeline.fetch_to_decode_valid ),
    .X(_03453_));
 sky130_fd_sc_hd__a22o_1 _06801_ (.A1(_03317_),
    .A2(net626),
    .B1(net466),
    .B2(\core_pipeline.decode_to_execute_rd_address[4] ),
    .X(_03454_));
 sky130_fd_sc_hd__o22a_1 _06802_ (.A1(_03317_),
    .A2(net626),
    .B1(net480),
    .B2(\core_pipeline.decode_to_execute_rd_address[2] ),
    .X(_03455_));
 sky130_fd_sc_hd__o221a_1 _06803_ (.A1(\core_pipeline.decode_to_execute_rd_address[1] ),
    .A2(net485),
    .B1(net581),
    .B2(_03319_),
    .C1(_03455_),
    .X(_03456_));
 sky130_fd_sc_hd__a221o_1 _06804_ (.A1(\core_pipeline.decode_to_execute_rd_address[3] ),
    .A2(net471),
    .B1(net569),
    .B2(_03320_),
    .C1(_03454_),
    .X(_03457_));
 sky130_fd_sc_hd__a221oi_1 _06805_ (.A1(\core_pipeline.decode_to_execute_rd_address[1] ),
    .A2(_03323_),
    .B1(net575),
    .B2(_03318_),
    .C1(_03457_),
    .Y(_03458_));
 sky130_fd_sc_hd__and3_1 _06806_ (.A(_03453_),
    .B(_03456_),
    .C(_03458_),
    .X(_03459_));
 sky130_fd_sc_hd__and2_2 _06807_ (.A(\core_pipeline.fetch_to_decode_instruction[4] ),
    .B(_03443_),
    .X(_03460_));
 sky130_fd_sc_hd__and3_2 _06808_ (.A(\core_pipeline.fetch_to_decode_instruction[5] ),
    .B(\core_pipeline.fetch_to_decode_instruction[4] ),
    .C(_03443_),
    .X(_03461_));
 sky130_fd_sc_hd__o21a_1 _06809_ (.A1(_03442_),
    .A2(_03461_),
    .B1(\core_pipeline.fetch_to_decode_valid ),
    .X(_03462_));
 sky130_fd_sc_hd__a22o_1 _06810_ (.A1(\core_pipeline.decode_to_execute_rd_address[0] ),
    .A2(_03327_),
    .B1(net512),
    .B2(_03320_),
    .X(_03463_));
 sky130_fd_sc_hd__a22o_1 _06811_ (.A1(_03317_),
    .A2(net565),
    .B1(net465),
    .B2(\core_pipeline.decode_to_execute_rd_address[2] ),
    .X(_03464_));
 sky130_fd_sc_hd__o22a_1 _06812_ (.A1(\core_pipeline.decode_to_execute_rd_address[1] ),
    .A2(_03328_),
    .B1(net517),
    .B2(_03318_),
    .X(_03465_));
 sky130_fd_sc_hd__a221o_1 _06813_ (.A1(\core_pipeline.decode_to_execute_rd_address[1] ),
    .A2(_03328_),
    .B1(net524),
    .B2(_03319_),
    .C1(_03464_),
    .X(_03466_));
 sky130_fd_sc_hd__a211oi_1 _06814_ (.A1(_03318_),
    .A2(net517),
    .B1(_03463_),
    .C1(_03466_),
    .Y(_03467_));
 sky130_fd_sc_hd__o2111a_1 _06815_ (.A1(_03320_),
    .A2(net512),
    .B1(_03462_),
    .C1(_03465_),
    .D1(_03467_),
    .X(_03468_));
 sky130_fd_sc_hd__or4_1 _06816_ (.A(\core_pipeline.decode_to_execute_rd_address[0] ),
    .B(\core_pipeline.decode_to_execute_rd_address[3] ),
    .C(\core_pipeline.decode_to_execute_rd_address[2] ),
    .D(\core_pipeline.decode_to_execute_rd_address[4] ),
    .X(_03469_));
 sky130_fd_sc_hd__or2_1 _06817_ (.A(\core_pipeline.decode_to_execute_rd_address[1] ),
    .B(_03469_),
    .X(_03470_));
 sky130_fd_sc_hd__o211a_1 _06818_ (.A1(_03459_),
    .A2(_03468_),
    .B1(_03470_),
    .C1(\core_pipeline.decode_to_execute_valid ),
    .X(_03471_));
 sky130_fd_sc_hd__and3_1 _06819_ (.A(\core_pipeline.pipeline_csr.ie ),
    .B(\core_pipeline.pipeline_csr.mtie ),
    .C(\core_pipeline.pipeline_csr.mtip ),
    .X(_03472_));
 sky130_fd_sc_hd__nand3_2 _06820_ (.A(\core_pipeline.pipeline_csr.msie ),
    .B(\core_pipeline.pipeline_csr.ie ),
    .C(\core_pipeline.pipeline_csr.msip ),
    .Y(_03473_));
 sky130_fd_sc_hd__and2b_1 _06821_ (.A_N(_03472_),
    .B(_03473_),
    .X(_03474_));
 sky130_fd_sc_hd__nand3_4 _06822_ (.A(\core_pipeline.pipeline_csr.ie ),
    .B(\core_pipeline.pipeline_csr.meie ),
    .C(net34),
    .Y(_03475_));
 sky130_fd_sc_hd__nand2_1 _06823_ (.A(_03474_),
    .B(_03475_),
    .Y(_03476_));
 sky130_fd_sc_hd__nand2_4 _06824_ (.A(\core_pipeline.memory_to_writeback_valid ),
    .B(\core_pipeline.memory_to_writeback_exception ),
    .Y(_03477_));
 sky130_fd_sc_hd__and4b_4 _06825_ (.A_N(_03472_),
    .B(_03473_),
    .C(_03475_),
    .D(_03477_),
    .X(_03478_));
 sky130_fd_sc_hd__nand2b_4 _06826_ (.A_N(_03476_),
    .B(_03477_),
    .Y(_03479_));
 sky130_fd_sc_hd__and2_4 _06827_ (.A(\core_pipeline.memory_to_writeback_valid ),
    .B(net400),
    .X(_03480_));
 sky130_fd_sc_hd__and3_2 _06828_ (.A(\core_pipeline.memory_to_writeback_valid ),
    .B(\core_pipeline.memory_to_writeback_csr_write ),
    .C(net400),
    .X(_03481_));
 sky130_fd_sc_hd__nand2_4 _06829_ (.A(\core_pipeline.memory_to_writeback_csr_write ),
    .B(_03480_),
    .Y(_03482_));
 sky130_fd_sc_hd__a221o_1 _06830_ (.A1(\core_pipeline.decode_to_execute_valid ),
    .A2(\core_pipeline.decode_to_execute_csr_write ),
    .B1(\core_pipeline.execute_to_memory_csr_write ),
    .B2(\core_pipeline.execute_to_memory_valid ),
    .C1(_03481_),
    .X(_03483_));
 sky130_fd_sc_hd__and2_2 _06831_ (.A(_03448_),
    .B(_03451_),
    .X(_03484_));
 sky130_fd_sc_hd__or3_1 _06832_ (.A(\core_pipeline.fetch_to_decode_instruction[11] ),
    .B(\core_pipeline.fetch_to_decode_instruction[8] ),
    .C(\core_pipeline.fetch_to_decode_instruction[10] ),
    .X(_03485_));
 sky130_fd_sc_hd__or4_1 _06833_ (.A(\core_pipeline.fetch_to_decode_instruction[13] ),
    .B(\core_pipeline.fetch_to_decode_instruction[7] ),
    .C(\core_pipeline.fetch_to_decode_instruction[9] ),
    .D(_03485_),
    .X(_03486_));
 sky130_fd_sc_hd__nand2_1 _06834_ (.A(net517),
    .B(_03333_),
    .Y(_03487_));
 sky130_fd_sc_hd__o221a_1 _06835_ (.A1(_03328_),
    .A2(\core_pipeline.execute_to_memory_rd_address[1] ),
    .B1(\core_pipeline.execute_to_memory_rd_address[4] ),
    .B2(net460),
    .C1(_03487_),
    .X(_03488_));
 sky130_fd_sc_hd__xnor2_1 _06836_ (.A(net524),
    .B(\core_pipeline.execute_to_memory_rd_address[2] ),
    .Y(_03489_));
 sky130_fd_sc_hd__o221a_1 _06837_ (.A1(net565),
    .A2(_03332_),
    .B1(_03333_),
    .B2(net517),
    .C1(_03489_),
    .X(_03490_));
 sky130_fd_sc_hd__o22a_1 _06838_ (.A1(net542),
    .A2(_03331_),
    .B1(_03335_),
    .B2(net513),
    .X(_03491_));
 sky130_fd_sc_hd__o211a_1 _06839_ (.A1(_03327_),
    .A2(\core_pipeline.execute_to_memory_rd_address[0] ),
    .B1(_03490_),
    .C1(_03491_),
    .X(_03492_));
 sky130_fd_sc_hd__o2111a_1 _06840_ (.A1(_03442_),
    .A2(_03461_),
    .B1(_03488_),
    .C1(_03492_),
    .D1(\core_pipeline.fetch_to_decode_valid ),
    .X(_03493_));
 sky130_fd_sc_hd__o22a_1 _06841_ (.A1(net575),
    .A2(_03333_),
    .B1(_03335_),
    .B2(net569),
    .X(_03494_));
 sky130_fd_sc_hd__o221a_1 _06842_ (.A1(net602),
    .A2(_03331_),
    .B1(\core_pipeline.execute_to_memory_rd_address[2] ),
    .B2(net480),
    .C1(_03494_),
    .X(_03495_));
 sky130_fd_sc_hd__xnor2_1 _06843_ (.A(net626),
    .B(\core_pipeline.execute_to_memory_rd_address[0] ),
    .Y(_03496_));
 sky130_fd_sc_hd__o211a_1 _06844_ (.A1(net581),
    .A2(_03334_),
    .B1(_03495_),
    .C1(_03496_),
    .X(_03497_));
 sky130_fd_sc_hd__nand2_1 _06845_ (.A(net602),
    .B(_03331_),
    .Y(_03498_));
 sky130_fd_sc_hd__o221a_1 _06846_ (.A1(net471),
    .A2(\core_pipeline.execute_to_memory_rd_address[3] ),
    .B1(\core_pipeline.execute_to_memory_rd_address[4] ),
    .B2(_03326_),
    .C1(_03498_),
    .X(_03499_));
 sky130_fd_sc_hd__a31o_1 _06847_ (.A1(_03453_),
    .A2(_03497_),
    .A3(_03499_),
    .B1(_03493_),
    .X(_03500_));
 sky130_fd_sc_hd__or4_1 _06848_ (.A(\core_pipeline.execute_to_memory_rd_address[0] ),
    .B(\core_pipeline.execute_to_memory_rd_address[3] ),
    .C(\core_pipeline.execute_to_memory_rd_address[2] ),
    .D(\core_pipeline.execute_to_memory_rd_address[4] ),
    .X(_03501_));
 sky130_fd_sc_hd__o2111a_1 _06849_ (.A1(\core_pipeline.execute_to_memory_rd_address[1] ),
    .A2(_03501_),
    .B1(_03336_),
    .C1(\core_pipeline.execute_to_memory_valid ),
    .D1(_03500_),
    .X(_03502_));
 sky130_fd_sc_hd__a41o_1 _06850_ (.A1(\core_pipeline.fetch_to_decode_valid ),
    .A2(_03483_),
    .A3(_03484_),
    .A4(_03486_),
    .B1(_03502_),
    .X(_03503_));
 sky130_fd_sc_hd__nor2_1 _06851_ (.A(_03471_),
    .B(_03503_),
    .Y(_03504_));
 sky130_fd_sc_hd__nand2_2 _06852_ (.A(net147),
    .B(_03504_),
    .Y(_03505_));
 sky130_fd_sc_hd__inv_8 _06853_ (.A(net111),
    .Y(_03506_));
 sky130_fd_sc_hd__xor2_1 _06854_ (.A(\core_pipeline.pipeline_execute.ex_cmp.negate ),
    .B(\core_pipeline.pipeline_execute.ex_cmp.quasi_result ),
    .X(_03507_));
 sky130_fd_sc_hd__o21ai_2 _06855_ (.A1(\core_pipeline.execute_to_memory_jump ),
    .A2(_03507_),
    .B1(\core_pipeline.execute_to_memory_branch ),
    .Y(_03508_));
 sky130_fd_sc_hd__nor2_8 _06856_ (.A(net492),
    .B(net494),
    .Y(_03509_));
 sky130_fd_sc_hd__or4b_4 _06857_ (.A(net492),
    .B(net494),
    .C(_03508_),
    .D_N(\core_pipeline.execute_to_memory_valid ),
    .X(_03510_));
 sky130_fd_sc_hd__inv_4 _06858_ (.A(net351),
    .Y(_03511_));
 sky130_fd_sc_hd__and2_4 _06859_ (.A(\core_pipeline.memory_to_writeback_valid ),
    .B(\core_pipeline.memory_to_writeback_mret ),
    .X(_03512_));
 sky130_fd_sc_hd__nand2_8 _06860_ (.A(\core_pipeline.memory_to_writeback_valid ),
    .B(\core_pipeline.memory_to_writeback_mret ),
    .Y(_03513_));
 sky130_fd_sc_hd__nor2_8 _06861_ (.A(_03479_),
    .B(_03512_),
    .Y(_03514_));
 sky130_fd_sc_hd__nand2_2 _06862_ (.A(net400),
    .B(net445),
    .Y(_03515_));
 sky130_fd_sc_hd__or2_4 _06863_ (.A(_03511_),
    .B(_03515_),
    .X(_03516_));
 sky130_fd_sc_hd__nor2_4 _06864_ (.A(net35),
    .B(_03516_),
    .Y(_03517_));
 sky130_fd_sc_hd__and4_2 _06865_ (.A(net33),
    .B(net66),
    .C(_03506_),
    .D(_03517_),
    .X(_00004_));
 sky130_fd_sc_hd__a2bb2o_1 _06866_ (.A1_N(_03349_),
    .A2_N(\core_pipeline.pipeline_csr.mtimecmp[60] ),
    .B1(\core_pipeline.pipeline_csr.cycle[61] ),
    .B2(_03346_),
    .X(_03518_));
 sky130_fd_sc_hd__a22o_1 _06867_ (.A1(_03351_),
    .A2(\core_pipeline.pipeline_csr.cycle[59] ),
    .B1(_03354_),
    .B2(\core_pipeline.pipeline_csr.cycle[58] ),
    .X(_03519_));
 sky130_fd_sc_hd__a22o_1 _06868_ (.A1(_03340_),
    .A2(\core_pipeline.pipeline_csr.cycle[63] ),
    .B1(_03343_),
    .B2(\core_pipeline.pipeline_csr.cycle[62] ),
    .X(_03520_));
 sky130_fd_sc_hd__o22a_1 _06869_ (.A1(\core_pipeline.pipeline_csr.mtimecmp[57] ),
    .A2(_03357_),
    .B1(\core_pipeline.pipeline_csr.mtimecmp[56] ),
    .B2(_03359_),
    .X(_03521_));
 sky130_fd_sc_hd__a2bb2o_1 _06870_ (.A1_N(_03354_),
    .A2_N(\core_pipeline.pipeline_csr.cycle[58] ),
    .B1(\core_pipeline.pipeline_csr.mtimecmp[57] ),
    .B2(_03357_),
    .X(_03522_));
 sky130_fd_sc_hd__nor2_1 _06871_ (.A(_03521_),
    .B(_03522_),
    .Y(_03523_));
 sky130_fd_sc_hd__or2_1 _06872_ (.A(_03340_),
    .B(\core_pipeline.pipeline_csr.cycle[63] ),
    .X(_03524_));
 sky130_fd_sc_hd__nand2_1 _06873_ (.A(\core_pipeline.pipeline_csr.mtimecmp[60] ),
    .B(_03349_),
    .Y(_03525_));
 sky130_fd_sc_hd__or2_1 _06874_ (.A(_03343_),
    .B(\core_pipeline.pipeline_csr.cycle[62] ),
    .X(_03526_));
 sky130_fd_sc_hd__o221a_1 _06875_ (.A1(_03351_),
    .A2(\core_pipeline.pipeline_csr.cycle[59] ),
    .B1(_03519_),
    .B2(_03523_),
    .C1(_03525_),
    .X(_03527_));
 sky130_fd_sc_hd__o221a_1 _06876_ (.A1(_03346_),
    .A2(\core_pipeline.pipeline_csr.cycle[61] ),
    .B1(_03518_),
    .B2(_03527_),
    .C1(_03526_),
    .X(_03528_));
 sky130_fd_sc_hd__or2_1 _06877_ (.A(_03520_),
    .B(_03528_),
    .X(_03529_));
 sky130_fd_sc_hd__a2bb2o_1 _06878_ (.A1_N(_03346_),
    .A2_N(\core_pipeline.pipeline_csr.cycle[61] ),
    .B1(\core_pipeline.pipeline_csr.mtimecmp[55] ),
    .B2(_03361_),
    .X(_03530_));
 sky130_fd_sc_hd__nand3_1 _06879_ (.A(_03521_),
    .B(_03524_),
    .C(_03526_),
    .Y(_03531_));
 sky130_fd_sc_hd__a221o_1 _06880_ (.A1(\core_pipeline.pipeline_csr.mtimecmp[60] ),
    .A2(_03349_),
    .B1(\core_pipeline.pipeline_csr.mtimecmp[59] ),
    .B2(_03352_),
    .C1(_03522_),
    .X(_03532_));
 sky130_fd_sc_hd__a2111o_1 _06881_ (.A1(\core_pipeline.pipeline_csr.mtimecmp[56] ),
    .A2(_03359_),
    .B1(_03530_),
    .C1(_03531_),
    .D1(_03532_),
    .X(_03533_));
 sky130_fd_sc_hd__nor4_1 _06882_ (.A(_03518_),
    .B(_03519_),
    .C(_03520_),
    .D(_03533_),
    .Y(_03534_));
 sky130_fd_sc_hd__o22a_1 _06883_ (.A1(\core_pipeline.pipeline_csr.mtimecmp[31] ),
    .A2(_03342_),
    .B1(\core_pipeline.pipeline_csr.mtimecmp[30] ),
    .B2(_03345_),
    .X(_03535_));
 sky130_fd_sc_hd__o22a_1 _06884_ (.A1(\core_pipeline.pipeline_csr.mtimecmp[29] ),
    .A2(_03348_),
    .B1(\core_pipeline.pipeline_csr.mtimecmp[28] ),
    .B2(_03350_),
    .X(_03536_));
 sky130_fd_sc_hd__a22o_1 _06885_ (.A1(\core_pipeline.pipeline_csr.mtimecmp[28] ),
    .A2(_03350_),
    .B1(\core_pipeline.pipeline_csr.mtimecmp[27] ),
    .B2(_03353_),
    .X(_03537_));
 sky130_fd_sc_hd__o2bb2a_1 _06886_ (.A1_N(\core_pipeline.pipeline_csr.mtimecmp[26] ),
    .A2_N(_03355_),
    .B1(_03356_),
    .B2(\core_pipeline.pipeline_csr.cycle[25] ),
    .X(_03538_));
 sky130_fd_sc_hd__a22o_1 _06887_ (.A1(_03356_),
    .A2(\core_pipeline.pipeline_csr.cycle[25] ),
    .B1(_03358_),
    .B2(\core_pipeline.pipeline_csr.cycle[24] ),
    .X(_03539_));
 sky130_fd_sc_hd__nand2_1 _06888_ (.A(_03538_),
    .B(_03539_),
    .Y(_03540_));
 sky130_fd_sc_hd__o221a_1 _06889_ (.A1(\core_pipeline.pipeline_csr.mtimecmp[27] ),
    .A2(_03353_),
    .B1(\core_pipeline.pipeline_csr.mtimecmp[26] ),
    .B2(_03355_),
    .C1(_03540_),
    .X(_03541_));
 sky130_fd_sc_hd__o21a_1 _06890_ (.A1(_03537_),
    .A2(_03541_),
    .B1(_03536_),
    .X(_03542_));
 sky130_fd_sc_hd__a221o_1 _06891_ (.A1(\core_pipeline.pipeline_csr.mtimecmp[30] ),
    .A2(_03345_),
    .B1(\core_pipeline.pipeline_csr.mtimecmp[29] ),
    .B2(_03348_),
    .C1(_03542_),
    .X(_03543_));
 sky130_fd_sc_hd__a22o_1 _06892_ (.A1(\core_pipeline.pipeline_csr.mtimecmp[31] ),
    .A2(_03342_),
    .B1(_03535_),
    .B2(_03543_),
    .X(_03544_));
 sky130_fd_sc_hd__o22a_1 _06893_ (.A1(\core_pipeline.pipeline_csr.mtimecmp[15] ),
    .A2(_03377_),
    .B1(\core_pipeline.pipeline_csr.mtimecmp[14] ),
    .B2(_03379_),
    .X(_03545_));
 sky130_fd_sc_hd__and2_1 _06894_ (.A(\core_pipeline.pipeline_csr.mtimecmp[15] ),
    .B(_03377_),
    .X(_03546_));
 sky130_fd_sc_hd__o211a_1 _06895_ (.A1(\core_pipeline.pipeline_csr.mtimecmp[1] ),
    .A2(_03409_),
    .B1(\core_pipeline.pipeline_csr.mtimecmp[0] ),
    .C1(_03411_),
    .X(_03547_));
 sky130_fd_sc_hd__a221o_1 _06896_ (.A1(\core_pipeline.pipeline_csr.mtimecmp[2] ),
    .A2(_03406_),
    .B1(\core_pipeline.pipeline_csr.mtimecmp[1] ),
    .B2(_03409_),
    .C1(_03547_),
    .X(_03548_));
 sky130_fd_sc_hd__o221a_1 _06897_ (.A1(\core_pipeline.pipeline_csr.mtimecmp[3] ),
    .A2(_03403_),
    .B1(\core_pipeline.pipeline_csr.mtimecmp[2] ),
    .B2(_03406_),
    .C1(_03548_),
    .X(_03549_));
 sky130_fd_sc_hd__a221o_1 _06898_ (.A1(\core_pipeline.pipeline_csr.mtimecmp[4] ),
    .A2(_03401_),
    .B1(\core_pipeline.pipeline_csr.mtimecmp[3] ),
    .B2(_03403_),
    .C1(_03549_),
    .X(_03550_));
 sky130_fd_sc_hd__o221a_1 _06899_ (.A1(\core_pipeline.pipeline_csr.mtimecmp[5] ),
    .A2(_03398_),
    .B1(\core_pipeline.pipeline_csr.mtimecmp[4] ),
    .B2(_03401_),
    .C1(_03550_),
    .X(_03551_));
 sky130_fd_sc_hd__a221o_1 _06900_ (.A1(\core_pipeline.pipeline_csr.mtimecmp[6] ),
    .A2(_03395_),
    .B1(\core_pipeline.pipeline_csr.mtimecmp[5] ),
    .B2(_03398_),
    .C1(_03551_),
    .X(_03552_));
 sky130_fd_sc_hd__o221a_1 _06901_ (.A1(\core_pipeline.pipeline_csr.mtimecmp[7] ),
    .A2(_03393_),
    .B1(\core_pipeline.pipeline_csr.mtimecmp[6] ),
    .B2(_03395_),
    .C1(_03552_),
    .X(_03553_));
 sky130_fd_sc_hd__a221o_1 _06902_ (.A1(\core_pipeline.pipeline_csr.mtimecmp[8] ),
    .A2(_03391_),
    .B1(\core_pipeline.pipeline_csr.mtimecmp[7] ),
    .B2(_03393_),
    .C1(_03553_),
    .X(_03554_));
 sky130_fd_sc_hd__o221a_1 _06903_ (.A1(\core_pipeline.pipeline_csr.mtimecmp[9] ),
    .A2(_03389_),
    .B1(\core_pipeline.pipeline_csr.mtimecmp[8] ),
    .B2(_03391_),
    .C1(_03554_),
    .X(_03555_));
 sky130_fd_sc_hd__a221o_1 _06904_ (.A1(\core_pipeline.pipeline_csr.mtimecmp[10] ),
    .A2(_03387_),
    .B1(\core_pipeline.pipeline_csr.mtimecmp[9] ),
    .B2(_03389_),
    .C1(_03555_),
    .X(_03556_));
 sky130_fd_sc_hd__o221a_1 _06905_ (.A1(\core_pipeline.pipeline_csr.mtimecmp[11] ),
    .A2(_03385_),
    .B1(\core_pipeline.pipeline_csr.mtimecmp[10] ),
    .B2(_03387_),
    .C1(_03556_),
    .X(_03557_));
 sky130_fd_sc_hd__a221o_1 _06906_ (.A1(\core_pipeline.pipeline_csr.mtimecmp[12] ),
    .A2(_03383_),
    .B1(\core_pipeline.pipeline_csr.mtimecmp[11] ),
    .B2(_03385_),
    .C1(_03557_),
    .X(_03558_));
 sky130_fd_sc_hd__o22a_1 _06907_ (.A1(\core_pipeline.pipeline_csr.mtimecmp[13] ),
    .A2(_03381_),
    .B1(\core_pipeline.pipeline_csr.mtimecmp[12] ),
    .B2(_03383_),
    .X(_03559_));
 sky130_fd_sc_hd__a221o_1 _06908_ (.A1(\core_pipeline.pipeline_csr.mtimecmp[14] ),
    .A2(_03379_),
    .B1(\core_pipeline.pipeline_csr.mtimecmp[13] ),
    .B2(_03381_),
    .C1(_03546_),
    .X(_03560_));
 sky130_fd_sc_hd__a21o_1 _06909_ (.A1(_03558_),
    .A2(_03559_),
    .B1(_03560_),
    .X(_03561_));
 sky130_fd_sc_hd__mux2_1 _06910_ (.A0(_03546_),
    .A1(_03561_),
    .S(_03545_),
    .X(_03562_));
 sky130_fd_sc_hd__o22a_1 _06911_ (.A1(_03371_),
    .A2(\core_pipeline.pipeline_csr.cycle[18] ),
    .B1(_03373_),
    .B2(\core_pipeline.pipeline_csr.cycle[17] ),
    .X(_03563_));
 sky130_fd_sc_hd__a22o_1 _06912_ (.A1(_03373_),
    .A2(\core_pipeline.pipeline_csr.cycle[17] ),
    .B1(_03375_),
    .B2(\core_pipeline.pipeline_csr.cycle[16] ),
    .X(_03564_));
 sky130_fd_sc_hd__a2bb2o_1 _06913_ (.A1_N(_03363_),
    .A2_N(\core_pipeline.pipeline_csr.mtimecmp[22] ),
    .B1(\core_pipeline.pipeline_csr.cycle[23] ),
    .B2(_03360_),
    .X(_03565_));
 sky130_fd_sc_hd__a22o_1 _06914_ (.A1(\core_pipeline.pipeline_csr.mtimecmp[22] ),
    .A2(_03363_),
    .B1(\core_pipeline.pipeline_csr.mtimecmp[21] ),
    .B2(_03365_),
    .X(_03566_));
 sky130_fd_sc_hd__a22o_1 _06915_ (.A1(_03368_),
    .A2(\core_pipeline.pipeline_csr.cycle[19] ),
    .B1(_03371_),
    .B2(\core_pipeline.pipeline_csr.cycle[18] ),
    .X(_03567_));
 sky130_fd_sc_hd__o22a_1 _06916_ (.A1(_03366_),
    .A2(\core_pipeline.pipeline_csr.cycle[20] ),
    .B1(_03368_),
    .B2(\core_pipeline.pipeline_csr.cycle[19] ),
    .X(_03568_));
 sky130_fd_sc_hd__a2bb2o_1 _06917_ (.A1_N(\core_pipeline.pipeline_csr.mtimecmp[21] ),
    .A2_N(_03365_),
    .B1(_03366_),
    .B2(\core_pipeline.pipeline_csr.cycle[20] ),
    .X(_03569_));
 sky130_fd_sc_hd__or2_1 _06918_ (.A(_03360_),
    .B(\core_pipeline.pipeline_csr.cycle[23] ),
    .X(_03570_));
 sky130_fd_sc_hd__nor2_1 _06919_ (.A(_03375_),
    .B(\core_pipeline.pipeline_csr.cycle[16] ),
    .Y(_03571_));
 sky130_fd_sc_hd__or3b_2 _06920_ (.A(_03565_),
    .B(_03566_),
    .C_N(_03570_),
    .X(_03572_));
 sky130_fd_sc_hd__or4bb_1 _06921_ (.A(_03571_),
    .B(_03569_),
    .C_N(_03568_),
    .D_N(_03563_),
    .X(_03573_));
 sky130_fd_sc_hd__or3_1 _06922_ (.A(_03567_),
    .B(_03572_),
    .C(_03573_),
    .X(_03574_));
 sky130_fd_sc_hd__or3_2 _06923_ (.A(_03562_),
    .B(_03564_),
    .C(_03574_),
    .X(_03575_));
 sky130_fd_sc_hd__a21o_1 _06924_ (.A1(_03563_),
    .A2(_03564_),
    .B1(_03567_),
    .X(_03576_));
 sky130_fd_sc_hd__a21oi_1 _06925_ (.A1(_03568_),
    .A2(_03576_),
    .B1(_03569_),
    .Y(_03577_));
 sky130_fd_sc_hd__o2bb2a_1 _06926_ (.A1_N(_03565_),
    .A2_N(_03570_),
    .B1(_03572_),
    .B2(_03577_),
    .X(_03578_));
 sky130_fd_sc_hd__o221a_1 _06927_ (.A1(\core_pipeline.pipeline_csr.mtimecmp[27] ),
    .A2(_03353_),
    .B1(\core_pipeline.pipeline_csr.mtimecmp[26] ),
    .B2(_03355_),
    .C1(_03538_),
    .X(_03579_));
 sky130_fd_sc_hd__o221a_1 _06928_ (.A1(_03341_),
    .A2(\core_pipeline.pipeline_csr.cycle[31] ),
    .B1(_03358_),
    .B2(\core_pipeline.pipeline_csr.cycle[24] ),
    .C1(_03535_),
    .X(_03580_));
 sky130_fd_sc_hd__or3b_1 _06929_ (.A(_03537_),
    .B(_03539_),
    .C_N(_03579_),
    .X(_03581_));
 sky130_fd_sc_hd__o221a_1 _06930_ (.A1(_03344_),
    .A2(\core_pipeline.pipeline_csr.cycle[30] ),
    .B1(_03347_),
    .B2(\core_pipeline.pipeline_csr.cycle[29] ),
    .C1(_03536_),
    .X(_03582_));
 sky130_fd_sc_hd__nand2_1 _06931_ (.A(_03580_),
    .B(_03582_),
    .Y(_03583_));
 sky130_fd_sc_hd__a211o_1 _06932_ (.A1(_03575_),
    .A2(_03578_),
    .B1(_03581_),
    .C1(_03583_),
    .X(_03584_));
 sky130_fd_sc_hd__a22o_2 _06933_ (.A1(_03388_),
    .A2(\core_pipeline.pipeline_csr.cycle[41] ),
    .B1(_03390_),
    .B2(\core_pipeline.pipeline_csr.cycle[40] ),
    .X(_03585_));
 sky130_fd_sc_hd__o2bb2a_1 _06934_ (.A1_N(_03384_),
    .A2_N(\core_pipeline.pipeline_csr.cycle[43] ),
    .B1(\core_pipeline.pipeline_csr.mtimecmp[42] ),
    .B2(_03386_),
    .X(_03586_));
 sky130_fd_sc_hd__o22a_1 _06935_ (.A1(\core_pipeline.pipeline_csr.mtimecmp[47] ),
    .A2(_03376_),
    .B1(\core_pipeline.pipeline_csr.mtimecmp[46] ),
    .B2(_03378_),
    .X(_03587_));
 sky130_fd_sc_hd__nand2_1 _06936_ (.A(\core_pipeline.pipeline_csr.mtimecmp[47] ),
    .B(_03376_),
    .Y(_03588_));
 sky130_fd_sc_hd__o221a_1 _06937_ (.A1(_03390_),
    .A2(\core_pipeline.pipeline_csr.cycle[40] ),
    .B1(_03392_),
    .B2(\core_pipeline.pipeline_csr.cycle[39] ),
    .C1(_03588_),
    .X(_03589_));
 sky130_fd_sc_hd__o2bb2a_1 _06938_ (.A1_N(\core_pipeline.pipeline_csr.mtimecmp[42] ),
    .A2_N(_03386_),
    .B1(_03388_),
    .B2(\core_pipeline.pipeline_csr.cycle[41] ),
    .X(_03590_));
 sky130_fd_sc_hd__o2bb2a_1 _06939_ (.A1_N(\core_pipeline.pipeline_csr.cycle[44] ),
    .A2_N(_03382_),
    .B1(_03380_),
    .B2(\core_pipeline.pipeline_csr.mtimecmp[45] ),
    .X(_03591_));
 sky130_fd_sc_hd__a22o_2 _06940_ (.A1(\core_pipeline.pipeline_csr.mtimecmp[46] ),
    .A2(_03378_),
    .B1(\core_pipeline.pipeline_csr.mtimecmp[45] ),
    .B2(_03380_),
    .X(_03592_));
 sky130_fd_sc_hd__nand3_2 _06941_ (.A(_03587_),
    .B(_03590_),
    .C(_03591_),
    .Y(_03593_));
 sky130_fd_sc_hd__o221a_1 _06942_ (.A1(_03382_),
    .A2(\core_pipeline.pipeline_csr.cycle[44] ),
    .B1(_03384_),
    .B2(\core_pipeline.pipeline_csr.cycle[43] ),
    .C1(_03586_),
    .X(_03594_));
 sky130_fd_sc_hd__nand2_1 _06943_ (.A(_03589_),
    .B(_03594_),
    .Y(_03595_));
 sky130_fd_sc_hd__nor4_4 _06944_ (.A(_03585_),
    .B(_03592_),
    .C(_03593_),
    .D(_03595_),
    .Y(_03596_));
 sky130_fd_sc_hd__inv_2 _06945_ (.A(_03596_),
    .Y(_03597_));
 sky130_fd_sc_hd__a22o_2 _06946_ (.A1(_03392_),
    .A2(\core_pipeline.pipeline_csr.cycle[39] ),
    .B1(_03394_),
    .B2(\core_pipeline.pipeline_csr.cycle[38] ),
    .X(_03598_));
 sky130_fd_sc_hd__a221o_1 _06947_ (.A1(_03396_),
    .A2(\core_pipeline.pipeline_csr.cycle[37] ),
    .B1(_03399_),
    .B2(\core_pipeline.pipeline_csr.cycle[36] ),
    .C1(_03598_),
    .X(_03599_));
 sky130_fd_sc_hd__a2bb2o_1 _06948_ (.A1_N(_03410_),
    .A2_N(\core_pipeline.pipeline_csr.mtimecmp[32] ),
    .B1(\core_pipeline.pipeline_csr.cycle[33] ),
    .B2(_03407_),
    .X(_03600_));
 sky130_fd_sc_hd__a2bb2o_1 _06949_ (.A1_N(_03394_),
    .A2_N(\core_pipeline.pipeline_csr.cycle[38] ),
    .B1(\core_pipeline.pipeline_csr.mtimecmp[37] ),
    .B2(_03397_),
    .X(_03601_));
 sky130_fd_sc_hd__a2bb2o_1 _06950_ (.A1_N(\core_pipeline.pipeline_csr.mtimecmp[35] ),
    .A2_N(_03402_),
    .B1(_03404_),
    .B2(\core_pipeline.pipeline_csr.cycle[34] ),
    .X(_03602_));
 sky130_fd_sc_hd__a221o_1 _06951_ (.A1(\core_pipeline.pipeline_csr.mtimecmp[34] ),
    .A2(_03405_),
    .B1(\core_pipeline.pipeline_csr.mtimecmp[33] ),
    .B2(_03408_),
    .C1(_03602_),
    .X(_03603_));
 sky130_fd_sc_hd__a221o_1 _06952_ (.A1(\core_pipeline.pipeline_csr.mtimecmp[36] ),
    .A2(_03400_),
    .B1(\core_pipeline.pipeline_csr.mtimecmp[35] ),
    .B2(_03402_),
    .C1(_03600_),
    .X(_03604_));
 sky130_fd_sc_hd__a2111o_1 _06953_ (.A1(\core_pipeline.pipeline_csr.mtimecmp[32] ),
    .A2(_03410_),
    .B1(_03599_),
    .C1(_03601_),
    .D1(_03604_),
    .X(_03605_));
 sky130_fd_sc_hd__a2111o_2 _06954_ (.A1(_03544_),
    .A2(_03584_),
    .B1(_03597_),
    .C1(_03603_),
    .D1(_03605_),
    .X(_03606_));
 sky130_fd_sc_hd__a21bo_1 _06955_ (.A1(_03585_),
    .A2(_03590_),
    .B1_N(_03586_),
    .X(_03607_));
 sky130_fd_sc_hd__o221ai_4 _06956_ (.A1(_03382_),
    .A2(\core_pipeline.pipeline_csr.cycle[44] ),
    .B1(_03384_),
    .B2(\core_pipeline.pipeline_csr.cycle[43] ),
    .C1(_03607_),
    .Y(_03608_));
 sky130_fd_sc_hd__a21o_1 _06957_ (.A1(_03591_),
    .A2(_03608_),
    .B1(_03592_),
    .X(_03609_));
 sky130_fd_sc_hd__a21bo_1 _06958_ (.A1(_03587_),
    .A2(_03609_),
    .B1_N(_03588_),
    .X(_03610_));
 sky130_fd_sc_hd__o221a_1 _06959_ (.A1(_03404_),
    .A2(\core_pipeline.pipeline_csr.cycle[34] ),
    .B1(_03407_),
    .B2(\core_pipeline.pipeline_csr.cycle[33] ),
    .C1(_03600_),
    .X(_03611_));
 sky130_fd_sc_hd__nor2_1 _06960_ (.A(_03602_),
    .B(_03611_),
    .Y(_03612_));
 sky130_fd_sc_hd__a221o_1 _06961_ (.A1(\core_pipeline.pipeline_csr.mtimecmp[36] ),
    .A2(_03400_),
    .B1(\core_pipeline.pipeline_csr.mtimecmp[35] ),
    .B2(_03402_),
    .C1(_03612_),
    .X(_03613_));
 sky130_fd_sc_hd__o221a_1 _06962_ (.A1(\core_pipeline.pipeline_csr.mtimecmp[37] ),
    .A2(_03397_),
    .B1(\core_pipeline.pipeline_csr.mtimecmp[36] ),
    .B2(_03400_),
    .C1(_03613_),
    .X(_03614_));
 sky130_fd_sc_hd__nor2_1 _06963_ (.A(_03601_),
    .B(_03614_),
    .Y(_03615_));
 sky130_fd_sc_hd__o21ai_2 _06964_ (.A1(_03598_),
    .A2(_03615_),
    .B1(_03596_),
    .Y(_03616_));
 sky130_fd_sc_hd__a22o_1 _06965_ (.A1(\core_pipeline.pipeline_csr.mtimecmp[52] ),
    .A2(_03367_),
    .B1(\core_pipeline.pipeline_csr.mtimecmp[51] ),
    .B2(_03369_),
    .X(_03617_));
 sky130_fd_sc_hd__a2bb2o_1 _06966_ (.A1_N(\core_pipeline.pipeline_csr.mtimecmp[51] ),
    .A2_N(_03369_),
    .B1(_03370_),
    .B2(\core_pipeline.pipeline_csr.cycle[50] ),
    .X(_03618_));
 sky130_fd_sc_hd__a22o_1 _06967_ (.A1(_03372_),
    .A2(\core_pipeline.pipeline_csr.cycle[49] ),
    .B1(_03374_),
    .B2(\core_pipeline.pipeline_csr.cycle[48] ),
    .X(_03619_));
 sky130_fd_sc_hd__o22ai_2 _06968_ (.A1(_03370_),
    .A2(\core_pipeline.pipeline_csr.cycle[50] ),
    .B1(_03372_),
    .B2(\core_pipeline.pipeline_csr.cycle[49] ),
    .Y(_03620_));
 sky130_fd_sc_hd__or4_1 _06969_ (.A(_03617_),
    .B(_03618_),
    .C(_03619_),
    .D(_03620_),
    .X(_03621_));
 sky130_fd_sc_hd__a2bb2o_1 _06970_ (.A1_N(\core_pipeline.pipeline_csr.mtimecmp[55] ),
    .A2_N(_03361_),
    .B1(_03362_),
    .B2(\core_pipeline.pipeline_csr.cycle[54] ),
    .X(_03622_));
 sky130_fd_sc_hd__o22a_1 _06971_ (.A1(_03362_),
    .A2(\core_pipeline.pipeline_csr.cycle[54] ),
    .B1(_03364_),
    .B2(\core_pipeline.pipeline_csr.cycle[53] ),
    .X(_03623_));
 sky130_fd_sc_hd__o2bb2a_1 _06972_ (.A1_N(_03364_),
    .A2_N(\core_pipeline.pipeline_csr.cycle[53] ),
    .B1(\core_pipeline.pipeline_csr.mtimecmp[52] ),
    .B2(_03367_),
    .X(_03624_));
 sky130_fd_sc_hd__o211a_1 _06973_ (.A1(_03374_),
    .A2(\core_pipeline.pipeline_csr.cycle[48] ),
    .B1(_03623_),
    .C1(_03624_),
    .X(_03625_));
 sky130_fd_sc_hd__or3b_2 _06974_ (.A(_03621_),
    .B(_03622_),
    .C_N(_03625_),
    .X(_03626_));
 sky130_fd_sc_hd__a31oi_2 _06975_ (.A1(_03606_),
    .A2(_03610_),
    .A3(_03616_),
    .B1(_03626_),
    .Y(_03627_));
 sky130_fd_sc_hd__and2b_1 _06976_ (.A_N(_03620_),
    .B(_03619_),
    .X(_03628_));
 sky130_fd_sc_hd__nor2_1 _06977_ (.A(_03618_),
    .B(_03628_),
    .Y(_03629_));
 sky130_fd_sc_hd__o21ai_1 _06978_ (.A1(_03617_),
    .A2(_03629_),
    .B1(_03624_),
    .Y(_03630_));
 sky130_fd_sc_hd__a211o_1 _06979_ (.A1(_03623_),
    .A2(_03630_),
    .B1(_03627_),
    .C1(_03622_),
    .X(_03631_));
 sky130_fd_sc_hd__a22o_2 _06980_ (.A1(_03524_),
    .A2(_03529_),
    .B1(_03534_),
    .B2(_03631_),
    .X(_00003_));
 sky130_fd_sc_hd__and2_4 _06981_ (.A(net142),
    .B(_03451_),
    .X(_03632_));
 sky130_fd_sc_hd__a22o_1 _06982_ (.A1(net501),
    .A2(net126),
    .B1(_03632_),
    .B2(\core_pipeline.fetch_to_decode_instruction[13] ),
    .X(_00002_));
 sky130_fd_sc_hd__a211o_1 _06983_ (.A1(\core_pipeline.fetch_to_decode_instruction[13] ),
    .A2(_03451_),
    .B1(_03461_),
    .C1(net126),
    .X(_03633_));
 sky130_fd_sc_hd__a21bo_1 _06984_ (.A1(net503),
    .A2(net126),
    .B1_N(_03633_),
    .X(_00001_));
 sky130_fd_sc_hd__nand2_1 _06985_ (.A(\core_pipeline.fetch_to_decode_instruction[3] ),
    .B(_03436_),
    .Y(_03634_));
 sky130_fd_sc_hd__and2_1 _06986_ (.A(\core_pipeline.fetch_to_decode_instruction[3] ),
    .B(_03437_),
    .X(_03635_));
 sky130_fd_sc_hd__and4bb_4 _06987_ (.A_N(\core_pipeline.fetch_to_decode_instruction[3] ),
    .B_N(\core_pipeline.fetch_to_decode_instruction[6] ),
    .C(\core_pipeline.fetch_to_decode_instruction[4] ),
    .D(_03436_),
    .X(_03636_));
 sky130_fd_sc_hd__or2_4 _06988_ (.A(_03635_),
    .B(_03636_),
    .X(_03637_));
 sky130_fd_sc_hd__a21o_1 _06989_ (.A1(_03322_),
    .A2(_03636_),
    .B1(_03635_),
    .X(_03638_));
 sky130_fd_sc_hd__nor2_1 _06990_ (.A(_03452_),
    .B(_03638_),
    .Y(_03639_));
 sky130_fd_sc_hd__and2_1 _06991_ (.A(net142),
    .B(_03639_),
    .X(_03640_));
 sky130_fd_sc_hd__a221o_1 _06992_ (.A1(net628),
    .A2(net126),
    .B1(_03450_),
    .B2(_03632_),
    .C1(_03640_),
    .X(_00000_));
 sky130_fd_sc_hd__o2111a_1 _06993_ (.A1(\core_pipeline.execute_to_memory_valid ),
    .A2(net458),
    .B1(_03514_),
    .C1(net638),
    .D1(_03430_),
    .X(_00040_));
 sky130_fd_sc_hd__or2_1 _06994_ (.A(\core_pipeline.execute_to_memory_valid ),
    .B(net147),
    .X(_03641_));
 sky130_fd_sc_hd__o211a_1 _06995_ (.A1(\core_pipeline.decode_to_execute_valid ),
    .A2(net133),
    .B1(_03517_),
    .C1(_03641_),
    .X(_00038_));
 sky130_fd_sc_hd__mux2_1 _06996_ (.A0(\core_pipeline.decode_to_execute_valid ),
    .A1(\core_pipeline.fetch_to_decode_valid ),
    .S(net147),
    .X(_03642_));
 sky130_fd_sc_hd__and3_1 _06997_ (.A(_03504_),
    .B(_03517_),
    .C(_03642_),
    .X(_00037_));
 sky130_fd_sc_hd__or4bb_4 _06998_ (.A(\core_pipeline.memory_to_writeback_csr_address[10] ),
    .B(\core_pipeline.memory_to_writeback_csr_address[11] ),
    .C_N(\core_pipeline.memory_to_writeback_csr_address[9] ),
    .D_N(\core_pipeline.memory_to_writeback_csr_address[8] ),
    .X(_03643_));
 sky130_fd_sc_hd__or3b_4 _06999_ (.A(\core_pipeline.memory_to_writeback_csr_address[5] ),
    .B(\core_pipeline.memory_to_writeback_csr_address[4] ),
    .C_N(\core_pipeline.memory_to_writeback_csr_address[6] ),
    .X(_03644_));
 sky130_fd_sc_hd__nor3_4 _07000_ (.A(\core_pipeline.memory_to_writeback_csr_address[7] ),
    .B(_03643_),
    .C(_03644_),
    .Y(_03645_));
 sky130_fd_sc_hd__or2_4 _07001_ (.A(\core_pipeline.memory_to_writeback_csr_address[3] ),
    .B(\core_pipeline.memory_to_writeback_csr_address[2] ),
    .X(_03646_));
 sky130_fd_sc_hd__nor3_4 _07002_ (.A(\core_pipeline.memory_to_writeback_csr_address[1] ),
    .B(_03482_),
    .C(_03646_),
    .Y(_03647_));
 sky130_fd_sc_hd__or3_2 _07003_ (.A(\core_pipeline.memory_to_writeback_csr_address[1] ),
    .B(_03482_),
    .C(_03646_),
    .X(_03648_));
 sky130_fd_sc_hd__and3_4 _07004_ (.A(\core_pipeline.memory_to_writeback_csr_address[0] ),
    .B(_03645_),
    .C(_03647_),
    .X(_03649_));
 sky130_fd_sc_hd__mux2_1 _07005_ (.A0(\core_pipeline.memory_to_writeback_next_pc[0] ),
    .A1(\core_pipeline.csr_to_fetch_mret_vector[0] ),
    .S(net400),
    .X(_03650_));
 sky130_fd_sc_hd__mux2_1 _07006_ (.A0(_03650_),
    .A1(\core_pipeline.memory_to_writeback_alu_data[0] ),
    .S(net237),
    .X(_00005_));
 sky130_fd_sc_hd__mux2_1 _07007_ (.A0(\core_pipeline.memory_to_writeback_next_pc[1] ),
    .A1(\core_pipeline.csr_to_fetch_mret_vector[1] ),
    .S(net400),
    .X(_03651_));
 sky130_fd_sc_hd__mux2_1 _07008_ (.A0(_03651_),
    .A1(\core_pipeline.memory_to_writeback_alu_data[1] ),
    .S(net237),
    .X(_00016_));
 sky130_fd_sc_hd__mux2_1 _07009_ (.A0(\core_pipeline.memory_to_writeback_pc[2] ),
    .A1(\core_pipeline.memory_to_writeback_next_pc[2] ),
    .S(net505),
    .X(_03652_));
 sky130_fd_sc_hd__mux2_1 _07010_ (.A0(_03652_),
    .A1(\core_pipeline.csr_to_fetch_mret_vector[2] ),
    .S(net401),
    .X(_03653_));
 sky130_fd_sc_hd__mux2_1 _07011_ (.A0(_03653_),
    .A1(\core_pipeline.memory_to_writeback_alu_data[2] ),
    .S(net237),
    .X(_00027_));
 sky130_fd_sc_hd__mux2_1 _07012_ (.A0(\core_pipeline.memory_to_writeback_pc[3] ),
    .A1(\core_pipeline.memory_to_writeback_next_pc[3] ),
    .S(net505),
    .X(_03654_));
 sky130_fd_sc_hd__mux2_1 _07013_ (.A0(_03654_),
    .A1(\core_pipeline.csr_to_fetch_mret_vector[3] ),
    .S(net400),
    .X(_03655_));
 sky130_fd_sc_hd__mux2_1 _07014_ (.A0(_03655_),
    .A1(\core_pipeline.memory_to_writeback_alu_data[3] ),
    .S(net237),
    .X(_00030_));
 sky130_fd_sc_hd__mux2_1 _07015_ (.A0(\core_pipeline.memory_to_writeback_pc[4] ),
    .A1(\core_pipeline.memory_to_writeback_next_pc[4] ),
    .S(net505),
    .X(_03656_));
 sky130_fd_sc_hd__mux2_1 _07016_ (.A0(_03656_),
    .A1(\core_pipeline.csr_to_fetch_mret_vector[4] ),
    .S(net400),
    .X(_03657_));
 sky130_fd_sc_hd__mux2_1 _07017_ (.A0(_03657_),
    .A1(\core_pipeline.memory_to_writeback_alu_data[4] ),
    .S(net237),
    .X(_00031_));
 sky130_fd_sc_hd__mux2_1 _07018_ (.A0(\core_pipeline.memory_to_writeback_pc[5] ),
    .A1(\core_pipeline.memory_to_writeback_next_pc[5] ),
    .S(net505),
    .X(_03658_));
 sky130_fd_sc_hd__mux2_1 _07019_ (.A0(_03658_),
    .A1(\core_pipeline.csr_to_fetch_mret_vector[5] ),
    .S(net400),
    .X(_03659_));
 sky130_fd_sc_hd__mux2_1 _07020_ (.A0(_03659_),
    .A1(\core_pipeline.memory_to_writeback_alu_data[5] ),
    .S(net237),
    .X(_00032_));
 sky130_fd_sc_hd__mux2_1 _07021_ (.A0(\core_pipeline.memory_to_writeback_pc[6] ),
    .A1(\core_pipeline.memory_to_writeback_next_pc[6] ),
    .S(net505),
    .X(_03660_));
 sky130_fd_sc_hd__mux2_1 _07022_ (.A0(_03660_),
    .A1(\core_pipeline.csr_to_fetch_mret_vector[6] ),
    .S(net401),
    .X(_03661_));
 sky130_fd_sc_hd__mux2_1 _07023_ (.A0(_03661_),
    .A1(\core_pipeline.memory_to_writeback_alu_data[6] ),
    .S(net237),
    .X(_00033_));
 sky130_fd_sc_hd__mux2_1 _07024_ (.A0(\core_pipeline.memory_to_writeback_pc[7] ),
    .A1(\core_pipeline.memory_to_writeback_next_pc[7] ),
    .S(net505),
    .X(_03662_));
 sky130_fd_sc_hd__mux2_1 _07025_ (.A0(_03662_),
    .A1(\core_pipeline.csr_to_fetch_mret_vector[7] ),
    .S(net401),
    .X(_03663_));
 sky130_fd_sc_hd__mux2_1 _07026_ (.A0(_03663_),
    .A1(\core_pipeline.memory_to_writeback_alu_data[7] ),
    .S(net237),
    .X(_00034_));
 sky130_fd_sc_hd__mux2_1 _07027_ (.A0(\core_pipeline.memory_to_writeback_pc[8] ),
    .A1(\core_pipeline.memory_to_writeback_next_pc[8] ),
    .S(net504),
    .X(_03664_));
 sky130_fd_sc_hd__mux2_1 _07028_ (.A0(_03664_),
    .A1(\core_pipeline.csr_to_fetch_mret_vector[8] ),
    .S(net403),
    .X(_03665_));
 sky130_fd_sc_hd__mux2_1 _07029_ (.A0(_03665_),
    .A1(\core_pipeline.memory_to_writeback_alu_data[8] ),
    .S(net237),
    .X(_00035_));
 sky130_fd_sc_hd__mux2_1 _07030_ (.A0(\core_pipeline.memory_to_writeback_pc[9] ),
    .A1(\core_pipeline.memory_to_writeback_next_pc[9] ),
    .S(net504),
    .X(_03666_));
 sky130_fd_sc_hd__mux2_1 _07031_ (.A0(_03666_),
    .A1(\core_pipeline.csr_to_fetch_mret_vector[9] ),
    .S(net402),
    .X(_03667_));
 sky130_fd_sc_hd__mux2_1 _07032_ (.A0(_03667_),
    .A1(\core_pipeline.memory_to_writeback_alu_data[9] ),
    .S(net238),
    .X(_00036_));
 sky130_fd_sc_hd__mux2_1 _07033_ (.A0(\core_pipeline.memory_to_writeback_pc[10] ),
    .A1(\core_pipeline.memory_to_writeback_next_pc[10] ),
    .S(net504),
    .X(_03668_));
 sky130_fd_sc_hd__mux2_1 _07034_ (.A0(_03668_),
    .A1(\core_pipeline.csr_to_fetch_mret_vector[10] ),
    .S(net402),
    .X(_03669_));
 sky130_fd_sc_hd__mux2_1 _07035_ (.A0(_03669_),
    .A1(\core_pipeline.memory_to_writeback_alu_data[10] ),
    .S(net238),
    .X(_00006_));
 sky130_fd_sc_hd__mux2_1 _07036_ (.A0(\core_pipeline.memory_to_writeback_pc[11] ),
    .A1(\core_pipeline.memory_to_writeback_next_pc[11] ),
    .S(net504),
    .X(_03670_));
 sky130_fd_sc_hd__mux2_1 _07037_ (.A0(_03670_),
    .A1(\core_pipeline.csr_to_fetch_mret_vector[11] ),
    .S(net402),
    .X(_03671_));
 sky130_fd_sc_hd__mux2_1 _07038_ (.A0(_03671_),
    .A1(\core_pipeline.memory_to_writeback_alu_data[11] ),
    .S(net238),
    .X(_00007_));
 sky130_fd_sc_hd__mux2_1 _07039_ (.A0(\core_pipeline.memory_to_writeback_pc[12] ),
    .A1(\core_pipeline.memory_to_writeback_next_pc[12] ),
    .S(net504),
    .X(_03672_));
 sky130_fd_sc_hd__mux2_1 _07040_ (.A0(_03672_),
    .A1(\core_pipeline.csr_to_fetch_mret_vector[12] ),
    .S(net402),
    .X(_03673_));
 sky130_fd_sc_hd__mux2_1 _07041_ (.A0(_03673_),
    .A1(\core_pipeline.memory_to_writeback_alu_data[12] ),
    .S(net238),
    .X(_00008_));
 sky130_fd_sc_hd__mux2_1 _07042_ (.A0(\core_pipeline.memory_to_writeback_pc[13] ),
    .A1(\core_pipeline.memory_to_writeback_next_pc[13] ),
    .S(net504),
    .X(_03674_));
 sky130_fd_sc_hd__mux2_1 _07043_ (.A0(_03674_),
    .A1(\core_pipeline.csr_to_fetch_mret_vector[13] ),
    .S(net402),
    .X(_03675_));
 sky130_fd_sc_hd__mux2_1 _07044_ (.A0(_03675_),
    .A1(\core_pipeline.memory_to_writeback_alu_data[13] ),
    .S(net238),
    .X(_00009_));
 sky130_fd_sc_hd__mux2_1 _07045_ (.A0(\core_pipeline.memory_to_writeback_pc[14] ),
    .A1(\core_pipeline.memory_to_writeback_next_pc[14] ),
    .S(net504),
    .X(_03676_));
 sky130_fd_sc_hd__mux2_1 _07046_ (.A0(_03676_),
    .A1(\core_pipeline.csr_to_fetch_mret_vector[14] ),
    .S(net402),
    .X(_03677_));
 sky130_fd_sc_hd__mux2_1 _07047_ (.A0(_03677_),
    .A1(\core_pipeline.memory_to_writeback_alu_data[14] ),
    .S(net238),
    .X(_00010_));
 sky130_fd_sc_hd__mux2_1 _07048_ (.A0(\core_pipeline.memory_to_writeback_pc[15] ),
    .A1(\core_pipeline.memory_to_writeback_next_pc[15] ),
    .S(net504),
    .X(_03678_));
 sky130_fd_sc_hd__mux2_1 _07049_ (.A0(_03678_),
    .A1(\core_pipeline.csr_to_fetch_mret_vector[15] ),
    .S(net402),
    .X(_03679_));
 sky130_fd_sc_hd__mux2_1 _07050_ (.A0(_03679_),
    .A1(\core_pipeline.memory_to_writeback_alu_data[15] ),
    .S(net238),
    .X(_00011_));
 sky130_fd_sc_hd__mux2_1 _07051_ (.A0(\core_pipeline.memory_to_writeback_pc[16] ),
    .A1(\core_pipeline.memory_to_writeback_next_pc[16] ),
    .S(net504),
    .X(_03680_));
 sky130_fd_sc_hd__mux2_1 _07052_ (.A0(_03680_),
    .A1(\core_pipeline.csr_to_fetch_mret_vector[16] ),
    .S(net402),
    .X(_03681_));
 sky130_fd_sc_hd__mux2_1 _07053_ (.A0(_03681_),
    .A1(\core_pipeline.memory_to_writeback_alu_data[16] ),
    .S(net238),
    .X(_00012_));
 sky130_fd_sc_hd__mux2_1 _07054_ (.A0(\core_pipeline.memory_to_writeback_pc[17] ),
    .A1(\core_pipeline.memory_to_writeback_next_pc[17] ),
    .S(net504),
    .X(_03682_));
 sky130_fd_sc_hd__mux2_1 _07055_ (.A0(_03682_),
    .A1(\core_pipeline.csr_to_fetch_mret_vector[17] ),
    .S(net403),
    .X(_03683_));
 sky130_fd_sc_hd__mux2_1 _07056_ (.A0(_03683_),
    .A1(\core_pipeline.memory_to_writeback_alu_data[17] ),
    .S(net238),
    .X(_00013_));
 sky130_fd_sc_hd__mux2_1 _07057_ (.A0(\core_pipeline.memory_to_writeback_pc[18] ),
    .A1(\core_pipeline.memory_to_writeback_next_pc[18] ),
    .S(net504),
    .X(_03684_));
 sky130_fd_sc_hd__mux2_1 _07058_ (.A0(_03684_),
    .A1(\core_pipeline.csr_to_fetch_mret_vector[18] ),
    .S(net403),
    .X(_03685_));
 sky130_fd_sc_hd__mux2_1 _07059_ (.A0(_03685_),
    .A1(\core_pipeline.memory_to_writeback_alu_data[18] ),
    .S(net238),
    .X(_00014_));
 sky130_fd_sc_hd__mux2_1 _07060_ (.A0(\core_pipeline.memory_to_writeback_pc[19] ),
    .A1(\core_pipeline.memory_to_writeback_next_pc[19] ),
    .S(net504),
    .X(_03686_));
 sky130_fd_sc_hd__mux2_1 _07061_ (.A0(_03686_),
    .A1(\core_pipeline.csr_to_fetch_mret_vector[19] ),
    .S(net402),
    .X(_03687_));
 sky130_fd_sc_hd__mux2_1 _07062_ (.A0(_03687_),
    .A1(\core_pipeline.memory_to_writeback_alu_data[19] ),
    .S(net237),
    .X(_00015_));
 sky130_fd_sc_hd__mux2_1 _07063_ (.A0(\core_pipeline.memory_to_writeback_pc[20] ),
    .A1(\core_pipeline.memory_to_writeback_next_pc[20] ),
    .S(net504),
    .X(_03688_));
 sky130_fd_sc_hd__mux2_1 _07064_ (.A0(_03688_),
    .A1(\core_pipeline.csr_to_fetch_mret_vector[20] ),
    .S(net403),
    .X(_03689_));
 sky130_fd_sc_hd__mux2_1 _07065_ (.A0(_03689_),
    .A1(\core_pipeline.memory_to_writeback_alu_data[20] ),
    .S(net238),
    .X(_00017_));
 sky130_fd_sc_hd__mux2_1 _07066_ (.A0(\core_pipeline.memory_to_writeback_pc[21] ),
    .A1(\core_pipeline.memory_to_writeback_next_pc[21] ),
    .S(net505),
    .X(_03690_));
 sky130_fd_sc_hd__mux2_1 _07067_ (.A0(_03690_),
    .A1(\core_pipeline.csr_to_fetch_mret_vector[21] ),
    .S(net403),
    .X(_03691_));
 sky130_fd_sc_hd__mux2_1 _07068_ (.A0(_03691_),
    .A1(\core_pipeline.memory_to_writeback_alu_data[21] ),
    .S(net238),
    .X(_00018_));
 sky130_fd_sc_hd__mux2_1 _07069_ (.A0(\core_pipeline.memory_to_writeback_pc[22] ),
    .A1(\core_pipeline.memory_to_writeback_next_pc[22] ),
    .S(net504),
    .X(_03692_));
 sky130_fd_sc_hd__mux2_1 _07070_ (.A0(_03692_),
    .A1(\core_pipeline.csr_to_fetch_mret_vector[22] ),
    .S(net403),
    .X(_03693_));
 sky130_fd_sc_hd__mux2_1 _07071_ (.A0(_03693_),
    .A1(\core_pipeline.memory_to_writeback_alu_data[22] ),
    .S(net238),
    .X(_00019_));
 sky130_fd_sc_hd__mux2_2 _07072_ (.A0(\core_pipeline.memory_to_writeback_pc[23] ),
    .A1(\core_pipeline.memory_to_writeback_next_pc[23] ),
    .S(net504),
    .X(_03694_));
 sky130_fd_sc_hd__mux2_1 _07073_ (.A0(_03694_),
    .A1(\core_pipeline.csr_to_fetch_mret_vector[23] ),
    .S(net403),
    .X(_03695_));
 sky130_fd_sc_hd__mux2_1 _07074_ (.A0(_03695_),
    .A1(\core_pipeline.memory_to_writeback_alu_data[23] ),
    .S(net238),
    .X(_00020_));
 sky130_fd_sc_hd__mux2_1 _07075_ (.A0(\core_pipeline.memory_to_writeback_pc[24] ),
    .A1(\core_pipeline.memory_to_writeback_next_pc[24] ),
    .S(net504),
    .X(_03696_));
 sky130_fd_sc_hd__mux2_1 _07076_ (.A0(_03696_),
    .A1(\core_pipeline.csr_to_fetch_mret_vector[24] ),
    .S(net403),
    .X(_03697_));
 sky130_fd_sc_hd__mux2_1 _07077_ (.A0(_03697_),
    .A1(\core_pipeline.memory_to_writeback_alu_data[24] ),
    .S(net238),
    .X(_00021_));
 sky130_fd_sc_hd__mux2_2 _07078_ (.A0(\core_pipeline.memory_to_writeback_pc[25] ),
    .A1(\core_pipeline.memory_to_writeback_next_pc[25] ),
    .S(net504),
    .X(_03698_));
 sky130_fd_sc_hd__mux2_1 _07079_ (.A0(_03698_),
    .A1(\core_pipeline.csr_to_fetch_mret_vector[25] ),
    .S(net403),
    .X(_03699_));
 sky130_fd_sc_hd__mux2_1 _07080_ (.A0(_03699_),
    .A1(\core_pipeline.memory_to_writeback_alu_data[25] ),
    .S(net237),
    .X(_00022_));
 sky130_fd_sc_hd__mux2_1 _07081_ (.A0(\core_pipeline.memory_to_writeback_pc[26] ),
    .A1(\core_pipeline.memory_to_writeback_next_pc[26] ),
    .S(net505),
    .X(_03700_));
 sky130_fd_sc_hd__mux2_1 _07082_ (.A0(_03700_),
    .A1(\core_pipeline.csr_to_fetch_mret_vector[26] ),
    .S(net401),
    .X(_03701_));
 sky130_fd_sc_hd__mux2_1 _07083_ (.A0(_03701_),
    .A1(\core_pipeline.memory_to_writeback_alu_data[26] ),
    .S(net237),
    .X(_00023_));
 sky130_fd_sc_hd__mux2_1 _07084_ (.A0(\core_pipeline.memory_to_writeback_pc[27] ),
    .A1(\core_pipeline.memory_to_writeback_next_pc[27] ),
    .S(net505),
    .X(_03702_));
 sky130_fd_sc_hd__mux2_1 _07085_ (.A0(_03702_),
    .A1(\core_pipeline.csr_to_fetch_mret_vector[27] ),
    .S(net401),
    .X(_03703_));
 sky130_fd_sc_hd__mux2_1 _07086_ (.A0(_03703_),
    .A1(\core_pipeline.memory_to_writeback_alu_data[27] ),
    .S(net237),
    .X(_00024_));
 sky130_fd_sc_hd__mux2_1 _07087_ (.A0(\core_pipeline.memory_to_writeback_pc[28] ),
    .A1(\core_pipeline.memory_to_writeback_next_pc[28] ),
    .S(net505),
    .X(_03704_));
 sky130_fd_sc_hd__mux2_1 _07088_ (.A0(_03704_),
    .A1(\core_pipeline.csr_to_fetch_mret_vector[28] ),
    .S(net401),
    .X(_03705_));
 sky130_fd_sc_hd__mux2_1 _07089_ (.A0(_03705_),
    .A1(\core_pipeline.memory_to_writeback_alu_data[28] ),
    .S(net237),
    .X(_00025_));
 sky130_fd_sc_hd__mux2_1 _07090_ (.A0(\core_pipeline.memory_to_writeback_pc[29] ),
    .A1(\core_pipeline.memory_to_writeback_next_pc[29] ),
    .S(net505),
    .X(_03706_));
 sky130_fd_sc_hd__mux2_1 _07091_ (.A0(_03706_),
    .A1(\core_pipeline.csr_to_fetch_mret_vector[29] ),
    .S(net401),
    .X(_03707_));
 sky130_fd_sc_hd__mux2_1 _07092_ (.A0(_03707_),
    .A1(\core_pipeline.memory_to_writeback_alu_data[29] ),
    .S(net237),
    .X(_00026_));
 sky130_fd_sc_hd__mux2_2 _07093_ (.A0(\core_pipeline.memory_to_writeback_pc[30] ),
    .A1(\core_pipeline.memory_to_writeback_next_pc[30] ),
    .S(net505),
    .X(_03708_));
 sky130_fd_sc_hd__mux2_1 _07094_ (.A0(_03708_),
    .A1(\core_pipeline.csr_to_fetch_mret_vector[30] ),
    .S(net401),
    .X(_03709_));
 sky130_fd_sc_hd__mux2_1 _07095_ (.A0(_03709_),
    .A1(\core_pipeline.memory_to_writeback_alu_data[30] ),
    .S(net237),
    .X(_00028_));
 sky130_fd_sc_hd__mux2_1 _07096_ (.A0(\core_pipeline.memory_to_writeback_pc[31] ),
    .A1(\core_pipeline.memory_to_writeback_next_pc[31] ),
    .S(net505),
    .X(_03710_));
 sky130_fd_sc_hd__mux2_1 _07097_ (.A0(_03710_),
    .A1(\core_pipeline.csr_to_fetch_mret_vector[31] ),
    .S(net400),
    .X(_03711_));
 sky130_fd_sc_hd__mux2_1 _07098_ (.A0(_03711_),
    .A1(\core_pipeline.memory_to_writeback_alu_data[31] ),
    .S(net237),
    .X(_00029_));
 sky130_fd_sc_hd__and4b_4 _07099_ (.A_N(\core_pipeline.execute_to_memory_exception ),
    .B(\core_pipeline.execute_to_memory_valid ),
    .C(\core_pipeline.execute_to_memory_store ),
    .D(_03426_),
    .X(_03712_));
 sky130_fd_sc_hd__and2b_4 _07100_ (.A_N(net492),
    .B(net275),
    .X(_03713_));
 sky130_fd_sc_hd__and2_4 _07101_ (.A(_03509_),
    .B(net275),
    .X(net99));
 sky130_fd_sc_hd__or2_1 _07102_ (.A(\core_busio.mem_address[0] ),
    .B(_03424_),
    .X(_03714_));
 sky130_fd_sc_hd__and2_4 _07103_ (.A(_03713_),
    .B(_03714_),
    .X(net100));
 sky130_fd_sc_hd__and3b_4 _07104_ (.A_N(net493),
    .B(net275),
    .C(net492),
    .X(_03715_));
 sky130_fd_sc_hd__a21o_4 _07105_ (.A1(\core_busio.mem_size[1] ),
    .A2(net275),
    .B1(_03715_),
    .X(net101));
 sky130_fd_sc_hd__nand2_1 _07106_ (.A(\core_busio.mem_size[1] ),
    .B(\core_busio.mem_size[0] ),
    .Y(_03716_));
 sky130_fd_sc_hd__o2111a_4 _07107_ (.A1(\core_busio.mem_size[1] ),
    .A2(net490),
    .B1(net275),
    .C1(_03714_),
    .D1(_03716_),
    .X(net102));
 sky130_fd_sc_hd__and3_4 _07108_ (.A(\core_busio.mem_store_data[0] ),
    .B(_03509_),
    .C(net275),
    .X(net67));
 sky130_fd_sc_hd__and3_4 _07109_ (.A(\core_busio.mem_store_data[1] ),
    .B(_03509_),
    .C(net275),
    .X(net78));
 sky130_fd_sc_hd__and3_4 _07110_ (.A(\core_busio.mem_store_data[2] ),
    .B(_03509_),
    .C(net275),
    .X(net89));
 sky130_fd_sc_hd__and3_4 _07111_ (.A(\core_busio.mem_store_data[3] ),
    .B(_03509_),
    .C(net275),
    .X(net92));
 sky130_fd_sc_hd__and3_2 _07112_ (.A(\core_busio.mem_store_data[4] ),
    .B(_03509_),
    .C(net275),
    .X(net93));
 sky130_fd_sc_hd__and3_4 _07113_ (.A(\core_busio.mem_store_data[5] ),
    .B(_03509_),
    .C(_03712_),
    .X(net94));
 sky130_fd_sc_hd__and3_4 _07114_ (.A(\core_busio.mem_store_data[6] ),
    .B(_03509_),
    .C(_03712_),
    .X(net95));
 sky130_fd_sc_hd__and3_4 _07115_ (.A(\core_busio.mem_store_data[7] ),
    .B(_03509_),
    .C(net275),
    .X(net96));
 sky130_fd_sc_hd__mux2_1 _07116_ (.A0(\core_busio.mem_store_data[8] ),
    .A1(\core_busio.mem_store_data[0] ),
    .S(net493),
    .X(_03717_));
 sky130_fd_sc_hd__and2_2 _07117_ (.A(_03713_),
    .B(_03717_),
    .X(net97));
 sky130_fd_sc_hd__mux2_1 _07118_ (.A0(\core_busio.mem_store_data[9] ),
    .A1(\core_busio.mem_store_data[1] ),
    .S(net494),
    .X(_03718_));
 sky130_fd_sc_hd__and2_4 _07119_ (.A(_03713_),
    .B(_03718_),
    .X(net98));
 sky130_fd_sc_hd__mux2_1 _07120_ (.A0(\core_busio.mem_store_data[10] ),
    .A1(\core_busio.mem_store_data[2] ),
    .S(net493),
    .X(_03719_));
 sky130_fd_sc_hd__and2_2 _07121_ (.A(_03713_),
    .B(_03719_),
    .X(net68));
 sky130_fd_sc_hd__mux2_1 _07122_ (.A0(\core_busio.mem_store_data[11] ),
    .A1(\core_busio.mem_store_data[3] ),
    .S(net493),
    .X(_03720_));
 sky130_fd_sc_hd__and2_2 _07123_ (.A(_03713_),
    .B(_03720_),
    .X(net69));
 sky130_fd_sc_hd__mux2_1 _07124_ (.A0(\core_busio.mem_store_data[12] ),
    .A1(\core_busio.mem_store_data[4] ),
    .S(net494),
    .X(_03721_));
 sky130_fd_sc_hd__and2_4 _07125_ (.A(_03713_),
    .B(_03721_),
    .X(net70));
 sky130_fd_sc_hd__mux2_1 _07126_ (.A0(\core_busio.mem_store_data[13] ),
    .A1(\core_busio.mem_store_data[5] ),
    .S(net495),
    .X(_03722_));
 sky130_fd_sc_hd__and2_4 _07127_ (.A(_03713_),
    .B(_03722_),
    .X(net71));
 sky130_fd_sc_hd__mux2_1 _07128_ (.A0(\core_busio.mem_store_data[14] ),
    .A1(\core_busio.mem_store_data[6] ),
    .S(net494),
    .X(_03723_));
 sky130_fd_sc_hd__and2_4 _07129_ (.A(_03713_),
    .B(_03723_),
    .X(net72));
 sky130_fd_sc_hd__mux2_1 _07130_ (.A0(\core_busio.mem_store_data[15] ),
    .A1(\core_busio.mem_store_data[7] ),
    .S(net495),
    .X(_03724_));
 sky130_fd_sc_hd__and2_4 _07131_ (.A(_03713_),
    .B(_03724_),
    .X(net73));
 sky130_fd_sc_hd__mux2_1 _07132_ (.A0(\core_busio.mem_store_data[16] ),
    .A1(\core_busio.mem_store_data[8] ),
    .S(net493),
    .X(_03725_));
 sky130_fd_sc_hd__a22o_4 _07133_ (.A1(\core_busio.mem_store_data[0] ),
    .A2(_03715_),
    .B1(_03725_),
    .B2(_03713_),
    .X(net74));
 sky130_fd_sc_hd__mux2_1 _07134_ (.A0(\core_busio.mem_store_data[17] ),
    .A1(\core_busio.mem_store_data[9] ),
    .S(net493),
    .X(_03726_));
 sky130_fd_sc_hd__a22o_4 _07135_ (.A1(\core_busio.mem_store_data[1] ),
    .A2(_03715_),
    .B1(_03726_),
    .B2(_03713_),
    .X(net75));
 sky130_fd_sc_hd__mux2_1 _07136_ (.A0(\core_busio.mem_store_data[18] ),
    .A1(\core_busio.mem_store_data[10] ),
    .S(net493),
    .X(_03727_));
 sky130_fd_sc_hd__a22o_2 _07137_ (.A1(\core_busio.mem_store_data[2] ),
    .A2(_03715_),
    .B1(_03727_),
    .B2(_03713_),
    .X(net76));
 sky130_fd_sc_hd__mux2_1 _07138_ (.A0(\core_busio.mem_store_data[19] ),
    .A1(\core_busio.mem_store_data[11] ),
    .S(net493),
    .X(_03728_));
 sky130_fd_sc_hd__a22o_4 _07139_ (.A1(\core_busio.mem_store_data[3] ),
    .A2(_03715_),
    .B1(_03728_),
    .B2(_03713_),
    .X(net77));
 sky130_fd_sc_hd__mux2_1 _07140_ (.A0(\core_busio.mem_store_data[20] ),
    .A1(\core_busio.mem_store_data[12] ),
    .S(net493),
    .X(_03729_));
 sky130_fd_sc_hd__a22o_4 _07141_ (.A1(\core_busio.mem_store_data[4] ),
    .A2(_03715_),
    .B1(_03729_),
    .B2(_03713_),
    .X(net79));
 sky130_fd_sc_hd__mux2_1 _07142_ (.A0(\core_busio.mem_store_data[21] ),
    .A1(\core_busio.mem_store_data[13] ),
    .S(net495),
    .X(_03730_));
 sky130_fd_sc_hd__a22o_4 _07143_ (.A1(\core_busio.mem_store_data[5] ),
    .A2(_03715_),
    .B1(_03730_),
    .B2(_03713_),
    .X(net80));
 sky130_fd_sc_hd__mux2_1 _07144_ (.A0(\core_busio.mem_store_data[22] ),
    .A1(\core_busio.mem_store_data[14] ),
    .S(net494),
    .X(_03731_));
 sky130_fd_sc_hd__a22o_4 _07145_ (.A1(\core_busio.mem_store_data[6] ),
    .A2(_03715_),
    .B1(_03731_),
    .B2(_03713_),
    .X(net81));
 sky130_fd_sc_hd__mux2_1 _07146_ (.A0(\core_busio.mem_store_data[23] ),
    .A1(\core_busio.mem_store_data[15] ),
    .S(net493),
    .X(_03732_));
 sky130_fd_sc_hd__a22o_4 _07147_ (.A1(\core_busio.mem_store_data[7] ),
    .A2(_03715_),
    .B1(_03732_),
    .B2(_03713_),
    .X(net82));
 sky130_fd_sc_hd__mux4_1 _07148_ (.A0(\core_busio.mem_store_data[24] ),
    .A1(\core_busio.mem_store_data[16] ),
    .A2(\core_busio.mem_store_data[8] ),
    .A3(\core_busio.mem_store_data[0] ),
    .S0(net493),
    .S1(net492),
    .X(_03733_));
 sky130_fd_sc_hd__and2_4 _07149_ (.A(net275),
    .B(_03733_),
    .X(net83));
 sky130_fd_sc_hd__mux4_1 _07150_ (.A0(\core_busio.mem_store_data[25] ),
    .A1(\core_busio.mem_store_data[17] ),
    .A2(\core_busio.mem_store_data[9] ),
    .A3(\core_busio.mem_store_data[1] ),
    .S0(net493),
    .S1(net492),
    .X(_03734_));
 sky130_fd_sc_hd__and2_4 _07151_ (.A(net275),
    .B(_03734_),
    .X(net84));
 sky130_fd_sc_hd__mux4_1 _07152_ (.A0(\core_busio.mem_store_data[26] ),
    .A1(\core_busio.mem_store_data[18] ),
    .A2(\core_busio.mem_store_data[10] ),
    .A3(\core_busio.mem_store_data[2] ),
    .S0(net493),
    .S1(net492),
    .X(_03735_));
 sky130_fd_sc_hd__and2_4 _07153_ (.A(net275),
    .B(_03735_),
    .X(net85));
 sky130_fd_sc_hd__mux4_2 _07154_ (.A0(\core_busio.mem_store_data[27] ),
    .A1(\core_busio.mem_store_data[19] ),
    .A2(\core_busio.mem_store_data[11] ),
    .A3(\core_busio.mem_store_data[3] ),
    .S0(net493),
    .S1(net492),
    .X(_03736_));
 sky130_fd_sc_hd__and2_4 _07155_ (.A(_03712_),
    .B(_03736_),
    .X(net86));
 sky130_fd_sc_hd__mux4_1 _07156_ (.A0(\core_busio.mem_store_data[28] ),
    .A1(\core_busio.mem_store_data[20] ),
    .A2(\core_busio.mem_store_data[12] ),
    .A3(\core_busio.mem_store_data[4] ),
    .S0(net494),
    .S1(net492),
    .X(_03737_));
 sky130_fd_sc_hd__and2_2 _07157_ (.A(_03712_),
    .B(_03737_),
    .X(net87));
 sky130_fd_sc_hd__mux4_1 _07158_ (.A0(\core_busio.mem_store_data[29] ),
    .A1(\core_busio.mem_store_data[21] ),
    .A2(\core_busio.mem_store_data[13] ),
    .A3(\core_busio.mem_store_data[5] ),
    .S0(net495),
    .S1(net490),
    .X(_03738_));
 sky130_fd_sc_hd__and2_4 _07159_ (.A(net275),
    .B(_03738_),
    .X(net88));
 sky130_fd_sc_hd__mux4_1 _07160_ (.A0(\core_busio.mem_store_data[30] ),
    .A1(\core_busio.mem_store_data[22] ),
    .A2(\core_busio.mem_store_data[14] ),
    .A3(\core_busio.mem_store_data[6] ),
    .S0(net494),
    .S1(net492),
    .X(_03739_));
 sky130_fd_sc_hd__and2_4 _07161_ (.A(net275),
    .B(_03739_),
    .X(net90));
 sky130_fd_sc_hd__mux4_1 _07162_ (.A0(\core_busio.mem_store_data[31] ),
    .A1(\core_busio.mem_store_data[23] ),
    .A2(\core_busio.mem_store_data[15] ),
    .A3(\core_busio.mem_store_data[7] ),
    .S0(net493),
    .S1(net490),
    .X(_03740_));
 sky130_fd_sc_hd__and2_4 _07163_ (.A(net275),
    .B(_03740_),
    .X(net91));
 sky130_fd_sc_hd__mux2_8 _07164_ (.A0(\core_pipeline.pipeline_fetch.pc[2] ),
    .A1(\core_busio.mem_address[2] ),
    .S(net262),
    .X(net56));
 sky130_fd_sc_hd__mux2_4 _07165_ (.A0(\core_pipeline.pipeline_fetch.pc[3] ),
    .A1(\core_busio.mem_address[3] ),
    .S(net262),
    .X(net59));
 sky130_fd_sc_hd__mux2_4 _07166_ (.A0(\core_pipeline.pipeline_fetch.pc[4] ),
    .A1(\core_busio.mem_address[4] ),
    .S(net262),
    .X(net60));
 sky130_fd_sc_hd__mux2_8 _07167_ (.A0(\core_pipeline.pipeline_fetch.pc[5] ),
    .A1(\core_busio.mem_address[5] ),
    .S(net262),
    .X(net61));
 sky130_fd_sc_hd__mux2_8 _07168_ (.A0(\core_pipeline.pipeline_fetch.pc[6] ),
    .A1(\core_busio.mem_address[6] ),
    .S(net262),
    .X(net62));
 sky130_fd_sc_hd__mux2_8 _07169_ (.A0(\core_pipeline.pipeline_fetch.pc[7] ),
    .A1(\core_busio.mem_address[7] ),
    .S(net262),
    .X(net63));
 sky130_fd_sc_hd__mux2_8 _07170_ (.A0(\core_pipeline.pipeline_fetch.pc[8] ),
    .A1(\core_busio.mem_address[8] ),
    .S(net261),
    .X(net64));
 sky130_fd_sc_hd__mux2_8 _07171_ (.A0(\core_pipeline.pipeline_fetch.pc[9] ),
    .A1(\core_busio.mem_address[9] ),
    .S(net261),
    .X(net65));
 sky130_fd_sc_hd__mux2_8 _07172_ (.A0(\core_pipeline.pipeline_fetch.pc[10] ),
    .A1(\core_busio.mem_address[10] ),
    .S(net261),
    .X(net36));
 sky130_fd_sc_hd__mux2_8 _07173_ (.A0(\core_pipeline.pipeline_fetch.pc[11] ),
    .A1(\core_busio.mem_address[11] ),
    .S(net261),
    .X(net37));
 sky130_fd_sc_hd__mux2_8 _07174_ (.A0(\core_pipeline.pipeline_fetch.pc[12] ),
    .A1(\core_busio.mem_address[12] ),
    .S(net261),
    .X(net38));
 sky130_fd_sc_hd__mux2_1 _07175_ (.A0(\core_pipeline.pipeline_fetch.pc[13] ),
    .A1(\core_busio.mem_address[13] ),
    .S(net262),
    .X(net39));
 sky130_fd_sc_hd__mux2_2 _07176_ (.A0(\core_pipeline.pipeline_fetch.pc[14] ),
    .A1(\core_busio.mem_address[14] ),
    .S(net261),
    .X(net40));
 sky130_fd_sc_hd__mux2_8 _07177_ (.A0(\core_pipeline.pipeline_fetch.pc[15] ),
    .A1(\core_busio.mem_address[15] ),
    .S(net261),
    .X(net41));
 sky130_fd_sc_hd__mux2_8 _07178_ (.A0(\core_pipeline.pipeline_fetch.pc[16] ),
    .A1(\core_busio.mem_address[16] ),
    .S(net261),
    .X(net42));
 sky130_fd_sc_hd__mux2_8 _07179_ (.A0(\core_pipeline.pipeline_fetch.pc[17] ),
    .A1(\core_busio.mem_address[17] ),
    .S(net261),
    .X(net43));
 sky130_fd_sc_hd__mux2_8 _07180_ (.A0(\core_pipeline.pipeline_fetch.pc[18] ),
    .A1(\core_busio.mem_address[18] ),
    .S(net261),
    .X(net44));
 sky130_fd_sc_hd__mux2_8 _07181_ (.A0(\core_pipeline.pipeline_fetch.pc[19] ),
    .A1(\core_busio.mem_address[19] ),
    .S(net261),
    .X(net45));
 sky130_fd_sc_hd__mux2_8 _07182_ (.A0(\core_pipeline.pipeline_fetch.pc[20] ),
    .A1(\core_busio.mem_address[20] ),
    .S(net261),
    .X(net46));
 sky130_fd_sc_hd__mux2_8 _07183_ (.A0(\core_pipeline.pipeline_fetch.pc[21] ),
    .A1(\core_busio.mem_address[21] ),
    .S(net262),
    .X(net47));
 sky130_fd_sc_hd__mux2_8 _07184_ (.A0(\core_pipeline.pipeline_fetch.pc[22] ),
    .A1(\core_busio.mem_address[22] ),
    .S(net261),
    .X(net48));
 sky130_fd_sc_hd__mux2_2 _07185_ (.A0(\core_pipeline.pipeline_fetch.pc[23] ),
    .A1(\core_busio.mem_address[23] ),
    .S(net262),
    .X(net49));
 sky130_fd_sc_hd__mux2_4 _07186_ (.A0(\core_pipeline.pipeline_fetch.pc[24] ),
    .A1(\core_busio.mem_address[24] ),
    .S(net261),
    .X(net50));
 sky130_fd_sc_hd__mux2_2 _07187_ (.A0(\core_pipeline.pipeline_fetch.pc[25] ),
    .A1(\core_busio.mem_address[25] ),
    .S(net261),
    .X(net51));
 sky130_fd_sc_hd__mux2_8 _07188_ (.A0(\core_pipeline.pipeline_fetch.pc[26] ),
    .A1(\core_busio.mem_address[26] ),
    .S(net261),
    .X(net52));
 sky130_fd_sc_hd__mux2_2 _07189_ (.A0(\core_pipeline.pipeline_fetch.pc[27] ),
    .A1(\core_busio.mem_address[27] ),
    .S(net262),
    .X(net53));
 sky130_fd_sc_hd__mux2_8 _07190_ (.A0(\core_pipeline.pipeline_fetch.pc[28] ),
    .A1(\core_busio.mem_address[28] ),
    .S(net262),
    .X(net54));
 sky130_fd_sc_hd__mux2_4 _07191_ (.A0(\core_pipeline.pipeline_fetch.pc[29] ),
    .A1(\core_busio.mem_address[29] ),
    .S(net262),
    .X(net55));
 sky130_fd_sc_hd__mux2_8 _07192_ (.A0(\core_pipeline.pipeline_fetch.pc[30] ),
    .A1(\core_busio.mem_address[30] ),
    .S(net262),
    .X(net57));
 sky130_fd_sc_hd__mux2_8 _07193_ (.A0(\core_pipeline.pipeline_fetch.pc[31] ),
    .A1(\core_busio.mem_address[31] ),
    .S(net262),
    .X(net58));
 sky130_fd_sc_hd__mux2_8 _07194_ (.A0(\core_pipeline.decode_to_execute_rs2_data[31] ),
    .A1(\core_pipeline.decode_to_execute_rs2_bypass[31] ),
    .S(net487),
    .X(_03741_));
 sky130_fd_sc_hd__inv_2 _07195_ (.A(_03741_),
    .Y(_03742_));
 sky130_fd_sc_hd__mux2_8 _07196_ (.A0(\core_pipeline.decode_to_execute_rs1_data[31] ),
    .A1(\core_pipeline.decode_to_execute_rs1_bypass[31] ),
    .S(net489),
    .X(_03743_));
 sky130_fd_sc_hd__xor2_1 _07197_ (.A(_03741_),
    .B(_03743_),
    .X(_03744_));
 sky130_fd_sc_hd__a21bo_1 _07198_ (.A1(_03422_),
    .A2(_03744_),
    .B1_N(\core_pipeline.decode_to_execute_cmp_function[2] ),
    .X(_03745_));
 sky130_fd_sc_hd__mux2_8 _07199_ (.A0(\core_pipeline.decode_to_execute_rs2_data[29] ),
    .A1(\core_pipeline.decode_to_execute_rs2_bypass[29] ),
    .S(net487),
    .X(_03746_));
 sky130_fd_sc_hd__mux2_8 _07200_ (.A0(\core_pipeline.decode_to_execute_rs1_data[29] ),
    .A1(\core_pipeline.decode_to_execute_rs1_bypass[29] ),
    .S(net489),
    .X(_03747_));
 sky130_fd_sc_hd__inv_2 _07201_ (.A(_03747_),
    .Y(_03748_));
 sky130_fd_sc_hd__mux2_8 _07202_ (.A0(\core_pipeline.decode_to_execute_rs2_data[28] ),
    .A1(\core_pipeline.decode_to_execute_rs2_bypass[28] ),
    .S(net487),
    .X(_03749_));
 sky130_fd_sc_hd__mux2_8 _07203_ (.A0(\core_pipeline.decode_to_execute_rs1_data[28] ),
    .A1(\core_pipeline.decode_to_execute_rs1_bypass[28] ),
    .S(net489),
    .X(_03750_));
 sky130_fd_sc_hd__inv_2 _07204_ (.A(_03750_),
    .Y(_03751_));
 sky130_fd_sc_hd__a22o_1 _07205_ (.A1(_03746_),
    .A2(_03748_),
    .B1(_03749_),
    .B2(_03751_),
    .X(_03752_));
 sky130_fd_sc_hd__mux2_8 _07206_ (.A0(\core_pipeline.decode_to_execute_rs2_data[25] ),
    .A1(\core_pipeline.decode_to_execute_rs2_bypass[25] ),
    .S(net486),
    .X(_03753_));
 sky130_fd_sc_hd__mux2_4 _07207_ (.A0(\core_pipeline.decode_to_execute_rs1_data[25] ),
    .A1(\core_pipeline.decode_to_execute_rs1_bypass[25] ),
    .S(net488),
    .X(_03754_));
 sky130_fd_sc_hd__inv_2 _07208_ (.A(_03754_),
    .Y(_03755_));
 sky130_fd_sc_hd__mux2_8 _07209_ (.A0(\core_pipeline.decode_to_execute_rs2_data[26] ),
    .A1(\core_pipeline.decode_to_execute_rs2_bypass[26] ),
    .S(net486),
    .X(_03756_));
 sky130_fd_sc_hd__inv_2 _07210_ (.A(_03756_),
    .Y(_03757_));
 sky130_fd_sc_hd__mux2_4 _07211_ (.A0(\core_pipeline.decode_to_execute_rs1_data[26] ),
    .A1(\core_pipeline.decode_to_execute_rs1_bypass[26] ),
    .S(net488),
    .X(_03758_));
 sky130_fd_sc_hd__a2bb2o_1 _07212_ (.A1_N(_03753_),
    .A2_N(_03755_),
    .B1(_03757_),
    .B2(_03758_),
    .X(_03759_));
 sky130_fd_sc_hd__mux2_8 _07213_ (.A0(\core_pipeline.decode_to_execute_rs2_data[27] ),
    .A1(\core_pipeline.decode_to_execute_rs2_bypass[27] ),
    .S(net487),
    .X(_03760_));
 sky130_fd_sc_hd__mux2_8 _07214_ (.A0(\core_pipeline.decode_to_execute_rs1_data[27] ),
    .A1(\core_pipeline.decode_to_execute_rs1_bypass[27] ),
    .S(net489),
    .X(_03761_));
 sky130_fd_sc_hd__inv_2 _07215_ (.A(_03761_),
    .Y(_03762_));
 sky130_fd_sc_hd__o22a_1 _07216_ (.A1(_03749_),
    .A2(_03751_),
    .B1(_03760_),
    .B2(_03762_),
    .X(_03763_));
 sky130_fd_sc_hd__o2bb2a_1 _07217_ (.A1_N(_03762_),
    .A2_N(_03760_),
    .B1(_03758_),
    .B2(_03757_),
    .X(_03764_));
 sky130_fd_sc_hd__inv_2 _07218_ (.A(_03764_),
    .Y(_03765_));
 sky130_fd_sc_hd__mux2_8 _07219_ (.A0(\core_pipeline.decode_to_execute_rs2_data[24] ),
    .A1(\core_pipeline.decode_to_execute_rs2_bypass[24] ),
    .S(net486),
    .X(_03766_));
 sky130_fd_sc_hd__mux2_8 _07220_ (.A0(\core_pipeline.decode_to_execute_rs1_data[24] ),
    .A1(\core_pipeline.decode_to_execute_rs1_bypass[24] ),
    .S(net488),
    .X(_03767_));
 sky130_fd_sc_hd__inv_2 _07221_ (.A(_03767_),
    .Y(_03768_));
 sky130_fd_sc_hd__a221o_1 _07222_ (.A1(_03753_),
    .A2(_03755_),
    .B1(_03766_),
    .B2(_03768_),
    .C1(_03765_),
    .X(_03769_));
 sky130_fd_sc_hd__mux2_8 _07223_ (.A0(\core_pipeline.decode_to_execute_rs1_data[30] ),
    .A1(\core_pipeline.decode_to_execute_rs1_bypass[30] ),
    .S(net488),
    .X(_03770_));
 sky130_fd_sc_hd__mux2_8 _07224_ (.A0(\core_pipeline.decode_to_execute_rs2_data[30] ),
    .A1(\core_pipeline.decode_to_execute_rs2_bypass[30] ),
    .S(\core_pipeline.decode_to_execute_rs2_bypassed ),
    .X(_03771_));
 sky130_fd_sc_hd__inv_2 _07225_ (.A(_03771_),
    .Y(_03772_));
 sky130_fd_sc_hd__a21o_1 _07226_ (.A1(_03770_),
    .A2(_03772_),
    .B1(_03744_),
    .X(_03773_));
 sky130_fd_sc_hd__nor2_1 _07227_ (.A(_03770_),
    .B(_03772_),
    .Y(_03774_));
 sky130_fd_sc_hd__or2_1 _07228_ (.A(_03746_),
    .B(_03748_),
    .X(_03775_));
 sky130_fd_sc_hd__o22a_1 _07229_ (.A1(_03766_),
    .A2(_03768_),
    .B1(_03770_),
    .B2(_03772_),
    .X(_03776_));
 sky130_fd_sc_hd__and4b_1 _07230_ (.A_N(_03752_),
    .B(_03763_),
    .C(_03775_),
    .D(_03776_),
    .X(_03777_));
 sky130_fd_sc_hd__or4b_1 _07231_ (.A(_03759_),
    .B(_03769_),
    .C(_03773_),
    .D_N(_03777_),
    .X(_03778_));
 sky130_fd_sc_hd__mux2_8 _07232_ (.A0(\core_pipeline.decode_to_execute_rs2_data[23] ),
    .A1(\core_pipeline.decode_to_execute_rs2_bypass[23] ),
    .S(\core_pipeline.decode_to_execute_rs2_bypassed ),
    .X(_03779_));
 sky130_fd_sc_hd__inv_2 _07233_ (.A(_03779_),
    .Y(_03780_));
 sky130_fd_sc_hd__mux2_8 _07234_ (.A0(\core_pipeline.decode_to_execute_rs1_data[23] ),
    .A1(\core_pipeline.decode_to_execute_rs1_bypass[23] ),
    .S(net489),
    .X(_03781_));
 sky130_fd_sc_hd__and2_1 _07235_ (.A(_03780_),
    .B(_03781_),
    .X(_03782_));
 sky130_fd_sc_hd__mux2_8 _07236_ (.A0(\core_pipeline.decode_to_execute_rs2_data[22] ),
    .A1(\core_pipeline.decode_to_execute_rs2_bypass[22] ),
    .S(net487),
    .X(_03783_));
 sky130_fd_sc_hd__inv_2 _07237_ (.A(_03783_),
    .Y(_03784_));
 sky130_fd_sc_hd__mux2_8 _07238_ (.A0(\core_pipeline.decode_to_execute_rs1_data[22] ),
    .A1(\core_pipeline.decode_to_execute_rs1_bypass[22] ),
    .S(net489),
    .X(_03785_));
 sky130_fd_sc_hd__mux2_8 _07239_ (.A0(\core_pipeline.decode_to_execute_rs2_data[20] ),
    .A1(\core_pipeline.decode_to_execute_rs2_bypass[20] ),
    .S(net487),
    .X(_03786_));
 sky130_fd_sc_hd__mux2_8 _07240_ (.A0(\core_pipeline.decode_to_execute_rs1_data[20] ),
    .A1(\core_pipeline.decode_to_execute_rs1_bypass[20] ),
    .S(net489),
    .X(_03787_));
 sky130_fd_sc_hd__inv_2 _07241_ (.A(_03787_),
    .Y(_03788_));
 sky130_fd_sc_hd__mux2_8 _07242_ (.A0(\core_pipeline.decode_to_execute_rs2_data[21] ),
    .A1(\core_pipeline.decode_to_execute_rs2_bypass[21] ),
    .S(net487),
    .X(_03789_));
 sky130_fd_sc_hd__mux2_8 _07243_ (.A0(\core_pipeline.decode_to_execute_rs1_data[21] ),
    .A1(\core_pipeline.decode_to_execute_rs1_bypass[21] ),
    .S(net489),
    .X(_03790_));
 sky130_fd_sc_hd__inv_2 _07244_ (.A(_03790_),
    .Y(_03791_));
 sky130_fd_sc_hd__a22o_1 _07245_ (.A1(_03786_),
    .A2(_03788_),
    .B1(_03789_),
    .B2(_03791_),
    .X(_03792_));
 sky130_fd_sc_hd__mux2_8 _07246_ (.A0(\core_pipeline.decode_to_execute_rs2_data[18] ),
    .A1(\core_pipeline.decode_to_execute_rs2_bypass[18] ),
    .S(net487),
    .X(_03793_));
 sky130_fd_sc_hd__mux2_8 _07247_ (.A0(\core_pipeline.decode_to_execute_rs1_data[18] ),
    .A1(\core_pipeline.decode_to_execute_rs1_bypass[18] ),
    .S(net489),
    .X(_03794_));
 sky130_fd_sc_hd__inv_2 _07248_ (.A(_03794_),
    .Y(_03795_));
 sky130_fd_sc_hd__mux2_8 _07249_ (.A0(\core_pipeline.decode_to_execute_rs2_data[19] ),
    .A1(\core_pipeline.decode_to_execute_rs2_bypass[19] ),
    .S(net487),
    .X(_03796_));
 sky130_fd_sc_hd__mux2_8 _07250_ (.A0(\core_pipeline.decode_to_execute_rs1_data[19] ),
    .A1(\core_pipeline.decode_to_execute_rs1_bypass[19] ),
    .S(net489),
    .X(_03797_));
 sky130_fd_sc_hd__inv_2 _07251_ (.A(_03797_),
    .Y(_03798_));
 sky130_fd_sc_hd__a22o_1 _07252_ (.A1(_03793_),
    .A2(_03795_),
    .B1(_03796_),
    .B2(_03798_),
    .X(_03799_));
 sky130_fd_sc_hd__mux2_8 _07253_ (.A0(\core_pipeline.decode_to_execute_rs2_data[17] ),
    .A1(\core_pipeline.decode_to_execute_rs2_bypass[17] ),
    .S(net487),
    .X(_03800_));
 sky130_fd_sc_hd__mux2_8 _07254_ (.A0(\core_pipeline.decode_to_execute_rs1_data[17] ),
    .A1(\core_pipeline.decode_to_execute_rs1_bypass[17] ),
    .S(net489),
    .X(_03801_));
 sky130_fd_sc_hd__inv_2 _07255_ (.A(_03801_),
    .Y(_03802_));
 sky130_fd_sc_hd__mux2_8 _07256_ (.A0(\core_pipeline.decode_to_execute_rs2_data[16] ),
    .A1(\core_pipeline.decode_to_execute_rs2_bypass[16] ),
    .S(net486),
    .X(_03803_));
 sky130_fd_sc_hd__mux2_8 _07257_ (.A0(\core_pipeline.decode_to_execute_rs1_data[16] ),
    .A1(\core_pipeline.decode_to_execute_rs1_bypass[16] ),
    .S(net488),
    .X(_03804_));
 sky130_fd_sc_hd__inv_2 _07258_ (.A(_03804_),
    .Y(_03805_));
 sky130_fd_sc_hd__a22o_1 _07259_ (.A1(_03800_),
    .A2(_03802_),
    .B1(_03803_),
    .B2(_03805_),
    .X(_03806_));
 sky130_fd_sc_hd__nor2_1 _07260_ (.A(_03793_),
    .B(_03795_),
    .Y(_03807_));
 sky130_fd_sc_hd__nor2_1 _07261_ (.A(_03800_),
    .B(_03802_),
    .Y(_03808_));
 sky130_fd_sc_hd__nor2_1 _07262_ (.A(_03807_),
    .B(_03808_),
    .Y(_03809_));
 sky130_fd_sc_hd__a21o_1 _07263_ (.A1(_03806_),
    .A2(_03809_),
    .B1(_03799_),
    .X(_03810_));
 sky130_fd_sc_hd__or2_1 _07264_ (.A(_03796_),
    .B(_03798_),
    .X(_03811_));
 sky130_fd_sc_hd__or2_1 _07265_ (.A(_03786_),
    .B(_03788_),
    .X(_03812_));
 sky130_fd_sc_hd__a31o_1 _07266_ (.A1(_03810_),
    .A2(_03811_),
    .A3(_03812_),
    .B1(_03792_),
    .X(_03813_));
 sky130_fd_sc_hd__o2bb2a_1 _07267_ (.A1_N(_03784_),
    .A2_N(_03785_),
    .B1(_03789_),
    .B2(_03791_),
    .X(_03814_));
 sky130_fd_sc_hd__nand2_1 _07268_ (.A(_03813_),
    .B(_03814_),
    .Y(_03815_));
 sky130_fd_sc_hd__o221a_1 _07269_ (.A1(_03780_),
    .A2(_03781_),
    .B1(_03784_),
    .B2(_03785_),
    .C1(_03815_),
    .X(_03816_));
 sky130_fd_sc_hd__or3_1 _07270_ (.A(_03806_),
    .B(_03807_),
    .C(_03808_),
    .X(_03817_));
 sky130_fd_sc_hd__o21a_1 _07271_ (.A1(_03803_),
    .A2(_03805_),
    .B1(_03811_),
    .X(_03818_));
 sky130_fd_sc_hd__o221a_1 _07272_ (.A1(_03780_),
    .A2(_03781_),
    .B1(_03784_),
    .B2(_03785_),
    .C1(_03814_),
    .X(_03819_));
 sky130_fd_sc_hd__and4b_1 _07273_ (.A_N(_03782_),
    .B(_03812_),
    .C(_03818_),
    .D(_03819_),
    .X(_03820_));
 sky130_fd_sc_hd__or4b_2 _07274_ (.A(_03792_),
    .B(_03799_),
    .C(_03817_),
    .D_N(_03820_),
    .X(_03821_));
 sky130_fd_sc_hd__mux2_4 _07275_ (.A0(\core_pipeline.decode_to_execute_rs2_data[15] ),
    .A1(\core_pipeline.decode_to_execute_rs2_bypass[15] ),
    .S(net486),
    .X(_03822_));
 sky130_fd_sc_hd__inv_2 _07276_ (.A(_03822_),
    .Y(_03823_));
 sky130_fd_sc_hd__mux2_4 _07277_ (.A0(\core_pipeline.decode_to_execute_rs1_data[15] ),
    .A1(\core_pipeline.decode_to_execute_rs1_bypass[15] ),
    .S(net488),
    .X(_03824_));
 sky130_fd_sc_hd__and2_1 _07278_ (.A(_03823_),
    .B(_03824_),
    .X(_03825_));
 sky130_fd_sc_hd__mux2_8 _07279_ (.A0(\core_pipeline.decode_to_execute_rs2_data[14] ),
    .A1(\core_pipeline.decode_to_execute_rs2_bypass[14] ),
    .S(net486),
    .X(_03826_));
 sky130_fd_sc_hd__inv_2 _07280_ (.A(_03826_),
    .Y(_03827_));
 sky130_fd_sc_hd__mux2_8 _07281_ (.A0(\core_pipeline.decode_to_execute_rs1_data[14] ),
    .A1(\core_pipeline.decode_to_execute_rs1_bypass[14] ),
    .S(net488),
    .X(_03828_));
 sky130_fd_sc_hd__o22a_1 _07282_ (.A1(_03823_),
    .A2(_03824_),
    .B1(_03827_),
    .B2(_03828_),
    .X(_03829_));
 sky130_fd_sc_hd__mux2_8 _07283_ (.A0(\core_pipeline.decode_to_execute_rs2_data[13] ),
    .A1(\core_pipeline.decode_to_execute_rs2_bypass[13] ),
    .S(net486),
    .X(_03830_));
 sky130_fd_sc_hd__inv_2 _07284_ (.A(_03830_),
    .Y(_03831_));
 sky130_fd_sc_hd__mux2_4 _07285_ (.A0(\core_pipeline.decode_to_execute_rs1_data[13] ),
    .A1(\core_pipeline.decode_to_execute_rs1_bypass[13] ),
    .S(net488),
    .X(_03832_));
 sky130_fd_sc_hd__a22o_1 _07286_ (.A1(_03827_),
    .A2(_03828_),
    .B1(_03831_),
    .B2(_03832_),
    .X(_03833_));
 sky130_fd_sc_hd__or2_1 _07287_ (.A(_03831_),
    .B(_03832_),
    .X(_03834_));
 sky130_fd_sc_hd__nand2b_2 _07288_ (.A_N(\core_pipeline.decode_to_execute_rs2_bypass[12] ),
    .B(net486),
    .Y(_03835_));
 sky130_fd_sc_hd__o21a_4 _07289_ (.A1(net486),
    .A2(\core_pipeline.decode_to_execute_rs2_data[12] ),
    .B1(_03835_),
    .X(_03836_));
 sky130_fd_sc_hd__o21ai_4 _07290_ (.A1(net486),
    .A2(\core_pipeline.decode_to_execute_rs2_data[12] ),
    .B1(_03835_),
    .Y(_03837_));
 sky130_fd_sc_hd__mux2_8 _07291_ (.A0(\core_pipeline.decode_to_execute_rs1_data[12] ),
    .A1(\core_pipeline.decode_to_execute_rs1_bypass[12] ),
    .S(net488),
    .X(_03838_));
 sky130_fd_sc_hd__nor2_1 _07292_ (.A(_03837_),
    .B(_03838_),
    .Y(_03839_));
 sky130_fd_sc_hd__mux2_8 _07293_ (.A0(\core_pipeline.decode_to_execute_rs2_data[10] ),
    .A1(\core_pipeline.decode_to_execute_rs2_bypass[10] ),
    .S(net486),
    .X(_03840_));
 sky130_fd_sc_hd__inv_2 _07294_ (.A(_03840_),
    .Y(_03841_));
 sky130_fd_sc_hd__mux2_4 _07295_ (.A0(\core_pipeline.decode_to_execute_rs1_data[10] ),
    .A1(\core_pipeline.decode_to_execute_rs1_bypass[10] ),
    .S(net488),
    .X(_03842_));
 sky130_fd_sc_hd__mux2_8 _07296_ (.A0(\core_pipeline.decode_to_execute_rs2_data[11] ),
    .A1(\core_pipeline.decode_to_execute_rs2_bypass[11] ),
    .S(net486),
    .X(_03843_));
 sky130_fd_sc_hd__inv_2 _07297_ (.A(_03843_),
    .Y(_03844_));
 sky130_fd_sc_hd__mux2_8 _07298_ (.A0(\core_pipeline.decode_to_execute_rs1_data[11] ),
    .A1(\core_pipeline.decode_to_execute_rs1_bypass[11] ),
    .S(net488),
    .X(_03845_));
 sky130_fd_sc_hd__o22a_1 _07299_ (.A1(_03841_),
    .A2(_03842_),
    .B1(_03844_),
    .B2(_03845_),
    .X(_03846_));
 sky130_fd_sc_hd__mux2_8 _07300_ (.A0(\core_pipeline.decode_to_execute_rs2_data[9] ),
    .A1(\core_pipeline.decode_to_execute_rs2_bypass[9] ),
    .S(net486),
    .X(_03847_));
 sky130_fd_sc_hd__inv_2 _07301_ (.A(_03847_),
    .Y(_03848_));
 sky130_fd_sc_hd__mux2_8 _07302_ (.A0(\core_pipeline.decode_to_execute_rs1_data[9] ),
    .A1(\core_pipeline.decode_to_execute_rs1_bypass[9] ),
    .S(net488),
    .X(_03849_));
 sky130_fd_sc_hd__a22o_1 _07303_ (.A1(_03841_),
    .A2(_03842_),
    .B1(_03848_),
    .B2(_03849_),
    .X(_03850_));
 sky130_fd_sc_hd__a22o_1 _07304_ (.A1(_03837_),
    .A2(_03838_),
    .B1(_03844_),
    .B2(_03845_),
    .X(_03851_));
 sky130_fd_sc_hd__mux2_8 _07305_ (.A0(\core_pipeline.decode_to_execute_rs2_data[8] ),
    .A1(\core_pipeline.decode_to_execute_rs2_bypass[8] ),
    .S(net487),
    .X(_03852_));
 sky130_fd_sc_hd__inv_2 _07306_ (.A(_03852_),
    .Y(_03853_));
 sky130_fd_sc_hd__mux2_8 _07307_ (.A0(\core_pipeline.decode_to_execute_rs1_data[8] ),
    .A1(\core_pipeline.decode_to_execute_rs1_bypass[8] ),
    .S(net488),
    .X(_03854_));
 sky130_fd_sc_hd__o22a_1 _07308_ (.A1(_03848_),
    .A2(_03849_),
    .B1(_03853_),
    .B2(_03854_),
    .X(_03855_));
 sky130_fd_sc_hd__o21a_1 _07309_ (.A1(_03850_),
    .A2(_03855_),
    .B1(_03846_),
    .X(_03856_));
 sky130_fd_sc_hd__o221a_1 _07310_ (.A1(_03837_),
    .A2(_03838_),
    .B1(_03851_),
    .B2(_03856_),
    .C1(_03834_),
    .X(_03857_));
 sky130_fd_sc_hd__o21a_1 _07311_ (.A1(_03833_),
    .A2(_03857_),
    .B1(_03829_),
    .X(_03858_));
 sky130_fd_sc_hd__mux2_8 _07312_ (.A0(\core_pipeline.decode_to_execute_rs2_data[6] ),
    .A1(\core_pipeline.decode_to_execute_rs2_bypass[6] ),
    .S(net487),
    .X(_03859_));
 sky130_fd_sc_hd__mux2_8 _07313_ (.A0(\core_pipeline.decode_to_execute_rs1_data[6] ),
    .A1(\core_pipeline.decode_to_execute_rs1_bypass[6] ),
    .S(net489),
    .X(_03860_));
 sky130_fd_sc_hd__inv_2 _07314_ (.A(_03860_),
    .Y(_03861_));
 sky130_fd_sc_hd__mux2_8 _07315_ (.A0(\core_pipeline.decode_to_execute_rs2_data[7] ),
    .A1(\core_pipeline.decode_to_execute_rs2_bypass[7] ),
    .S(net486),
    .X(_03862_));
 sky130_fd_sc_hd__mux2_4 _07316_ (.A0(\core_pipeline.decode_to_execute_rs1_data[7] ),
    .A1(\core_pipeline.decode_to_execute_rs1_bypass[7] ),
    .S(net488),
    .X(_03863_));
 sky130_fd_sc_hd__inv_2 _07317_ (.A(_03863_),
    .Y(_03864_));
 sky130_fd_sc_hd__a22o_1 _07318_ (.A1(_03859_),
    .A2(_03861_),
    .B1(_03862_),
    .B2(_03864_),
    .X(_03865_));
 sky130_fd_sc_hd__mux2_8 _07319_ (.A0(\core_pipeline.decode_to_execute_rs2_data[5] ),
    .A1(\core_pipeline.decode_to_execute_rs2_bypass[5] ),
    .S(net487),
    .X(_03866_));
 sky130_fd_sc_hd__mux2_4 _07320_ (.A0(\core_pipeline.decode_to_execute_rs1_data[5] ),
    .A1(\core_pipeline.decode_to_execute_rs1_bypass[5] ),
    .S(net489),
    .X(_03867_));
 sky130_fd_sc_hd__inv_2 _07321_ (.A(_03867_),
    .Y(_03868_));
 sky130_fd_sc_hd__mux2_8 _07322_ (.A0(\core_pipeline.decode_to_execute_rs2_data[4] ),
    .A1(\core_pipeline.decode_to_execute_rs2_bypass[4] ),
    .S(net486),
    .X(_03869_));
 sky130_fd_sc_hd__mux2_4 _07323_ (.A0(\core_pipeline.decode_to_execute_rs1_data[4] ),
    .A1(\core_pipeline.decode_to_execute_rs1_bypass[4] ),
    .S(net488),
    .X(_03870_));
 sky130_fd_sc_hd__inv_2 _07324_ (.A(_03870_),
    .Y(_03871_));
 sky130_fd_sc_hd__a22o_1 _07325_ (.A1(_03866_),
    .A2(_03868_),
    .B1(_03869_),
    .B2(_03871_),
    .X(_03872_));
 sky130_fd_sc_hd__mux2_8 _07326_ (.A0(\core_pipeline.decode_to_execute_rs2_data[1] ),
    .A1(\core_pipeline.decode_to_execute_rs2_bypass[1] ),
    .S(net487),
    .X(_03873_));
 sky130_fd_sc_hd__inv_2 _07327_ (.A(_03873_),
    .Y(_03874_));
 sky130_fd_sc_hd__mux2_4 _07328_ (.A0(\core_pipeline.decode_to_execute_rs1_data[1] ),
    .A1(\core_pipeline.decode_to_execute_rs1_bypass[1] ),
    .S(net489),
    .X(_03875_));
 sky130_fd_sc_hd__inv_2 _07329_ (.A(_03875_),
    .Y(_03876_));
 sky130_fd_sc_hd__mux2_4 _07330_ (.A0(\core_pipeline.decode_to_execute_rs2_data[0] ),
    .A1(\core_pipeline.decode_to_execute_rs2_bypass[0] ),
    .S(net486),
    .X(_03877_));
 sky130_fd_sc_hd__inv_2 _07331_ (.A(_03877_),
    .Y(_03878_));
 sky130_fd_sc_hd__mux2_2 _07332_ (.A0(\core_pipeline.decode_to_execute_rs1_data[0] ),
    .A1(\core_pipeline.decode_to_execute_rs1_bypass[0] ),
    .S(net488),
    .X(_03879_));
 sky130_fd_sc_hd__o2bb2a_1 _07333_ (.A1_N(_03878_),
    .A2_N(_03879_),
    .B1(_03873_),
    .B2(_03876_),
    .X(_03880_));
 sky130_fd_sc_hd__mux2_8 _07334_ (.A0(\core_pipeline.decode_to_execute_rs2_data[2] ),
    .A1(\core_pipeline.decode_to_execute_rs2_bypass[2] ),
    .S(net487),
    .X(_03881_));
 sky130_fd_sc_hd__mux2_8 _07335_ (.A0(\core_pipeline.decode_to_execute_rs1_data[2] ),
    .A1(\core_pipeline.decode_to_execute_rs1_bypass[2] ),
    .S(net489),
    .X(_03882_));
 sky130_fd_sc_hd__inv_2 _07336_ (.A(_03882_),
    .Y(_03883_));
 sky130_fd_sc_hd__or2_1 _07337_ (.A(_03881_),
    .B(_03883_),
    .X(_03884_));
 sky130_fd_sc_hd__o211a_1 _07338_ (.A1(_03874_),
    .A2(_03875_),
    .B1(_03880_),
    .C1(_03884_),
    .X(_03885_));
 sky130_fd_sc_hd__mux2_8 _07339_ (.A0(\core_pipeline.decode_to_execute_rs2_data[3] ),
    .A1(\core_pipeline.decode_to_execute_rs2_bypass[3] ),
    .S(net486),
    .X(_03886_));
 sky130_fd_sc_hd__mux2_4 _07340_ (.A0(\core_pipeline.decode_to_execute_rs1_data[3] ),
    .A1(\core_pipeline.decode_to_execute_rs1_bypass[3] ),
    .S(net488),
    .X(_03887_));
 sky130_fd_sc_hd__inv_2 _07341_ (.A(_03887_),
    .Y(_03888_));
 sky130_fd_sc_hd__a22o_1 _07342_ (.A1(_03881_),
    .A2(_03883_),
    .B1(_03886_),
    .B2(_03888_),
    .X(_03889_));
 sky130_fd_sc_hd__a311o_1 _07343_ (.A1(_03873_),
    .A2(_03876_),
    .A3(_03884_),
    .B1(_03885_),
    .C1(_03889_),
    .X(_03890_));
 sky130_fd_sc_hd__o22a_1 _07344_ (.A1(_03869_),
    .A2(_03871_),
    .B1(_03886_),
    .B2(_03888_),
    .X(_03891_));
 sky130_fd_sc_hd__a21oi_1 _07345_ (.A1(_03890_),
    .A2(_03891_),
    .B1(_03872_),
    .Y(_03892_));
 sky130_fd_sc_hd__o22ai_2 _07346_ (.A1(_03859_),
    .A2(_03861_),
    .B1(_03866_),
    .B2(_03868_),
    .Y(_03893_));
 sky130_fd_sc_hd__o21ba_1 _07347_ (.A1(_03892_),
    .A2(_03893_),
    .B1_N(_03865_),
    .X(_03894_));
 sky130_fd_sc_hd__or3b_1 _07348_ (.A(_03839_),
    .B(_03833_),
    .C_N(_03834_),
    .X(_03895_));
 sky130_fd_sc_hd__a21oi_1 _07349_ (.A1(_03853_),
    .A2(_03854_),
    .B1(_03825_),
    .Y(_03896_));
 sky130_fd_sc_hd__and4_1 _07350_ (.A(_03829_),
    .B(_03846_),
    .C(_03855_),
    .D(_03896_),
    .X(_03897_));
 sky130_fd_sc_hd__or4b_2 _07351_ (.A(_03850_),
    .B(_03851_),
    .C(_03895_),
    .D_N(_03897_),
    .X(_03898_));
 sky130_fd_sc_hd__nor2_1 _07352_ (.A(_03862_),
    .B(_03864_),
    .Y(_03899_));
 sky130_fd_sc_hd__o32a_1 _07353_ (.A1(_03894_),
    .A2(_03898_),
    .A3(_03899_),
    .B1(_03858_),
    .B2(_03825_),
    .X(_03900_));
 sky130_fd_sc_hd__o22a_1 _07354_ (.A1(_03782_),
    .A2(_03816_),
    .B1(_03821_),
    .B2(_03900_),
    .X(_03901_));
 sky130_fd_sc_hd__or2_1 _07355_ (.A(_03778_),
    .B(_03901_),
    .X(_03902_));
 sky130_fd_sc_hd__nand2_1 _07356_ (.A(_03759_),
    .B(_03764_),
    .Y(_03903_));
 sky130_fd_sc_hd__a31o_1 _07357_ (.A1(_03763_),
    .A2(_03769_),
    .A3(_03903_),
    .B1(_03752_),
    .X(_03904_));
 sky130_fd_sc_hd__a21oi_1 _07358_ (.A1(_03775_),
    .A2(_03904_),
    .B1(_03774_),
    .Y(_03905_));
 sky130_fd_sc_hd__o221a_1 _07359_ (.A1(_03742_),
    .A2(_03743_),
    .B1(_03773_),
    .B2(_03905_),
    .C1(\core_pipeline.decode_to_execute_cmp_function[2] ),
    .X(_03906_));
 sky130_fd_sc_hd__or4_1 _07360_ (.A(_03865_),
    .B(_03872_),
    .C(_03889_),
    .D(_03893_),
    .X(_03907_));
 sky130_fd_sc_hd__o221a_1 _07361_ (.A1(_03862_),
    .A2(_03864_),
    .B1(_03878_),
    .B2(_03879_),
    .C1(_03891_),
    .X(_03908_));
 sky130_fd_sc_hd__nand2_1 _07362_ (.A(_03885_),
    .B(_03908_),
    .Y(_03909_));
 sky130_fd_sc_hd__or4_1 _07363_ (.A(_03821_),
    .B(_03898_),
    .C(_03907_),
    .D(_03909_),
    .X(_03910_));
 sky130_fd_sc_hd__a2bb2o_1 _07364_ (.A1_N(_03778_),
    .A2_N(_03910_),
    .B1(_03906_),
    .B2(_03902_),
    .X(_03911_));
 sky130_fd_sc_hd__xnor2_1 _07365_ (.A(_03745_),
    .B(_03911_),
    .Y(_00039_));
 sky130_fd_sc_hd__nand2_8 _07366_ (.A(\core_pipeline.memory_to_writeback_rd_address[4] ),
    .B(_03480_),
    .Y(_03912_));
 sky130_fd_sc_hd__nand2_8 _07367_ (.A(\core_pipeline.memory_to_writeback_rd_address[0] ),
    .B(_03480_),
    .Y(_03913_));
 sky130_fd_sc_hd__nand2_4 _07368_ (.A(\core_pipeline.memory_to_writeback_rd_address[1] ),
    .B(_03480_),
    .Y(_03914_));
 sky130_fd_sc_hd__nand3_4 _07369_ (.A(\core_pipeline.memory_to_writeback_rd_address[0] ),
    .B(\core_pipeline.memory_to_writeback_rd_address[1] ),
    .C(_03480_),
    .Y(_03915_));
 sky130_fd_sc_hd__or4_4 _07370_ (.A(\core_pipeline.memory_to_writeback_rd_address[2] ),
    .B(\core_pipeline.memory_to_writeback_rd_address[3] ),
    .C(_03912_),
    .D(_03915_),
    .X(_03916_));
 sky130_fd_sc_hd__and3_1 _07371_ (.A(\core_pipeline.memory_to_writeback_next_pc[0] ),
    .B(net508),
    .C(net510),
    .X(_03917_));
 sky130_fd_sc_hd__and2b_2 _07372_ (.A_N(net509),
    .B(net506),
    .X(_03918_));
 sky130_fd_sc_hd__or2_2 _07373_ (.A(net508),
    .B(net510),
    .X(_03919_));
 sky130_fd_sc_hd__and2b_1 _07374_ (.A_N(net506),
    .B(net510),
    .X(_03920_));
 sky130_fd_sc_hd__a221o_1 _07375_ (.A1(\core_pipeline.memory_to_writeback_load_data[0] ),
    .A2(net444),
    .B1(net440),
    .B2(\core_pipeline.memory_to_writeback_csr_data[0] ),
    .C1(_03917_),
    .X(_03921_));
 sky130_fd_sc_hd__mux2_8 _07376_ (.A0(\core_pipeline.memory_to_writeback_alu_data[0] ),
    .A1(_03921_),
    .S(net442),
    .X(_03922_));
 sky130_fd_sc_hd__mux2_1 _07377_ (.A0(net348),
    .A1(\core_pipeline.pipeline_registers.registers[19][0] ),
    .S(net259),
    .X(_00041_));
 sky130_fd_sc_hd__and3_1 _07378_ (.A(\core_pipeline.memory_to_writeback_next_pc[1] ),
    .B(net508),
    .C(net510),
    .X(_03923_));
 sky130_fd_sc_hd__a221o_1 _07379_ (.A1(\core_pipeline.memory_to_writeback_load_data[1] ),
    .A2(net444),
    .B1(net440),
    .B2(\core_pipeline.memory_to_writeback_csr_data[1] ),
    .C1(_03923_),
    .X(_03924_));
 sky130_fd_sc_hd__mux2_8 _07380_ (.A0(\core_pipeline.memory_to_writeback_alu_data[1] ),
    .A1(_03924_),
    .S(net442),
    .X(_03925_));
 sky130_fd_sc_hd__mux2_1 _07381_ (.A0(net346),
    .A1(\core_pipeline.pipeline_registers.registers[19][1] ),
    .S(net260),
    .X(_00042_));
 sky130_fd_sc_hd__and3_1 _07382_ (.A(\core_pipeline.memory_to_writeback_next_pc[2] ),
    .B(net508),
    .C(net510),
    .X(_03926_));
 sky130_fd_sc_hd__a221o_1 _07383_ (.A1(\core_pipeline.memory_to_writeback_load_data[2] ),
    .A2(net444),
    .B1(net440),
    .B2(\core_pipeline.memory_to_writeback_csr_data[2] ),
    .C1(_03926_),
    .X(_03927_));
 sky130_fd_sc_hd__mux2_8 _07384_ (.A0(\core_pipeline.memory_to_writeback_alu_data[2] ),
    .A1(_03927_),
    .S(net442),
    .X(_03928_));
 sky130_fd_sc_hd__mux2_1 _07385_ (.A0(net344),
    .A1(\core_pipeline.pipeline_registers.registers[19][2] ),
    .S(net260),
    .X(_00043_));
 sky130_fd_sc_hd__and3_1 _07386_ (.A(\core_pipeline.memory_to_writeback_next_pc[3] ),
    .B(net508),
    .C(net510),
    .X(_03929_));
 sky130_fd_sc_hd__a221o_1 _07387_ (.A1(\core_pipeline.memory_to_writeback_load_data[3] ),
    .A2(net444),
    .B1(net440),
    .B2(\core_pipeline.memory_to_writeback_csr_data[3] ),
    .C1(_03929_),
    .X(_03930_));
 sky130_fd_sc_hd__mux2_8 _07388_ (.A0(\core_pipeline.memory_to_writeback_alu_data[3] ),
    .A1(_03930_),
    .S(net442),
    .X(_03931_));
 sky130_fd_sc_hd__mux2_1 _07389_ (.A0(net342),
    .A1(\core_pipeline.pipeline_registers.registers[19][3] ),
    .S(net259),
    .X(_00044_));
 sky130_fd_sc_hd__and3_1 _07390_ (.A(\core_pipeline.memory_to_writeback_next_pc[4] ),
    .B(net508),
    .C(net510),
    .X(_03932_));
 sky130_fd_sc_hd__a221o_1 _07391_ (.A1(\core_pipeline.memory_to_writeback_load_data[4] ),
    .A2(net444),
    .B1(net440),
    .B2(\core_pipeline.memory_to_writeback_csr_data[4] ),
    .C1(_03932_),
    .X(_03933_));
 sky130_fd_sc_hd__mux2_8 _07392_ (.A0(\core_pipeline.memory_to_writeback_alu_data[4] ),
    .A1(_03933_),
    .S(net442),
    .X(_03934_));
 sky130_fd_sc_hd__mux2_1 _07393_ (.A0(net340),
    .A1(\core_pipeline.pipeline_registers.registers[19][4] ),
    .S(net259),
    .X(_00045_));
 sky130_fd_sc_hd__and3_1 _07394_ (.A(\core_pipeline.memory_to_writeback_next_pc[5] ),
    .B(net508),
    .C(net510),
    .X(_03935_));
 sky130_fd_sc_hd__a221o_1 _07395_ (.A1(\core_pipeline.memory_to_writeback_load_data[5] ),
    .A2(net444),
    .B1(net440),
    .B2(\core_pipeline.memory_to_writeback_csr_data[5] ),
    .C1(_03935_),
    .X(_03936_));
 sky130_fd_sc_hd__mux2_2 _07396_ (.A0(\core_pipeline.memory_to_writeback_alu_data[5] ),
    .A1(_03936_),
    .S(net442),
    .X(_03937_));
 sky130_fd_sc_hd__mux2_1 _07397_ (.A0(net339),
    .A1(\core_pipeline.pipeline_registers.registers[19][5] ),
    .S(net260),
    .X(_00046_));
 sky130_fd_sc_hd__and3_1 _07398_ (.A(\core_pipeline.memory_to_writeback_next_pc[6] ),
    .B(net508),
    .C(net510),
    .X(_03938_));
 sky130_fd_sc_hd__a221o_1 _07399_ (.A1(\core_pipeline.memory_to_writeback_load_data[6] ),
    .A2(net444),
    .B1(net440),
    .B2(\core_pipeline.memory_to_writeback_csr_data[6] ),
    .C1(_03938_),
    .X(_03939_));
 sky130_fd_sc_hd__mux2_8 _07400_ (.A0(\core_pipeline.memory_to_writeback_alu_data[6] ),
    .A1(_03939_),
    .S(net442),
    .X(_03940_));
 sky130_fd_sc_hd__mux2_1 _07401_ (.A0(net336),
    .A1(\core_pipeline.pipeline_registers.registers[19][6] ),
    .S(net260),
    .X(_00047_));
 sky130_fd_sc_hd__and3_1 _07402_ (.A(\core_pipeline.memory_to_writeback_next_pc[7] ),
    .B(net508),
    .C(net510),
    .X(_03941_));
 sky130_fd_sc_hd__a221o_1 _07403_ (.A1(\core_pipeline.memory_to_writeback_load_data[7] ),
    .A2(net444),
    .B1(net440),
    .B2(\core_pipeline.memory_to_writeback_csr_data[7] ),
    .C1(_03941_),
    .X(_03942_));
 sky130_fd_sc_hd__mux2_4 _07404_ (.A0(\core_pipeline.memory_to_writeback_alu_data[7] ),
    .A1(_03942_),
    .S(net442),
    .X(_03943_));
 sky130_fd_sc_hd__mux2_1 _07405_ (.A0(net333),
    .A1(\core_pipeline.pipeline_registers.registers[19][7] ),
    .S(net259),
    .X(_00048_));
 sky130_fd_sc_hd__and3_1 _07406_ (.A(\core_pipeline.memory_to_writeback_next_pc[8] ),
    .B(net507),
    .C(net509),
    .X(_03944_));
 sky130_fd_sc_hd__a221o_1 _07407_ (.A1(\core_pipeline.memory_to_writeback_load_data[8] ),
    .A2(net443),
    .B1(net439),
    .B2(\core_pipeline.memory_to_writeback_csr_data[8] ),
    .C1(_03944_),
    .X(_03945_));
 sky130_fd_sc_hd__mux2_8 _07408_ (.A0(\core_pipeline.memory_to_writeback_alu_data[8] ),
    .A1(_03945_),
    .S(net441),
    .X(_03946_));
 sky130_fd_sc_hd__mux2_1 _07409_ (.A0(net331),
    .A1(\core_pipeline.pipeline_registers.registers[19][8] ),
    .S(net259),
    .X(_00049_));
 sky130_fd_sc_hd__and3_1 _07410_ (.A(\core_pipeline.memory_to_writeback_next_pc[9] ),
    .B(net506),
    .C(net509),
    .X(_03947_));
 sky130_fd_sc_hd__a221o_1 _07411_ (.A1(\core_pipeline.memory_to_writeback_load_data[9] ),
    .A2(net443),
    .B1(net439),
    .B2(\core_pipeline.memory_to_writeback_csr_data[9] ),
    .C1(_03947_),
    .X(_03948_));
 sky130_fd_sc_hd__mux2_8 _07412_ (.A0(\core_pipeline.memory_to_writeback_alu_data[9] ),
    .A1(_03948_),
    .S(net441),
    .X(_03949_));
 sky130_fd_sc_hd__mux2_1 _07413_ (.A0(net330),
    .A1(\core_pipeline.pipeline_registers.registers[19][9] ),
    .S(net259),
    .X(_00050_));
 sky130_fd_sc_hd__and3_1 _07414_ (.A(\core_pipeline.memory_to_writeback_next_pc[10] ),
    .B(net506),
    .C(net509),
    .X(_03950_));
 sky130_fd_sc_hd__a221o_1 _07415_ (.A1(\core_pipeline.memory_to_writeback_load_data[10] ),
    .A2(net443),
    .B1(net439),
    .B2(\core_pipeline.memory_to_writeback_csr_data[10] ),
    .C1(_03950_),
    .X(_03951_));
 sky130_fd_sc_hd__mux2_8 _07416_ (.A0(\core_pipeline.memory_to_writeback_alu_data[10] ),
    .A1(_03951_),
    .S(net441),
    .X(_03952_));
 sky130_fd_sc_hd__mux2_1 _07417_ (.A0(net327),
    .A1(\core_pipeline.pipeline_registers.registers[19][10] ),
    .S(net259),
    .X(_00051_));
 sky130_fd_sc_hd__and3_1 _07418_ (.A(\core_pipeline.memory_to_writeback_next_pc[11] ),
    .B(net506),
    .C(net509),
    .X(_03953_));
 sky130_fd_sc_hd__a221o_1 _07419_ (.A1(\core_pipeline.memory_to_writeback_load_data[11] ),
    .A2(net444),
    .B1(net440),
    .B2(\core_pipeline.memory_to_writeback_csr_data[11] ),
    .C1(_03953_),
    .X(_03954_));
 sky130_fd_sc_hd__mux2_8 _07420_ (.A0(\core_pipeline.memory_to_writeback_alu_data[11] ),
    .A1(_03954_),
    .S(net442),
    .X(_03955_));
 sky130_fd_sc_hd__mux2_1 _07421_ (.A0(net325),
    .A1(\core_pipeline.pipeline_registers.registers[19][11] ),
    .S(net259),
    .X(_00052_));
 sky130_fd_sc_hd__and3_1 _07422_ (.A(\core_pipeline.memory_to_writeback_next_pc[12] ),
    .B(net506),
    .C(net509),
    .X(_03956_));
 sky130_fd_sc_hd__a221o_1 _07423_ (.A1(\core_pipeline.memory_to_writeback_load_data[12] ),
    .A2(net443),
    .B1(net439),
    .B2(\core_pipeline.memory_to_writeback_csr_data[12] ),
    .C1(_03956_),
    .X(_03957_));
 sky130_fd_sc_hd__mux2_8 _07424_ (.A0(\core_pipeline.memory_to_writeback_alu_data[12] ),
    .A1(_03957_),
    .S(net441),
    .X(_03958_));
 sky130_fd_sc_hd__mux2_1 _07425_ (.A0(net323),
    .A1(\core_pipeline.pipeline_registers.registers[19][12] ),
    .S(net259),
    .X(_00053_));
 sky130_fd_sc_hd__and3_1 _07426_ (.A(\core_pipeline.memory_to_writeback_next_pc[13] ),
    .B(net506),
    .C(net509),
    .X(_03959_));
 sky130_fd_sc_hd__a221o_1 _07427_ (.A1(\core_pipeline.memory_to_writeback_load_data[13] ),
    .A2(net443),
    .B1(net439),
    .B2(\core_pipeline.memory_to_writeback_csr_data[13] ),
    .C1(_03959_),
    .X(_03960_));
 sky130_fd_sc_hd__mux2_8 _07428_ (.A0(\core_pipeline.memory_to_writeback_alu_data[13] ),
    .A1(_03960_),
    .S(net441),
    .X(_03961_));
 sky130_fd_sc_hd__mux2_1 _07429_ (.A0(net321),
    .A1(\core_pipeline.pipeline_registers.registers[19][13] ),
    .S(net259),
    .X(_00054_));
 sky130_fd_sc_hd__and3_1 _07430_ (.A(\core_pipeline.memory_to_writeback_next_pc[14] ),
    .B(net506),
    .C(net509),
    .X(_03962_));
 sky130_fd_sc_hd__a221o_1 _07431_ (.A1(\core_pipeline.memory_to_writeback_load_data[14] ),
    .A2(net443),
    .B1(net439),
    .B2(\core_pipeline.memory_to_writeback_csr_data[14] ),
    .C1(_03962_),
    .X(_03963_));
 sky130_fd_sc_hd__mux2_8 _07432_ (.A0(\core_pipeline.memory_to_writeback_alu_data[14] ),
    .A1(_03963_),
    .S(net441),
    .X(_03964_));
 sky130_fd_sc_hd__mux2_1 _07433_ (.A0(net319),
    .A1(\core_pipeline.pipeline_registers.registers[19][14] ),
    .S(net259),
    .X(_00055_));
 sky130_fd_sc_hd__and3_1 _07434_ (.A(\core_pipeline.memory_to_writeback_next_pc[15] ),
    .B(net506),
    .C(net509),
    .X(_03965_));
 sky130_fd_sc_hd__a221o_1 _07435_ (.A1(\core_pipeline.memory_to_writeback_load_data[15] ),
    .A2(net443),
    .B1(net439),
    .B2(\core_pipeline.memory_to_writeback_csr_data[15] ),
    .C1(_03965_),
    .X(_03966_));
 sky130_fd_sc_hd__mux2_8 _07436_ (.A0(\core_pipeline.memory_to_writeback_alu_data[15] ),
    .A1(_03966_),
    .S(net441),
    .X(_03967_));
 sky130_fd_sc_hd__mux2_1 _07437_ (.A0(net317),
    .A1(\core_pipeline.pipeline_registers.registers[19][15] ),
    .S(net259),
    .X(_00056_));
 sky130_fd_sc_hd__and3_1 _07438_ (.A(\core_pipeline.memory_to_writeback_next_pc[16] ),
    .B(net506),
    .C(net509),
    .X(_03968_));
 sky130_fd_sc_hd__a221o_1 _07439_ (.A1(\core_pipeline.memory_to_writeback_load_data[16] ),
    .A2(net443),
    .B1(net439),
    .B2(\core_pipeline.memory_to_writeback_csr_data[16] ),
    .C1(_03968_),
    .X(_03969_));
 sky130_fd_sc_hd__mux2_8 _07440_ (.A0(\core_pipeline.memory_to_writeback_alu_data[16] ),
    .A1(_03969_),
    .S(net441),
    .X(_03970_));
 sky130_fd_sc_hd__mux2_1 _07441_ (.A0(net316),
    .A1(\core_pipeline.pipeline_registers.registers[19][16] ),
    .S(net259),
    .X(_00057_));
 sky130_fd_sc_hd__and3_1 _07442_ (.A(\core_pipeline.memory_to_writeback_next_pc[17] ),
    .B(net506),
    .C(net509),
    .X(_03971_));
 sky130_fd_sc_hd__a221o_1 _07443_ (.A1(\core_pipeline.memory_to_writeback_load_data[17] ),
    .A2(net443),
    .B1(net439),
    .B2(\core_pipeline.memory_to_writeback_csr_data[17] ),
    .C1(_03971_),
    .X(_03972_));
 sky130_fd_sc_hd__mux2_8 _07444_ (.A0(\core_pipeline.memory_to_writeback_alu_data[17] ),
    .A1(_03972_),
    .S(net441),
    .X(_03973_));
 sky130_fd_sc_hd__mux2_1 _07445_ (.A0(net313),
    .A1(\core_pipeline.pipeline_registers.registers[19][17] ),
    .S(net260),
    .X(_00058_));
 sky130_fd_sc_hd__and3_1 _07446_ (.A(\core_pipeline.memory_to_writeback_next_pc[18] ),
    .B(net506),
    .C(net510),
    .X(_03974_));
 sky130_fd_sc_hd__a221o_1 _07447_ (.A1(\core_pipeline.memory_to_writeback_load_data[18] ),
    .A2(net443),
    .B1(net439),
    .B2(\core_pipeline.memory_to_writeback_csr_data[18] ),
    .C1(_03974_),
    .X(_03975_));
 sky130_fd_sc_hd__mux2_8 _07448_ (.A0(\core_pipeline.memory_to_writeback_alu_data[18] ),
    .A1(_03975_),
    .S(net441),
    .X(_03976_));
 sky130_fd_sc_hd__mux2_1 _07449_ (.A0(net310),
    .A1(\core_pipeline.pipeline_registers.registers[19][18] ),
    .S(net260),
    .X(_00059_));
 sky130_fd_sc_hd__and3_1 _07450_ (.A(\core_pipeline.memory_to_writeback_next_pc[19] ),
    .B(net506),
    .C(net509),
    .X(_03977_));
 sky130_fd_sc_hd__a221o_1 _07451_ (.A1(\core_pipeline.memory_to_writeback_load_data[19] ),
    .A2(net443),
    .B1(net439),
    .B2(\core_pipeline.memory_to_writeback_csr_data[19] ),
    .C1(_03977_),
    .X(_03978_));
 sky130_fd_sc_hd__mux2_8 _07452_ (.A0(\core_pipeline.memory_to_writeback_alu_data[19] ),
    .A1(_03978_),
    .S(net441),
    .X(_03979_));
 sky130_fd_sc_hd__mux2_1 _07453_ (.A0(net309),
    .A1(\core_pipeline.pipeline_registers.registers[19][19] ),
    .S(net260),
    .X(_00060_));
 sky130_fd_sc_hd__and3_1 _07454_ (.A(\core_pipeline.memory_to_writeback_next_pc[20] ),
    .B(net507),
    .C(\core_pipeline.memory_to_writeback_write_select[0] ),
    .X(_03980_));
 sky130_fd_sc_hd__a221o_1 _07455_ (.A1(\core_pipeline.memory_to_writeback_load_data[20] ),
    .A2(net443),
    .B1(net439),
    .B2(\core_pipeline.memory_to_writeback_csr_data[20] ),
    .C1(_03980_),
    .X(_03981_));
 sky130_fd_sc_hd__mux2_4 _07456_ (.A0(\core_pipeline.memory_to_writeback_alu_data[20] ),
    .A1(_03981_),
    .S(net441),
    .X(_03982_));
 sky130_fd_sc_hd__mux2_1 _07457_ (.A0(net306),
    .A1(\core_pipeline.pipeline_registers.registers[19][20] ),
    .S(net260),
    .X(_00061_));
 sky130_fd_sc_hd__and3_1 _07458_ (.A(\core_pipeline.memory_to_writeback_next_pc[21] ),
    .B(net507),
    .C(\core_pipeline.memory_to_writeback_write_select[0] ),
    .X(_03983_));
 sky130_fd_sc_hd__a221o_1 _07459_ (.A1(\core_pipeline.memory_to_writeback_load_data[21] ),
    .A2(net443),
    .B1(net439),
    .B2(\core_pipeline.memory_to_writeback_csr_data[21] ),
    .C1(_03983_),
    .X(_03984_));
 sky130_fd_sc_hd__mux2_8 _07460_ (.A0(\core_pipeline.memory_to_writeback_alu_data[21] ),
    .A1(_03984_),
    .S(net441),
    .X(_03985_));
 sky130_fd_sc_hd__mux2_1 _07461_ (.A0(net304),
    .A1(\core_pipeline.pipeline_registers.registers[19][21] ),
    .S(net260),
    .X(_00062_));
 sky130_fd_sc_hd__and3_1 _07462_ (.A(\core_pipeline.memory_to_writeback_next_pc[22] ),
    .B(net506),
    .C(net509),
    .X(_03986_));
 sky130_fd_sc_hd__a221o_1 _07463_ (.A1(\core_pipeline.memory_to_writeback_load_data[22] ),
    .A2(net444),
    .B1(net440),
    .B2(\core_pipeline.memory_to_writeback_csr_data[22] ),
    .C1(_03986_),
    .X(_03987_));
 sky130_fd_sc_hd__mux2_8 _07464_ (.A0(\core_pipeline.memory_to_writeback_alu_data[22] ),
    .A1(_03987_),
    .S(net441),
    .X(_03988_));
 sky130_fd_sc_hd__mux2_1 _07465_ (.A0(net302),
    .A1(\core_pipeline.pipeline_registers.registers[19][22] ),
    .S(net259),
    .X(_00063_));
 sky130_fd_sc_hd__and3_1 _07466_ (.A(\core_pipeline.memory_to_writeback_next_pc[23] ),
    .B(net506),
    .C(net509),
    .X(_03989_));
 sky130_fd_sc_hd__a221o_1 _07467_ (.A1(\core_pipeline.memory_to_writeback_load_data[23] ),
    .A2(net444),
    .B1(net440),
    .B2(\core_pipeline.memory_to_writeback_csr_data[23] ),
    .C1(_03989_),
    .X(_03990_));
 sky130_fd_sc_hd__mux2_8 _07468_ (.A0(\core_pipeline.memory_to_writeback_alu_data[23] ),
    .A1(_03990_),
    .S(net442),
    .X(_03991_));
 sky130_fd_sc_hd__mux2_1 _07469_ (.A0(net299),
    .A1(\core_pipeline.pipeline_registers.registers[19][23] ),
    .S(net260),
    .X(_00064_));
 sky130_fd_sc_hd__and3_1 _07470_ (.A(\core_pipeline.memory_to_writeback_next_pc[24] ),
    .B(net506),
    .C(net509),
    .X(_03992_));
 sky130_fd_sc_hd__a221o_1 _07471_ (.A1(\core_pipeline.memory_to_writeback_load_data[24] ),
    .A2(net443),
    .B1(net439),
    .B2(\core_pipeline.memory_to_writeback_csr_data[24] ),
    .C1(_03992_),
    .X(_03993_));
 sky130_fd_sc_hd__mux2_8 _07472_ (.A0(\core_pipeline.memory_to_writeback_alu_data[24] ),
    .A1(_03993_),
    .S(net441),
    .X(_03994_));
 sky130_fd_sc_hd__mux2_1 _07473_ (.A0(net298),
    .A1(\core_pipeline.pipeline_registers.registers[19][24] ),
    .S(net259),
    .X(_00065_));
 sky130_fd_sc_hd__and3_1 _07474_ (.A(\core_pipeline.memory_to_writeback_next_pc[25] ),
    .B(net506),
    .C(net509),
    .X(_03995_));
 sky130_fd_sc_hd__a221o_1 _07475_ (.A1(\core_pipeline.memory_to_writeback_load_data[25] ),
    .A2(net443),
    .B1(net439),
    .B2(\core_pipeline.memory_to_writeback_csr_data[25] ),
    .C1(_03995_),
    .X(_03996_));
 sky130_fd_sc_hd__mux2_8 _07476_ (.A0(\core_pipeline.memory_to_writeback_alu_data[25] ),
    .A1(_03996_),
    .S(net441),
    .X(_03997_));
 sky130_fd_sc_hd__mux2_1 _07477_ (.A0(net296),
    .A1(\core_pipeline.pipeline_registers.registers[19][25] ),
    .S(net259),
    .X(_00066_));
 sky130_fd_sc_hd__and3_1 _07478_ (.A(\core_pipeline.memory_to_writeback_next_pc[26] ),
    .B(net507),
    .C(\core_pipeline.memory_to_writeback_write_select[0] ),
    .X(_03998_));
 sky130_fd_sc_hd__a221o_1 _07479_ (.A1(\core_pipeline.memory_to_writeback_load_data[26] ),
    .A2(net443),
    .B1(net439),
    .B2(\core_pipeline.memory_to_writeback_csr_data[26] ),
    .C1(_03998_),
    .X(_03999_));
 sky130_fd_sc_hd__mux2_8 _07480_ (.A0(\core_pipeline.memory_to_writeback_alu_data[26] ),
    .A1(_03999_),
    .S(net441),
    .X(_04000_));
 sky130_fd_sc_hd__mux2_1 _07481_ (.A0(net293),
    .A1(\core_pipeline.pipeline_registers.registers[19][26] ),
    .S(net259),
    .X(_00067_));
 sky130_fd_sc_hd__and3_1 _07482_ (.A(\core_pipeline.memory_to_writeback_next_pc[27] ),
    .B(net507),
    .C(net509),
    .X(_04001_));
 sky130_fd_sc_hd__a221o_1 _07483_ (.A1(\core_pipeline.memory_to_writeback_load_data[27] ),
    .A2(net443),
    .B1(net439),
    .B2(\core_pipeline.memory_to_writeback_csr_data[27] ),
    .C1(_04001_),
    .X(_04002_));
 sky130_fd_sc_hd__mux2_8 _07484_ (.A0(\core_pipeline.memory_to_writeback_alu_data[27] ),
    .A1(_04002_),
    .S(net442),
    .X(_04003_));
 sky130_fd_sc_hd__mux2_1 _07485_ (.A0(net291),
    .A1(\core_pipeline.pipeline_registers.registers[19][27] ),
    .S(net260),
    .X(_00068_));
 sky130_fd_sc_hd__and3_1 _07486_ (.A(\core_pipeline.memory_to_writeback_next_pc[28] ),
    .B(net507),
    .C(net510),
    .X(_04004_));
 sky130_fd_sc_hd__a221o_1 _07487_ (.A1(\core_pipeline.memory_to_writeback_load_data[28] ),
    .A2(net444),
    .B1(net440),
    .B2(\core_pipeline.memory_to_writeback_csr_data[28] ),
    .C1(_04004_),
    .X(_04005_));
 sky130_fd_sc_hd__mux2_8 _07488_ (.A0(\core_pipeline.memory_to_writeback_alu_data[28] ),
    .A1(_04005_),
    .S(net442),
    .X(_04006_));
 sky130_fd_sc_hd__mux2_1 _07489_ (.A0(net290),
    .A1(\core_pipeline.pipeline_registers.registers[19][28] ),
    .S(net260),
    .X(_00069_));
 sky130_fd_sc_hd__and3_1 _07490_ (.A(\core_pipeline.memory_to_writeback_next_pc[29] ),
    .B(net507),
    .C(net510),
    .X(_04007_));
 sky130_fd_sc_hd__a221o_1 _07491_ (.A1(\core_pipeline.memory_to_writeback_load_data[29] ),
    .A2(net444),
    .B1(net440),
    .B2(\core_pipeline.memory_to_writeback_csr_data[29] ),
    .C1(_04007_),
    .X(_04008_));
 sky130_fd_sc_hd__mux2_4 _07492_ (.A0(\core_pipeline.memory_to_writeback_alu_data[29] ),
    .A1(_04008_),
    .S(net442),
    .X(_04009_));
 sky130_fd_sc_hd__mux2_1 _07493_ (.A0(net287),
    .A1(\core_pipeline.pipeline_registers.registers[19][29] ),
    .S(net260),
    .X(_00070_));
 sky130_fd_sc_hd__and3_1 _07494_ (.A(\core_pipeline.memory_to_writeback_next_pc[30] ),
    .B(net508),
    .C(net510),
    .X(_04010_));
 sky130_fd_sc_hd__a221o_1 _07495_ (.A1(\core_pipeline.memory_to_writeback_load_data[30] ),
    .A2(net444),
    .B1(net440),
    .B2(\core_pipeline.memory_to_writeback_csr_data[30] ),
    .C1(_04010_),
    .X(_04011_));
 sky130_fd_sc_hd__mux2_8 _07496_ (.A0(\core_pipeline.memory_to_writeback_alu_data[30] ),
    .A1(_04011_),
    .S(net442),
    .X(_04012_));
 sky130_fd_sc_hd__mux2_1 _07497_ (.A0(net285),
    .A1(\core_pipeline.pipeline_registers.registers[19][30] ),
    .S(net260),
    .X(_00071_));
 sky130_fd_sc_hd__and3_1 _07498_ (.A(\core_pipeline.memory_to_writeback_next_pc[31] ),
    .B(net508),
    .C(net510),
    .X(_04013_));
 sky130_fd_sc_hd__a221o_1 _07499_ (.A1(\core_pipeline.memory_to_writeback_load_data[31] ),
    .A2(net444),
    .B1(net440),
    .B2(\core_pipeline.memory_to_writeback_csr_data[31] ),
    .C1(_04013_),
    .X(_04014_));
 sky130_fd_sc_hd__mux2_8 _07500_ (.A0(\core_pipeline.memory_to_writeback_alu_data[31] ),
    .A1(_04014_),
    .S(net442),
    .X(_04015_));
 sky130_fd_sc_hd__mux2_1 _07501_ (.A0(net282),
    .A1(\core_pipeline.pipeline_registers.registers[19][31] ),
    .S(net260),
    .X(_00072_));
 sky130_fd_sc_hd__or4_1 _07502_ (.A(\core_pipeline.memory_to_writeback_csr_address[5] ),
    .B(\core_pipeline.memory_to_writeback_csr_address[4] ),
    .C(\core_pipeline.memory_to_writeback_csr_address[7] ),
    .D(\core_pipeline.memory_to_writeback_csr_address[6] ),
    .X(_04016_));
 sky130_fd_sc_hd__nand2b_2 _07503_ (.A_N(\core_pipeline.memory_to_writeback_csr_address[3] ),
    .B(\core_pipeline.memory_to_writeback_csr_address[2] ),
    .Y(_04017_));
 sky130_fd_sc_hd__or3_1 _07504_ (.A(_03482_),
    .B(_03643_),
    .C(_04016_),
    .X(_04018_));
 sky130_fd_sc_hd__or4b_4 _07505_ (.A(\core_pipeline.memory_to_writeback_csr_address[1] ),
    .B(_04017_),
    .C(_04018_),
    .D_N(\core_pipeline.memory_to_writeback_csr_address[0] ),
    .X(_04019_));
 sky130_fd_sc_hd__mux2_1 _07506_ (.A0(\core_pipeline.memory_to_writeback_alu_data[2] ),
    .A1(\core_pipeline.csr_to_fetch_trap_vector[2] ),
    .S(net236),
    .X(_00073_));
 sky130_fd_sc_hd__mux2_1 _07507_ (.A0(\core_pipeline.memory_to_writeback_alu_data[3] ),
    .A1(\core_pipeline.csr_to_fetch_trap_vector[3] ),
    .S(net236),
    .X(_00074_));
 sky130_fd_sc_hd__mux2_1 _07508_ (.A0(\core_pipeline.memory_to_writeback_alu_data[4] ),
    .A1(\core_pipeline.csr_to_fetch_trap_vector[4] ),
    .S(net236),
    .X(_00075_));
 sky130_fd_sc_hd__mux2_1 _07509_ (.A0(\core_pipeline.memory_to_writeback_alu_data[5] ),
    .A1(\core_pipeline.csr_to_fetch_trap_vector[5] ),
    .S(net236),
    .X(_00076_));
 sky130_fd_sc_hd__mux2_1 _07510_ (.A0(\core_pipeline.memory_to_writeback_alu_data[6] ),
    .A1(\core_pipeline.csr_to_fetch_trap_vector[6] ),
    .S(net236),
    .X(_00077_));
 sky130_fd_sc_hd__mux2_1 _07511_ (.A0(\core_pipeline.memory_to_writeback_alu_data[7] ),
    .A1(\core_pipeline.csr_to_fetch_trap_vector[7] ),
    .S(net236),
    .X(_00078_));
 sky130_fd_sc_hd__mux2_1 _07512_ (.A0(\core_pipeline.memory_to_writeback_alu_data[8] ),
    .A1(\core_pipeline.csr_to_fetch_trap_vector[8] ),
    .S(net235),
    .X(_00079_));
 sky130_fd_sc_hd__mux2_1 _07513_ (.A0(\core_pipeline.memory_to_writeback_alu_data[9] ),
    .A1(\core_pipeline.csr_to_fetch_trap_vector[9] ),
    .S(net235),
    .X(_00080_));
 sky130_fd_sc_hd__mux2_1 _07514_ (.A0(\core_pipeline.memory_to_writeback_alu_data[10] ),
    .A1(\core_pipeline.csr_to_fetch_trap_vector[10] ),
    .S(net235),
    .X(_00081_));
 sky130_fd_sc_hd__mux2_1 _07515_ (.A0(\core_pipeline.memory_to_writeback_alu_data[11] ),
    .A1(\core_pipeline.csr_to_fetch_trap_vector[11] ),
    .S(net235),
    .X(_00082_));
 sky130_fd_sc_hd__mux2_1 _07516_ (.A0(\core_pipeline.memory_to_writeback_alu_data[12] ),
    .A1(\core_pipeline.csr_to_fetch_trap_vector[12] ),
    .S(net235),
    .X(_00083_));
 sky130_fd_sc_hd__mux2_1 _07517_ (.A0(\core_pipeline.memory_to_writeback_alu_data[13] ),
    .A1(\core_pipeline.csr_to_fetch_trap_vector[13] ),
    .S(net235),
    .X(_00084_));
 sky130_fd_sc_hd__mux2_1 _07518_ (.A0(\core_pipeline.memory_to_writeback_alu_data[14] ),
    .A1(\core_pipeline.csr_to_fetch_trap_vector[14] ),
    .S(net235),
    .X(_00085_));
 sky130_fd_sc_hd__mux2_1 _07519_ (.A0(\core_pipeline.memory_to_writeback_alu_data[15] ),
    .A1(\core_pipeline.csr_to_fetch_trap_vector[15] ),
    .S(net235),
    .X(_00086_));
 sky130_fd_sc_hd__mux2_1 _07520_ (.A0(\core_pipeline.memory_to_writeback_alu_data[16] ),
    .A1(\core_pipeline.csr_to_fetch_trap_vector[16] ),
    .S(net235),
    .X(_00087_));
 sky130_fd_sc_hd__mux2_1 _07521_ (.A0(\core_pipeline.memory_to_writeback_alu_data[17] ),
    .A1(\core_pipeline.csr_to_fetch_trap_vector[17] ),
    .S(net235),
    .X(_00088_));
 sky130_fd_sc_hd__mux2_1 _07522_ (.A0(\core_pipeline.memory_to_writeback_alu_data[18] ),
    .A1(\core_pipeline.csr_to_fetch_trap_vector[18] ),
    .S(net235),
    .X(_00089_));
 sky130_fd_sc_hd__mux2_1 _07523_ (.A0(\core_pipeline.memory_to_writeback_alu_data[19] ),
    .A1(\core_pipeline.csr_to_fetch_trap_vector[19] ),
    .S(net235),
    .X(_00090_));
 sky130_fd_sc_hd__mux2_1 _07524_ (.A0(\core_pipeline.memory_to_writeback_alu_data[20] ),
    .A1(\core_pipeline.csr_to_fetch_trap_vector[20] ),
    .S(net236),
    .X(_00091_));
 sky130_fd_sc_hd__mux2_1 _07525_ (.A0(\core_pipeline.memory_to_writeback_alu_data[21] ),
    .A1(\core_pipeline.csr_to_fetch_trap_vector[21] ),
    .S(net235),
    .X(_00092_));
 sky130_fd_sc_hd__mux2_1 _07526_ (.A0(\core_pipeline.memory_to_writeback_alu_data[22] ),
    .A1(\core_pipeline.csr_to_fetch_trap_vector[22] ),
    .S(net235),
    .X(_00093_));
 sky130_fd_sc_hd__mux2_1 _07527_ (.A0(\core_pipeline.memory_to_writeback_alu_data[23] ),
    .A1(\core_pipeline.csr_to_fetch_trap_vector[23] ),
    .S(net235),
    .X(_00094_));
 sky130_fd_sc_hd__mux2_1 _07528_ (.A0(\core_pipeline.memory_to_writeback_alu_data[24] ),
    .A1(\core_pipeline.csr_to_fetch_trap_vector[24] ),
    .S(net235),
    .X(_00095_));
 sky130_fd_sc_hd__mux2_1 _07529_ (.A0(\core_pipeline.memory_to_writeback_alu_data[25] ),
    .A1(\core_pipeline.csr_to_fetch_trap_vector[25] ),
    .S(net235),
    .X(_00096_));
 sky130_fd_sc_hd__mux2_1 _07530_ (.A0(\core_pipeline.memory_to_writeback_alu_data[26] ),
    .A1(\core_pipeline.csr_to_fetch_trap_vector[26] ),
    .S(net236),
    .X(_00097_));
 sky130_fd_sc_hd__mux2_1 _07531_ (.A0(\core_pipeline.memory_to_writeback_alu_data[27] ),
    .A1(\core_pipeline.csr_to_fetch_trap_vector[27] ),
    .S(net236),
    .X(_00098_));
 sky130_fd_sc_hd__mux2_1 _07532_ (.A0(\core_pipeline.memory_to_writeback_alu_data[28] ),
    .A1(\core_pipeline.csr_to_fetch_trap_vector[28] ),
    .S(net236),
    .X(_00099_));
 sky130_fd_sc_hd__mux2_1 _07533_ (.A0(\core_pipeline.memory_to_writeback_alu_data[29] ),
    .A1(\core_pipeline.csr_to_fetch_trap_vector[29] ),
    .S(net236),
    .X(_00100_));
 sky130_fd_sc_hd__mux2_1 _07534_ (.A0(\core_pipeline.memory_to_writeback_alu_data[30] ),
    .A1(\core_pipeline.csr_to_fetch_trap_vector[30] ),
    .S(net236),
    .X(_00101_));
 sky130_fd_sc_hd__mux2_1 _07535_ (.A0(\core_pipeline.memory_to_writeback_alu_data[31] ),
    .A1(\core_pipeline.csr_to_fetch_trap_vector[31] ),
    .S(net236),
    .X(_00102_));
 sky130_fd_sc_hd__and4b_1 _07536_ (.A_N(\core_pipeline.memory_to_writeback_csr_address[10] ),
    .B(\core_pipeline.memory_to_writeback_csr_address[11] ),
    .C(\core_pipeline.memory_to_writeback_csr_address[9] ),
    .D(\core_pipeline.memory_to_writeback_csr_address[8] ),
    .X(_04020_));
 sky130_fd_sc_hd__nand2b_1 _07537_ (.A_N(_04016_),
    .B(_04020_),
    .Y(_04021_));
 sky130_fd_sc_hd__or2_4 _07538_ (.A(_03648_),
    .B(_04021_),
    .X(_04022_));
 sky130_fd_sc_hd__nand2_1 _07539_ (.A(\core_pipeline.pipeline_csr.cycle[0] ),
    .B(net231),
    .Y(_04023_));
 sky130_fd_sc_hd__o211a_1 _07540_ (.A1(\core_pipeline.memory_to_writeback_alu_data[0] ),
    .A2(net231),
    .B1(_04023_),
    .C1(net639),
    .X(_00103_));
 sky130_fd_sc_hd__xnor2_1 _07541_ (.A(\core_pipeline.pipeline_csr.cycle[1] ),
    .B(\core_pipeline.pipeline_csr.cycle[0] ),
    .Y(_04024_));
 sky130_fd_sc_hd__nand2_1 _07542_ (.A(net231),
    .B(_04024_),
    .Y(_04025_));
 sky130_fd_sc_hd__o211a_1 _07543_ (.A1(\core_pipeline.memory_to_writeback_alu_data[1] ),
    .A2(net231),
    .B1(_04025_),
    .C1(net639),
    .X(_00104_));
 sky130_fd_sc_hd__and3_1 _07544_ (.A(\core_pipeline.pipeline_csr.cycle[2] ),
    .B(\core_pipeline.pipeline_csr.cycle[1] ),
    .C(\core_pipeline.pipeline_csr.cycle[0] ),
    .X(_04026_));
 sky130_fd_sc_hd__a21oi_1 _07545_ (.A1(\core_pipeline.pipeline_csr.cycle[1] ),
    .A2(\core_pipeline.pipeline_csr.cycle[0] ),
    .B1(\core_pipeline.pipeline_csr.cycle[2] ),
    .Y(_04027_));
 sky130_fd_sc_hd__o21ai_1 _07546_ (.A1(_04026_),
    .A2(_04027_),
    .B1(net231),
    .Y(_04028_));
 sky130_fd_sc_hd__o211a_1 _07547_ (.A1(\core_pipeline.memory_to_writeback_alu_data[2] ),
    .A2(net231),
    .B1(_04028_),
    .C1(net639),
    .X(_00105_));
 sky130_fd_sc_hd__and4_2 _07548_ (.A(\core_pipeline.pipeline_csr.cycle[3] ),
    .B(\core_pipeline.pipeline_csr.cycle[2] ),
    .C(\core_pipeline.pipeline_csr.cycle[1] ),
    .D(\core_pipeline.pipeline_csr.cycle[0] ),
    .X(_04029_));
 sky130_fd_sc_hd__nor2_1 _07549_ (.A(\core_pipeline.pipeline_csr.cycle[3] ),
    .B(_04026_),
    .Y(_04030_));
 sky130_fd_sc_hd__o21ai_1 _07550_ (.A1(_04029_),
    .A2(_04030_),
    .B1(net231),
    .Y(_04031_));
 sky130_fd_sc_hd__o211a_1 _07551_ (.A1(\core_pipeline.memory_to_writeback_alu_data[3] ),
    .A2(net231),
    .B1(_04031_),
    .C1(net639),
    .X(_00106_));
 sky130_fd_sc_hd__xnor2_1 _07552_ (.A(\core_pipeline.pipeline_csr.cycle[4] ),
    .B(_04029_),
    .Y(_04032_));
 sky130_fd_sc_hd__nand2_1 _07553_ (.A(net231),
    .B(_04032_),
    .Y(_04033_));
 sky130_fd_sc_hd__o211a_1 _07554_ (.A1(\core_pipeline.memory_to_writeback_alu_data[4] ),
    .A2(net231),
    .B1(_04033_),
    .C1(net639),
    .X(_00107_));
 sky130_fd_sc_hd__and3_1 _07555_ (.A(\core_pipeline.pipeline_csr.cycle[5] ),
    .B(\core_pipeline.pipeline_csr.cycle[4] ),
    .C(_04029_),
    .X(_04034_));
 sky130_fd_sc_hd__a21oi_1 _07556_ (.A1(\core_pipeline.pipeline_csr.cycle[4] ),
    .A2(_04029_),
    .B1(\core_pipeline.pipeline_csr.cycle[5] ),
    .Y(_04035_));
 sky130_fd_sc_hd__o21ai_1 _07557_ (.A1(_04034_),
    .A2(_04035_),
    .B1(net232),
    .Y(_04036_));
 sky130_fd_sc_hd__o211a_1 _07558_ (.A1(\core_pipeline.memory_to_writeback_alu_data[5] ),
    .A2(net232),
    .B1(_04036_),
    .C1(net640),
    .X(_00108_));
 sky130_fd_sc_hd__and4_4 _07559_ (.A(\core_pipeline.pipeline_csr.cycle[6] ),
    .B(\core_pipeline.pipeline_csr.cycle[5] ),
    .C(\core_pipeline.pipeline_csr.cycle[4] ),
    .D(_04029_),
    .X(_04037_));
 sky130_fd_sc_hd__nor2_1 _07560_ (.A(\core_pipeline.pipeline_csr.cycle[6] ),
    .B(_04034_),
    .Y(_04038_));
 sky130_fd_sc_hd__o21ai_1 _07561_ (.A1(_04037_),
    .A2(_04038_),
    .B1(net232),
    .Y(_04039_));
 sky130_fd_sc_hd__o211a_1 _07562_ (.A1(\core_pipeline.memory_to_writeback_alu_data[6] ),
    .A2(net232),
    .B1(_04039_),
    .C1(net640),
    .X(_00109_));
 sky130_fd_sc_hd__nand2_2 _07563_ (.A(\core_pipeline.pipeline_csr.cycle[7] ),
    .B(_04037_),
    .Y(_04040_));
 sky130_fd_sc_hd__or2_1 _07564_ (.A(\core_pipeline.pipeline_csr.cycle[7] ),
    .B(_04037_),
    .X(_04041_));
 sky130_fd_sc_hd__a21bo_1 _07565_ (.A1(_04040_),
    .A2(_04041_),
    .B1_N(net231),
    .X(_04042_));
 sky130_fd_sc_hd__o211a_1 _07566_ (.A1(\core_pipeline.memory_to_writeback_alu_data[7] ),
    .A2(net231),
    .B1(_04042_),
    .C1(net638),
    .X(_00110_));
 sky130_fd_sc_hd__xnor2_1 _07567_ (.A(_03391_),
    .B(_04040_),
    .Y(_04043_));
 sky130_fd_sc_hd__nand2_1 _07568_ (.A(net234),
    .B(_04043_),
    .Y(_04044_));
 sky130_fd_sc_hd__o211a_1 _07569_ (.A1(\core_pipeline.memory_to_writeback_alu_data[8] ),
    .A2(net234),
    .B1(_04044_),
    .C1(net643),
    .X(_00111_));
 sky130_fd_sc_hd__o21a_1 _07570_ (.A1(_03391_),
    .A2(_04040_),
    .B1(_03389_),
    .X(_04045_));
 sky130_fd_sc_hd__nor2_1 _07571_ (.A(_03389_),
    .B(_03391_),
    .Y(_04046_));
 sky130_fd_sc_hd__and3_1 _07572_ (.A(\core_pipeline.pipeline_csr.cycle[7] ),
    .B(_04037_),
    .C(_04046_),
    .X(_04047_));
 sky130_fd_sc_hd__o21ai_1 _07573_ (.A1(_04045_),
    .A2(_04047_),
    .B1(net234),
    .Y(_04048_));
 sky130_fd_sc_hd__o211a_1 _07574_ (.A1(\core_pipeline.memory_to_writeback_alu_data[9] ),
    .A2(net234),
    .B1(_04048_),
    .C1(net637),
    .X(_00112_));
 sky130_fd_sc_hd__nor2_1 _07575_ (.A(\core_pipeline.pipeline_csr.cycle[10] ),
    .B(_04047_),
    .Y(_04049_));
 sky130_fd_sc_hd__and4_2 _07576_ (.A(\core_pipeline.pipeline_csr.cycle[10] ),
    .B(\core_pipeline.pipeline_csr.cycle[7] ),
    .C(_04037_),
    .D(_04046_),
    .X(_04050_));
 sky130_fd_sc_hd__o21ai_1 _07577_ (.A1(_04049_),
    .A2(_04050_),
    .B1(net234),
    .Y(_04051_));
 sky130_fd_sc_hd__o211a_1 _07578_ (.A1(\core_pipeline.memory_to_writeback_alu_data[10] ),
    .A2(net234),
    .B1(_04051_),
    .C1(net643),
    .X(_00113_));
 sky130_fd_sc_hd__nor2_1 _07579_ (.A(\core_pipeline.pipeline_csr.cycle[11] ),
    .B(_04050_),
    .Y(_04052_));
 sky130_fd_sc_hd__and2_1 _07580_ (.A(\core_pipeline.pipeline_csr.cycle[11] ),
    .B(_04050_),
    .X(_04053_));
 sky130_fd_sc_hd__o21ai_1 _07581_ (.A1(_04052_),
    .A2(_04053_),
    .B1(net233),
    .Y(_04054_));
 sky130_fd_sc_hd__o211a_1 _07582_ (.A1(\core_pipeline.memory_to_writeback_alu_data[11] ),
    .A2(net233),
    .B1(_04054_),
    .C1(net636),
    .X(_00114_));
 sky130_fd_sc_hd__nor2_1 _07583_ (.A(\core_pipeline.pipeline_csr.cycle[12] ),
    .B(_04053_),
    .Y(_04055_));
 sky130_fd_sc_hd__and3_1 _07584_ (.A(\core_pipeline.pipeline_csr.cycle[12] ),
    .B(\core_pipeline.pipeline_csr.cycle[11] ),
    .C(_04050_),
    .X(_04056_));
 sky130_fd_sc_hd__o21ai_1 _07585_ (.A1(_04055_),
    .A2(_04056_),
    .B1(net233),
    .Y(_04057_));
 sky130_fd_sc_hd__o211a_1 _07586_ (.A1(\core_pipeline.memory_to_writeback_alu_data[12] ),
    .A2(net233),
    .B1(_04057_),
    .C1(net636),
    .X(_00115_));
 sky130_fd_sc_hd__nor2_1 _07587_ (.A(\core_pipeline.pipeline_csr.cycle[13] ),
    .B(_04056_),
    .Y(_04058_));
 sky130_fd_sc_hd__and4_4 _07588_ (.A(\core_pipeline.pipeline_csr.cycle[13] ),
    .B(\core_pipeline.pipeline_csr.cycle[12] ),
    .C(\core_pipeline.pipeline_csr.cycle[11] ),
    .D(_04050_),
    .X(_04059_));
 sky130_fd_sc_hd__o21ai_1 _07589_ (.A1(_04058_),
    .A2(_04059_),
    .B1(net233),
    .Y(_04060_));
 sky130_fd_sc_hd__o211a_1 _07590_ (.A1(\core_pipeline.memory_to_writeback_alu_data[13] ),
    .A2(net233),
    .B1(_04060_),
    .C1(net636),
    .X(_00116_));
 sky130_fd_sc_hd__xnor2_1 _07591_ (.A(\core_pipeline.pipeline_csr.cycle[14] ),
    .B(_04059_),
    .Y(_04061_));
 sky130_fd_sc_hd__nand2_1 _07592_ (.A(net233),
    .B(_04061_),
    .Y(_04062_));
 sky130_fd_sc_hd__o211a_1 _07593_ (.A1(\core_pipeline.memory_to_writeback_alu_data[14] ),
    .A2(net233),
    .B1(_04062_),
    .C1(net646),
    .X(_00117_));
 sky130_fd_sc_hd__a21oi_1 _07594_ (.A1(\core_pipeline.pipeline_csr.cycle[14] ),
    .A2(_04059_),
    .B1(\core_pipeline.pipeline_csr.cycle[15] ),
    .Y(_04063_));
 sky130_fd_sc_hd__nor2_1 _07595_ (.A(_03377_),
    .B(_03379_),
    .Y(_04064_));
 sky130_fd_sc_hd__and2_2 _07596_ (.A(_04059_),
    .B(_04064_),
    .X(_04065_));
 sky130_fd_sc_hd__o21ai_1 _07597_ (.A1(_04063_),
    .A2(_04065_),
    .B1(net233),
    .Y(_04066_));
 sky130_fd_sc_hd__o211a_1 _07598_ (.A1(\core_pipeline.memory_to_writeback_alu_data[15] ),
    .A2(net233),
    .B1(_04066_),
    .C1(net646),
    .X(_00118_));
 sky130_fd_sc_hd__xnor2_1 _07599_ (.A(\core_pipeline.pipeline_csr.cycle[16] ),
    .B(_04065_),
    .Y(_04067_));
 sky130_fd_sc_hd__nand2_1 _07600_ (.A(net233),
    .B(_04067_),
    .Y(_04068_));
 sky130_fd_sc_hd__o211a_1 _07601_ (.A1(\core_pipeline.memory_to_writeback_alu_data[16] ),
    .A2(net233),
    .B1(_04068_),
    .C1(net643),
    .X(_00119_));
 sky130_fd_sc_hd__a21oi_1 _07602_ (.A1(\core_pipeline.pipeline_csr.cycle[16] ),
    .A2(_04065_),
    .B1(\core_pipeline.pipeline_csr.cycle[17] ),
    .Y(_04069_));
 sky130_fd_sc_hd__and4_2 _07603_ (.A(\core_pipeline.pipeline_csr.cycle[17] ),
    .B(\core_pipeline.pipeline_csr.cycle[16] ),
    .C(_04059_),
    .D(_04064_),
    .X(_04070_));
 sky130_fd_sc_hd__o21ai_1 _07604_ (.A1(_04069_),
    .A2(_04070_),
    .B1(net233),
    .Y(_04071_));
 sky130_fd_sc_hd__o211a_1 _07605_ (.A1(\core_pipeline.memory_to_writeback_alu_data[17] ),
    .A2(net233),
    .B1(_04071_),
    .C1(net643),
    .X(_00120_));
 sky130_fd_sc_hd__xnor2_1 _07606_ (.A(\core_pipeline.pipeline_csr.cycle[18] ),
    .B(_04070_),
    .Y(_04072_));
 sky130_fd_sc_hd__nand2_1 _07607_ (.A(net233),
    .B(_04072_),
    .Y(_04073_));
 sky130_fd_sc_hd__o211a_1 _07608_ (.A1(\core_pipeline.memory_to_writeback_alu_data[18] ),
    .A2(net233),
    .B1(_04073_),
    .C1(net645),
    .X(_00121_));
 sky130_fd_sc_hd__a21oi_1 _07609_ (.A1(\core_pipeline.pipeline_csr.cycle[18] ),
    .A2(_04070_),
    .B1(\core_pipeline.pipeline_csr.cycle[19] ),
    .Y(_04074_));
 sky130_fd_sc_hd__and3_2 _07610_ (.A(\core_pipeline.pipeline_csr.cycle[19] ),
    .B(\core_pipeline.pipeline_csr.cycle[18] ),
    .C(_04070_),
    .X(_04075_));
 sky130_fd_sc_hd__o21ai_1 _07611_ (.A1(_04074_),
    .A2(_04075_),
    .B1(_04022_),
    .Y(_04076_));
 sky130_fd_sc_hd__o211a_1 _07612_ (.A1(\core_pipeline.memory_to_writeback_alu_data[19] ),
    .A2(net233),
    .B1(_04076_),
    .C1(net645),
    .X(_00122_));
 sky130_fd_sc_hd__xnor2_1 _07613_ (.A(\core_pipeline.pipeline_csr.cycle[20] ),
    .B(_04075_),
    .Y(_04077_));
 sky130_fd_sc_hd__nand2_1 _07614_ (.A(_04022_),
    .B(_04077_),
    .Y(_04078_));
 sky130_fd_sc_hd__o211a_1 _07615_ (.A1(\core_pipeline.memory_to_writeback_alu_data[20] ),
    .A2(_04022_),
    .B1(_04078_),
    .C1(net645),
    .X(_00123_));
 sky130_fd_sc_hd__a21o_1 _07616_ (.A1(\core_pipeline.pipeline_csr.cycle[20] ),
    .A2(_04075_),
    .B1(\core_pipeline.pipeline_csr.cycle[21] ),
    .X(_04079_));
 sky130_fd_sc_hd__nand3_2 _07617_ (.A(\core_pipeline.pipeline_csr.cycle[21] ),
    .B(\core_pipeline.pipeline_csr.cycle[20] ),
    .C(_04075_),
    .Y(_04080_));
 sky130_fd_sc_hd__a21bo_1 _07618_ (.A1(_04079_),
    .A2(_04080_),
    .B1_N(net234),
    .X(_04081_));
 sky130_fd_sc_hd__o211a_1 _07619_ (.A1(\core_pipeline.memory_to_writeback_alu_data[21] ),
    .A2(net234),
    .B1(_04081_),
    .C1(net643),
    .X(_00124_));
 sky130_fd_sc_hd__and2_1 _07620_ (.A(_03363_),
    .B(_04080_),
    .X(_04082_));
 sky130_fd_sc_hd__nor2_1 _07621_ (.A(_03363_),
    .B(_04080_),
    .Y(_04083_));
 sky130_fd_sc_hd__o21ai_1 _07622_ (.A1(_04082_),
    .A2(_04083_),
    .B1(net234),
    .Y(_04084_));
 sky130_fd_sc_hd__o211a_1 _07623_ (.A1(\core_pipeline.memory_to_writeback_alu_data[22] ),
    .A2(net234),
    .B1(_04084_),
    .C1(net644),
    .X(_00125_));
 sky130_fd_sc_hd__nor2_1 _07624_ (.A(\core_pipeline.pipeline_csr.cycle[23] ),
    .B(_04083_),
    .Y(_04085_));
 sky130_fd_sc_hd__and2_2 _07625_ (.A(\core_pipeline.pipeline_csr.cycle[23] ),
    .B(_04083_),
    .X(_04086_));
 sky130_fd_sc_hd__o21ai_1 _07626_ (.A1(_04085_),
    .A2(_04086_),
    .B1(net234),
    .Y(_04087_));
 sky130_fd_sc_hd__o211a_1 _07627_ (.A1(\core_pipeline.memory_to_writeback_alu_data[23] ),
    .A2(net234),
    .B1(_04087_),
    .C1(net644),
    .X(_00126_));
 sky130_fd_sc_hd__xnor2_1 _07628_ (.A(\core_pipeline.pipeline_csr.cycle[24] ),
    .B(_04086_),
    .Y(_04088_));
 sky130_fd_sc_hd__nand2_1 _07629_ (.A(net234),
    .B(_04088_),
    .Y(_04089_));
 sky130_fd_sc_hd__o211a_1 _07630_ (.A1(\core_pipeline.memory_to_writeback_alu_data[24] ),
    .A2(net234),
    .B1(_04089_),
    .C1(net644),
    .X(_00127_));
 sky130_fd_sc_hd__a21oi_1 _07631_ (.A1(\core_pipeline.pipeline_csr.cycle[24] ),
    .A2(_04086_),
    .B1(\core_pipeline.pipeline_csr.cycle[25] ),
    .Y(_04090_));
 sky130_fd_sc_hd__and3_1 _07632_ (.A(\core_pipeline.pipeline_csr.cycle[25] ),
    .B(\core_pipeline.pipeline_csr.cycle[24] ),
    .C(_04086_),
    .X(_04091_));
 sky130_fd_sc_hd__o21ai_1 _07633_ (.A1(_04090_),
    .A2(_04091_),
    .B1(net234),
    .Y(_04092_));
 sky130_fd_sc_hd__o211a_1 _07634_ (.A1(\core_pipeline.memory_to_writeback_alu_data[25] ),
    .A2(net234),
    .B1(_04092_),
    .C1(net644),
    .X(_00128_));
 sky130_fd_sc_hd__xnor2_1 _07635_ (.A(\core_pipeline.pipeline_csr.cycle[26] ),
    .B(_04091_),
    .Y(_04093_));
 sky130_fd_sc_hd__nand2_1 _07636_ (.A(net232),
    .B(_04093_),
    .Y(_04094_));
 sky130_fd_sc_hd__o211a_1 _07637_ (.A1(\core_pipeline.memory_to_writeback_alu_data[26] ),
    .A2(net232),
    .B1(_04094_),
    .C1(net642),
    .X(_00129_));
 sky130_fd_sc_hd__a21oi_1 _07638_ (.A1(\core_pipeline.pipeline_csr.cycle[26] ),
    .A2(_04091_),
    .B1(\core_pipeline.pipeline_csr.cycle[27] ),
    .Y(_04095_));
 sky130_fd_sc_hd__and4_1 _07639_ (.A(\core_pipeline.pipeline_csr.cycle[27] ),
    .B(\core_pipeline.pipeline_csr.cycle[26] ),
    .C(\core_pipeline.pipeline_csr.cycle[25] ),
    .D(\core_pipeline.pipeline_csr.cycle[24] ),
    .X(_04096_));
 sky130_fd_sc_hd__and2_2 _07640_ (.A(_04086_),
    .B(_04096_),
    .X(_04097_));
 sky130_fd_sc_hd__o21ai_1 _07641_ (.A1(_04095_),
    .A2(_04097_),
    .B1(net232),
    .Y(_04098_));
 sky130_fd_sc_hd__o211a_1 _07642_ (.A1(\core_pipeline.memory_to_writeback_alu_data[27] ),
    .A2(net232),
    .B1(_04098_),
    .C1(net642),
    .X(_00130_));
 sky130_fd_sc_hd__xnor2_1 _07643_ (.A(\core_pipeline.pipeline_csr.cycle[28] ),
    .B(_04097_),
    .Y(_04099_));
 sky130_fd_sc_hd__nand2_1 _07644_ (.A(net231),
    .B(_04099_),
    .Y(_04100_));
 sky130_fd_sc_hd__o211a_1 _07645_ (.A1(\core_pipeline.memory_to_writeback_alu_data[28] ),
    .A2(net231),
    .B1(_04100_),
    .C1(net641),
    .X(_00131_));
 sky130_fd_sc_hd__a21oi_1 _07646_ (.A1(\core_pipeline.pipeline_csr.cycle[28] ),
    .A2(_04097_),
    .B1(\core_pipeline.pipeline_csr.cycle[29] ),
    .Y(_04101_));
 sky130_fd_sc_hd__and3_2 _07647_ (.A(\core_pipeline.pipeline_csr.cycle[29] ),
    .B(\core_pipeline.pipeline_csr.cycle[28] ),
    .C(_04097_),
    .X(_04102_));
 sky130_fd_sc_hd__o21ai_1 _07648_ (.A1(_04101_),
    .A2(_04102_),
    .B1(net232),
    .Y(_04103_));
 sky130_fd_sc_hd__o211a_1 _07649_ (.A1(\core_pipeline.memory_to_writeback_alu_data[29] ),
    .A2(net231),
    .B1(_04103_),
    .C1(net641),
    .X(_00132_));
 sky130_fd_sc_hd__xnor2_1 _07650_ (.A(\core_pipeline.pipeline_csr.cycle[30] ),
    .B(_04102_),
    .Y(_04104_));
 sky130_fd_sc_hd__nand2_1 _07651_ (.A(net232),
    .B(_04104_),
    .Y(_04105_));
 sky130_fd_sc_hd__o211a_1 _07652_ (.A1(\core_pipeline.memory_to_writeback_alu_data[30] ),
    .A2(net232),
    .B1(_04105_),
    .C1(net642),
    .X(_00133_));
 sky130_fd_sc_hd__a21oi_1 _07653_ (.A1(\core_pipeline.pipeline_csr.cycle[30] ),
    .A2(_04102_),
    .B1(\core_pipeline.pipeline_csr.cycle[31] ),
    .Y(_04106_));
 sky130_fd_sc_hd__and4_1 _07654_ (.A(\core_pipeline.pipeline_csr.cycle[31] ),
    .B(\core_pipeline.pipeline_csr.cycle[30] ),
    .C(\core_pipeline.pipeline_csr.cycle[29] ),
    .D(\core_pipeline.pipeline_csr.cycle[28] ),
    .X(_04107_));
 sky130_fd_sc_hd__and3_2 _07655_ (.A(_04086_),
    .B(_04096_),
    .C(_04107_),
    .X(_04108_));
 sky130_fd_sc_hd__o21ai_1 _07656_ (.A1(_04106_),
    .A2(_04108_),
    .B1(net231),
    .Y(_04109_));
 sky130_fd_sc_hd__o211a_1 _07657_ (.A1(\core_pipeline.memory_to_writeback_alu_data[31] ),
    .A2(net231),
    .B1(_04109_),
    .C1(net641),
    .X(_00134_));
 sky130_fd_sc_hd__nand2_2 _07658_ (.A(\core_pipeline.memory_to_writeback_csr_address[7] ),
    .B(_04020_),
    .Y(_04110_));
 sky130_fd_sc_hd__nor4_4 _07659_ (.A(\core_pipeline.memory_to_writeback_csr_address[5] ),
    .B(\core_pipeline.memory_to_writeback_csr_address[4] ),
    .C(\core_pipeline.memory_to_writeback_csr_address[6] ),
    .D(_04110_),
    .Y(_04111_));
 sky130_fd_sc_hd__nand2_8 _07660_ (.A(_03647_),
    .B(net281),
    .Y(_04112_));
 sky130_fd_sc_hd__xnor2_1 _07661_ (.A(\core_pipeline.pipeline_csr.cycle[32] ),
    .B(_04108_),
    .Y(_04113_));
 sky130_fd_sc_hd__nand2_1 _07662_ (.A(net227),
    .B(_04113_),
    .Y(_04114_));
 sky130_fd_sc_hd__o211a_1 _07663_ (.A1(\core_pipeline.memory_to_writeback_alu_data[0] ),
    .A2(net227),
    .B1(_04114_),
    .C1(net641),
    .X(_00135_));
 sky130_fd_sc_hd__a21oi_1 _07664_ (.A1(\core_pipeline.pipeline_csr.cycle[32] ),
    .A2(_04108_),
    .B1(\core_pipeline.pipeline_csr.cycle[33] ),
    .Y(_04115_));
 sky130_fd_sc_hd__and3_2 _07665_ (.A(\core_pipeline.pipeline_csr.cycle[33] ),
    .B(\core_pipeline.pipeline_csr.cycle[32] ),
    .C(_04108_),
    .X(_04116_));
 sky130_fd_sc_hd__o21ai_1 _07666_ (.A1(_04115_),
    .A2(_04116_),
    .B1(net227),
    .Y(_04117_));
 sky130_fd_sc_hd__o211a_1 _07667_ (.A1(\core_pipeline.memory_to_writeback_alu_data[1] ),
    .A2(net227),
    .B1(_04117_),
    .C1(net641),
    .X(_00136_));
 sky130_fd_sc_hd__xnor2_1 _07668_ (.A(\core_pipeline.pipeline_csr.cycle[34] ),
    .B(_04116_),
    .Y(_04118_));
 sky130_fd_sc_hd__nand2_1 _07669_ (.A(net227),
    .B(_04118_),
    .Y(_04119_));
 sky130_fd_sc_hd__o211a_1 _07670_ (.A1(\core_pipeline.memory_to_writeback_alu_data[2] ),
    .A2(net227),
    .B1(_04119_),
    .C1(net641),
    .X(_00137_));
 sky130_fd_sc_hd__a21oi_1 _07671_ (.A1(\core_pipeline.pipeline_csr.cycle[34] ),
    .A2(_04116_),
    .B1(\core_pipeline.pipeline_csr.cycle[35] ),
    .Y(_04120_));
 sky130_fd_sc_hd__and3_2 _07672_ (.A(\core_pipeline.pipeline_csr.cycle[35] ),
    .B(\core_pipeline.pipeline_csr.cycle[34] ),
    .C(_04116_),
    .X(_04121_));
 sky130_fd_sc_hd__o21ai_1 _07673_ (.A1(_04120_),
    .A2(_04121_),
    .B1(net228),
    .Y(_04122_));
 sky130_fd_sc_hd__o211a_1 _07674_ (.A1(\core_pipeline.memory_to_writeback_alu_data[3] ),
    .A2(net228),
    .B1(_04122_),
    .C1(net639),
    .X(_00138_));
 sky130_fd_sc_hd__xnor2_1 _07675_ (.A(\core_pipeline.pipeline_csr.cycle[36] ),
    .B(_04121_),
    .Y(_04123_));
 sky130_fd_sc_hd__nand2_1 _07676_ (.A(net228),
    .B(_04123_),
    .Y(_04124_));
 sky130_fd_sc_hd__o211a_1 _07677_ (.A1(\core_pipeline.memory_to_writeback_alu_data[4] ),
    .A2(net228),
    .B1(_04124_),
    .C1(net639),
    .X(_00139_));
 sky130_fd_sc_hd__a21oi_1 _07678_ (.A1(\core_pipeline.pipeline_csr.cycle[36] ),
    .A2(_04121_),
    .B1(\core_pipeline.pipeline_csr.cycle[37] ),
    .Y(_04125_));
 sky130_fd_sc_hd__and3_2 _07679_ (.A(\core_pipeline.pipeline_csr.cycle[37] ),
    .B(\core_pipeline.pipeline_csr.cycle[36] ),
    .C(_04121_),
    .X(_04126_));
 sky130_fd_sc_hd__o21ai_1 _07680_ (.A1(_04125_),
    .A2(_04126_),
    .B1(net228),
    .Y(_04127_));
 sky130_fd_sc_hd__o211a_1 _07681_ (.A1(\core_pipeline.memory_to_writeback_alu_data[5] ),
    .A2(net228),
    .B1(_04127_),
    .C1(net640),
    .X(_00140_));
 sky130_fd_sc_hd__nor2_1 _07682_ (.A(\core_pipeline.pipeline_csr.cycle[38] ),
    .B(_04126_),
    .Y(_04128_));
 sky130_fd_sc_hd__and2_1 _07683_ (.A(\core_pipeline.pipeline_csr.cycle[38] ),
    .B(_04126_),
    .X(_04129_));
 sky130_fd_sc_hd__o21ai_1 _07684_ (.A1(_04128_),
    .A2(_04129_),
    .B1(net228),
    .Y(_04130_));
 sky130_fd_sc_hd__o211a_1 _07685_ (.A1(\core_pipeline.memory_to_writeback_alu_data[6] ),
    .A2(net228),
    .B1(_04130_),
    .C1(net640),
    .X(_00141_));
 sky130_fd_sc_hd__nor2_1 _07686_ (.A(\core_pipeline.pipeline_csr.cycle[39] ),
    .B(_04129_),
    .Y(_04131_));
 sky130_fd_sc_hd__and3_4 _07687_ (.A(\core_pipeline.pipeline_csr.cycle[39] ),
    .B(\core_pipeline.pipeline_csr.cycle[38] ),
    .C(_04126_),
    .X(_04132_));
 sky130_fd_sc_hd__o21ai_1 _07688_ (.A1(_04131_),
    .A2(_04132_),
    .B1(net228),
    .Y(_04133_));
 sky130_fd_sc_hd__o211a_1 _07689_ (.A1(\core_pipeline.memory_to_writeback_alu_data[7] ),
    .A2(net228),
    .B1(_04133_),
    .C1(net640),
    .X(_00142_));
 sky130_fd_sc_hd__xnor2_1 _07690_ (.A(\core_pipeline.pipeline_csr.cycle[40] ),
    .B(_04132_),
    .Y(_04134_));
 sky130_fd_sc_hd__nand2_1 _07691_ (.A(net230),
    .B(_04134_),
    .Y(_04135_));
 sky130_fd_sc_hd__o211a_1 _07692_ (.A1(\core_pipeline.memory_to_writeback_alu_data[8] ),
    .A2(net230),
    .B1(_04135_),
    .C1(net643),
    .X(_00143_));
 sky130_fd_sc_hd__a21oi_1 _07693_ (.A1(\core_pipeline.pipeline_csr.cycle[40] ),
    .A2(_04132_),
    .B1(\core_pipeline.pipeline_csr.cycle[41] ),
    .Y(_04136_));
 sky130_fd_sc_hd__and3_2 _07694_ (.A(\core_pipeline.pipeline_csr.cycle[41] ),
    .B(\core_pipeline.pipeline_csr.cycle[40] ),
    .C(_04132_),
    .X(_04137_));
 sky130_fd_sc_hd__o21ai_1 _07695_ (.A1(_04136_),
    .A2(_04137_),
    .B1(net230),
    .Y(_04138_));
 sky130_fd_sc_hd__o211a_1 _07696_ (.A1(\core_pipeline.memory_to_writeback_alu_data[9] ),
    .A2(net230),
    .B1(_04138_),
    .C1(net643),
    .X(_00144_));
 sky130_fd_sc_hd__xnor2_1 _07697_ (.A(\core_pipeline.pipeline_csr.cycle[42] ),
    .B(_04137_),
    .Y(_04139_));
 sky130_fd_sc_hd__nand2_1 _07698_ (.A(net230),
    .B(_04139_),
    .Y(_04140_));
 sky130_fd_sc_hd__o211a_1 _07699_ (.A1(\core_pipeline.memory_to_writeback_alu_data[10] ),
    .A2(net230),
    .B1(_04140_),
    .C1(net643),
    .X(_00145_));
 sky130_fd_sc_hd__a21oi_1 _07700_ (.A1(\core_pipeline.pipeline_csr.cycle[42] ),
    .A2(_04137_),
    .B1(\core_pipeline.pipeline_csr.cycle[43] ),
    .Y(_04141_));
 sky130_fd_sc_hd__and4_1 _07701_ (.A(\core_pipeline.pipeline_csr.cycle[43] ),
    .B(\core_pipeline.pipeline_csr.cycle[42] ),
    .C(\core_pipeline.pipeline_csr.cycle[41] ),
    .D(\core_pipeline.pipeline_csr.cycle[40] ),
    .X(_04142_));
 sky130_fd_sc_hd__and2_2 _07702_ (.A(_04132_),
    .B(_04142_),
    .X(_04143_));
 sky130_fd_sc_hd__o21ai_1 _07703_ (.A1(_04141_),
    .A2(_04143_),
    .B1(net230),
    .Y(_04144_));
 sky130_fd_sc_hd__o211a_1 _07704_ (.A1(\core_pipeline.memory_to_writeback_alu_data[11] ),
    .A2(net230),
    .B1(_04144_),
    .C1(net643),
    .X(_00146_));
 sky130_fd_sc_hd__xnor2_1 _07705_ (.A(\core_pipeline.pipeline_csr.cycle[44] ),
    .B(_04143_),
    .Y(_04145_));
 sky130_fd_sc_hd__nand2_1 _07706_ (.A(net230),
    .B(_04145_),
    .Y(_04146_));
 sky130_fd_sc_hd__o211a_1 _07707_ (.A1(\core_pipeline.memory_to_writeback_alu_data[12] ),
    .A2(net230),
    .B1(_04146_),
    .C1(net643),
    .X(_00147_));
 sky130_fd_sc_hd__a21oi_1 _07708_ (.A1(\core_pipeline.pipeline_csr.cycle[44] ),
    .A2(_04143_),
    .B1(\core_pipeline.pipeline_csr.cycle[45] ),
    .Y(_04147_));
 sky130_fd_sc_hd__and3_2 _07709_ (.A(\core_pipeline.pipeline_csr.cycle[45] ),
    .B(\core_pipeline.pipeline_csr.cycle[44] ),
    .C(_04143_),
    .X(_04148_));
 sky130_fd_sc_hd__o21ai_1 _07710_ (.A1(_04147_),
    .A2(_04148_),
    .B1(net230),
    .Y(_04149_));
 sky130_fd_sc_hd__o211a_1 _07711_ (.A1(\core_pipeline.memory_to_writeback_alu_data[13] ),
    .A2(net230),
    .B1(_04149_),
    .C1(net643),
    .X(_00148_));
 sky130_fd_sc_hd__xnor2_1 _07712_ (.A(\core_pipeline.pipeline_csr.cycle[46] ),
    .B(_04148_),
    .Y(_04150_));
 sky130_fd_sc_hd__nand2_1 _07713_ (.A(net230),
    .B(_04150_),
    .Y(_04151_));
 sky130_fd_sc_hd__o211a_1 _07714_ (.A1(\core_pipeline.memory_to_writeback_alu_data[14] ),
    .A2(net230),
    .B1(_04151_),
    .C1(net643),
    .X(_00149_));
 sky130_fd_sc_hd__a21oi_1 _07715_ (.A1(\core_pipeline.pipeline_csr.cycle[46] ),
    .A2(_04148_),
    .B1(\core_pipeline.pipeline_csr.cycle[47] ),
    .Y(_04152_));
 sky130_fd_sc_hd__and4_1 _07716_ (.A(\core_pipeline.pipeline_csr.cycle[47] ),
    .B(\core_pipeline.pipeline_csr.cycle[46] ),
    .C(\core_pipeline.pipeline_csr.cycle[45] ),
    .D(\core_pipeline.pipeline_csr.cycle[44] ),
    .X(_04153_));
 sky130_fd_sc_hd__and3_2 _07717_ (.A(_04132_),
    .B(_04142_),
    .C(_04153_),
    .X(_04154_));
 sky130_fd_sc_hd__o21ai_1 _07718_ (.A1(_04152_),
    .A2(_04154_),
    .B1(net230),
    .Y(_04155_));
 sky130_fd_sc_hd__o211a_1 _07719_ (.A1(\core_pipeline.memory_to_writeback_alu_data[15] ),
    .A2(net230),
    .B1(_04155_),
    .C1(net643),
    .X(_00150_));
 sky130_fd_sc_hd__xnor2_1 _07720_ (.A(\core_pipeline.pipeline_csr.cycle[48] ),
    .B(_04154_),
    .Y(_04156_));
 sky130_fd_sc_hd__nand2_1 _07721_ (.A(net229),
    .B(_04156_),
    .Y(_04157_));
 sky130_fd_sc_hd__o211a_1 _07722_ (.A1(\core_pipeline.memory_to_writeback_alu_data[16] ),
    .A2(net229),
    .B1(_04157_),
    .C1(net645),
    .X(_00151_));
 sky130_fd_sc_hd__a21oi_1 _07723_ (.A1(\core_pipeline.pipeline_csr.cycle[48] ),
    .A2(_04154_),
    .B1(\core_pipeline.pipeline_csr.cycle[49] ),
    .Y(_04158_));
 sky130_fd_sc_hd__and3_2 _07724_ (.A(\core_pipeline.pipeline_csr.cycle[49] ),
    .B(\core_pipeline.pipeline_csr.cycle[48] ),
    .C(_04154_),
    .X(_04159_));
 sky130_fd_sc_hd__o21ai_1 _07725_ (.A1(_04158_),
    .A2(_04159_),
    .B1(net229),
    .Y(_04160_));
 sky130_fd_sc_hd__o211a_1 _07726_ (.A1(\core_pipeline.memory_to_writeback_alu_data[17] ),
    .A2(net229),
    .B1(_04160_),
    .C1(net645),
    .X(_00152_));
 sky130_fd_sc_hd__xnor2_1 _07727_ (.A(\core_pipeline.pipeline_csr.cycle[50] ),
    .B(_04159_),
    .Y(_04161_));
 sky130_fd_sc_hd__nand2_1 _07728_ (.A(net229),
    .B(_04161_),
    .Y(_04162_));
 sky130_fd_sc_hd__o211a_1 _07729_ (.A1(\core_pipeline.memory_to_writeback_alu_data[18] ),
    .A2(net229),
    .B1(_04162_),
    .C1(net645),
    .X(_00153_));
 sky130_fd_sc_hd__a21oi_1 _07730_ (.A1(\core_pipeline.pipeline_csr.cycle[50] ),
    .A2(_04159_),
    .B1(\core_pipeline.pipeline_csr.cycle[51] ),
    .Y(_04163_));
 sky130_fd_sc_hd__and4_1 _07731_ (.A(\core_pipeline.pipeline_csr.cycle[51] ),
    .B(\core_pipeline.pipeline_csr.cycle[50] ),
    .C(\core_pipeline.pipeline_csr.cycle[49] ),
    .D(\core_pipeline.pipeline_csr.cycle[48] ),
    .X(_04164_));
 sky130_fd_sc_hd__and3_2 _07732_ (.A(_04143_),
    .B(_04153_),
    .C(_04164_),
    .X(_04165_));
 sky130_fd_sc_hd__o21ai_1 _07733_ (.A1(_04163_),
    .A2(_04165_),
    .B1(net229),
    .Y(_04166_));
 sky130_fd_sc_hd__o211a_1 _07734_ (.A1(\core_pipeline.memory_to_writeback_alu_data[19] ),
    .A2(net229),
    .B1(_04166_),
    .C1(net645),
    .X(_00154_));
 sky130_fd_sc_hd__xnor2_1 _07735_ (.A(\core_pipeline.pipeline_csr.cycle[52] ),
    .B(_04165_),
    .Y(_04167_));
 sky130_fd_sc_hd__nand2_1 _07736_ (.A(_04112_),
    .B(_04167_),
    .Y(_04168_));
 sky130_fd_sc_hd__o211a_1 _07737_ (.A1(\core_pipeline.memory_to_writeback_alu_data[20] ),
    .A2(_04112_),
    .B1(_04168_),
    .C1(net644),
    .X(_00155_));
 sky130_fd_sc_hd__a21oi_1 _07738_ (.A1(\core_pipeline.pipeline_csr.cycle[52] ),
    .A2(_04165_),
    .B1(\core_pipeline.pipeline_csr.cycle[53] ),
    .Y(_04169_));
 sky130_fd_sc_hd__and3_2 _07739_ (.A(\core_pipeline.pipeline_csr.cycle[53] ),
    .B(\core_pipeline.pipeline_csr.cycle[52] ),
    .C(_04165_),
    .X(_04170_));
 sky130_fd_sc_hd__o21ai_1 _07740_ (.A1(_04169_),
    .A2(_04170_),
    .B1(net229),
    .Y(_04171_));
 sky130_fd_sc_hd__o211a_1 _07741_ (.A1(\core_pipeline.memory_to_writeback_alu_data[21] ),
    .A2(_04112_),
    .B1(_04171_),
    .C1(net644),
    .X(_00156_));
 sky130_fd_sc_hd__xnor2_1 _07742_ (.A(\core_pipeline.pipeline_csr.cycle[54] ),
    .B(_04170_),
    .Y(_04172_));
 sky130_fd_sc_hd__nand2_1 _07743_ (.A(net229),
    .B(_04172_),
    .Y(_04173_));
 sky130_fd_sc_hd__o211a_1 _07744_ (.A1(\core_pipeline.memory_to_writeback_alu_data[22] ),
    .A2(net229),
    .B1(_04173_),
    .C1(net644),
    .X(_00157_));
 sky130_fd_sc_hd__a21oi_1 _07745_ (.A1(\core_pipeline.pipeline_csr.cycle[54] ),
    .A2(_04170_),
    .B1(\core_pipeline.pipeline_csr.cycle[55] ),
    .Y(_04174_));
 sky130_fd_sc_hd__and3_2 _07746_ (.A(\core_pipeline.pipeline_csr.cycle[55] ),
    .B(\core_pipeline.pipeline_csr.cycle[54] ),
    .C(_04170_),
    .X(_04175_));
 sky130_fd_sc_hd__o21ai_1 _07747_ (.A1(_04174_),
    .A2(_04175_),
    .B1(net229),
    .Y(_04176_));
 sky130_fd_sc_hd__o211a_1 _07748_ (.A1(\core_pipeline.memory_to_writeback_alu_data[23] ),
    .A2(net229),
    .B1(_04176_),
    .C1(net644),
    .X(_00158_));
 sky130_fd_sc_hd__xnor2_1 _07749_ (.A(\core_pipeline.pipeline_csr.cycle[56] ),
    .B(_04175_),
    .Y(_04177_));
 sky130_fd_sc_hd__nand2_1 _07750_ (.A(net229),
    .B(_04177_),
    .Y(_04178_));
 sky130_fd_sc_hd__o211a_1 _07751_ (.A1(\core_pipeline.memory_to_writeback_alu_data[24] ),
    .A2(net229),
    .B1(_04178_),
    .C1(net644),
    .X(_00159_));
 sky130_fd_sc_hd__a21oi_1 _07752_ (.A1(\core_pipeline.pipeline_csr.cycle[56] ),
    .A2(_04175_),
    .B1(\core_pipeline.pipeline_csr.cycle[57] ),
    .Y(_04179_));
 sky130_fd_sc_hd__and3_1 _07753_ (.A(\core_pipeline.pipeline_csr.cycle[57] ),
    .B(\core_pipeline.pipeline_csr.cycle[56] ),
    .C(_04175_),
    .X(_04180_));
 sky130_fd_sc_hd__o21ai_1 _07754_ (.A1(_04179_),
    .A2(_04180_),
    .B1(net229),
    .Y(_04181_));
 sky130_fd_sc_hd__o211a_1 _07755_ (.A1(\core_pipeline.memory_to_writeback_alu_data[25] ),
    .A2(net229),
    .B1(_04181_),
    .C1(net642),
    .X(_00160_));
 sky130_fd_sc_hd__nor2_1 _07756_ (.A(\core_pipeline.pipeline_csr.cycle[58] ),
    .B(_04180_),
    .Y(_04182_));
 sky130_fd_sc_hd__and4_1 _07757_ (.A(\core_pipeline.pipeline_csr.cycle[58] ),
    .B(\core_pipeline.pipeline_csr.cycle[57] ),
    .C(\core_pipeline.pipeline_csr.cycle[56] ),
    .D(_04175_),
    .X(_04183_));
 sky130_fd_sc_hd__o21ai_1 _07758_ (.A1(_04182_),
    .A2(_04183_),
    .B1(net227),
    .Y(_04184_));
 sky130_fd_sc_hd__o211a_1 _07759_ (.A1(\core_pipeline.memory_to_writeback_alu_data[26] ),
    .A2(net227),
    .B1(_04184_),
    .C1(net641),
    .X(_00161_));
 sky130_fd_sc_hd__nor2_1 _07760_ (.A(\core_pipeline.pipeline_csr.cycle[59] ),
    .B(_04183_),
    .Y(_04185_));
 sky130_fd_sc_hd__and2_1 _07761_ (.A(\core_pipeline.pipeline_csr.cycle[59] ),
    .B(_04183_),
    .X(_04186_));
 sky130_fd_sc_hd__o21ai_1 _07762_ (.A1(_04185_),
    .A2(_04186_),
    .B1(net227),
    .Y(_04187_));
 sky130_fd_sc_hd__o211a_1 _07763_ (.A1(\core_pipeline.memory_to_writeback_alu_data[27] ),
    .A2(net227),
    .B1(_04187_),
    .C1(net642),
    .X(_00162_));
 sky130_fd_sc_hd__nor2_1 _07764_ (.A(\core_pipeline.pipeline_csr.cycle[60] ),
    .B(_04186_),
    .Y(_04188_));
 sky130_fd_sc_hd__and3_1 _07765_ (.A(\core_pipeline.pipeline_csr.cycle[60] ),
    .B(\core_pipeline.pipeline_csr.cycle[59] ),
    .C(_04183_),
    .X(_04189_));
 sky130_fd_sc_hd__o21ai_1 _07766_ (.A1(_04188_),
    .A2(_04189_),
    .B1(net227),
    .Y(_04190_));
 sky130_fd_sc_hd__o211a_1 _07767_ (.A1(\core_pipeline.memory_to_writeback_alu_data[28] ),
    .A2(net227),
    .B1(_04190_),
    .C1(net642),
    .X(_00163_));
 sky130_fd_sc_hd__nor2_1 _07768_ (.A(\core_pipeline.pipeline_csr.cycle[61] ),
    .B(_04189_),
    .Y(_04191_));
 sky130_fd_sc_hd__and2_2 _07769_ (.A(\core_pipeline.pipeline_csr.cycle[61] ),
    .B(_04189_),
    .X(_04192_));
 sky130_fd_sc_hd__o21ai_1 _07770_ (.A1(_04191_),
    .A2(_04192_),
    .B1(net228),
    .Y(_04193_));
 sky130_fd_sc_hd__o211a_1 _07771_ (.A1(\core_pipeline.memory_to_writeback_alu_data[29] ),
    .A2(net227),
    .B1(_04193_),
    .C1(net642),
    .X(_00164_));
 sky130_fd_sc_hd__xnor2_1 _07772_ (.A(\core_pipeline.pipeline_csr.cycle[62] ),
    .B(_04192_),
    .Y(_04194_));
 sky130_fd_sc_hd__nand2_1 _07773_ (.A(net227),
    .B(_04194_),
    .Y(_04195_));
 sky130_fd_sc_hd__o211a_1 _07774_ (.A1(\core_pipeline.memory_to_writeback_alu_data[30] ),
    .A2(net227),
    .B1(_04195_),
    .C1(net641),
    .X(_00165_));
 sky130_fd_sc_hd__a21bo_1 _07775_ (.A1(\core_pipeline.pipeline_csr.cycle[62] ),
    .A2(_04192_),
    .B1_N(\core_pipeline.pipeline_csr.cycle[63] ),
    .X(_04196_));
 sky130_fd_sc_hd__nand3b_1 _07776_ (.A_N(\core_pipeline.pipeline_csr.cycle[63] ),
    .B(\core_pipeline.pipeline_csr.cycle[62] ),
    .C(_04192_),
    .Y(_04197_));
 sky130_fd_sc_hd__nand3_1 _07777_ (.A(net227),
    .B(_04196_),
    .C(_04197_),
    .Y(_04198_));
 sky130_fd_sc_hd__o211a_1 _07778_ (.A1(\core_pipeline.memory_to_writeback_alu_data[31] ),
    .A2(net227),
    .B1(_04198_),
    .C1(net641),
    .X(_00166_));
 sky130_fd_sc_hd__and3_1 _07779_ (.A(_03314_),
    .B(\core_pipeline.pipeline_csr.instret[0] ),
    .C(_03480_),
    .X(_04199_));
 sky130_fd_sc_hd__a21oi_1 _07780_ (.A1(_03314_),
    .A2(_03480_),
    .B1(\core_pipeline.pipeline_csr.instret[0] ),
    .Y(_04200_));
 sky130_fd_sc_hd__or3b_4 _07781_ (.A(_03646_),
    .B(\core_pipeline.memory_to_writeback_csr_address[0] ),
    .C_N(\core_pipeline.memory_to_writeback_csr_address[1] ),
    .X(_04201_));
 sky130_fd_sc_hd__nor2_4 _07782_ (.A(_03482_),
    .B(_04201_),
    .Y(_04202_));
 sky130_fd_sc_hd__or3_4 _07783_ (.A(_03482_),
    .B(_04021_),
    .C(_04201_),
    .X(_04203_));
 sky130_fd_sc_hd__o21ai_1 _07784_ (.A1(_04199_),
    .A2(_04200_),
    .B1(net255),
    .Y(_04204_));
 sky130_fd_sc_hd__o211a_1 _07785_ (.A1(\core_pipeline.memory_to_writeback_alu_data[0] ),
    .A2(net255),
    .B1(_04204_),
    .C1(net638),
    .X(_00167_));
 sky130_fd_sc_hd__and2_1 _07786_ (.A(\core_pipeline.pipeline_csr.instret[1] ),
    .B(\core_pipeline.pipeline_csr.instret[0] ),
    .X(_04205_));
 sky130_fd_sc_hd__and4_2 _07787_ (.A(_03314_),
    .B(\core_pipeline.memory_to_writeback_valid ),
    .C(net400),
    .D(_04205_),
    .X(_04206_));
 sky130_fd_sc_hd__o21bai_1 _07788_ (.A1(\core_pipeline.pipeline_csr.instret[1] ),
    .A2(_04199_),
    .B1_N(_04206_),
    .Y(_04207_));
 sky130_fd_sc_hd__nand2_1 _07789_ (.A(net255),
    .B(_04207_),
    .Y(_04208_));
 sky130_fd_sc_hd__o211a_1 _07790_ (.A1(\core_pipeline.memory_to_writeback_alu_data[1] ),
    .A2(net255),
    .B1(_04208_),
    .C1(net639),
    .X(_00168_));
 sky130_fd_sc_hd__xnor2_1 _07791_ (.A(\core_pipeline.pipeline_csr.instret[2] ),
    .B(_04206_),
    .Y(_04209_));
 sky130_fd_sc_hd__nand2_1 _07792_ (.A(net255),
    .B(_04209_),
    .Y(_04210_));
 sky130_fd_sc_hd__o211a_1 _07793_ (.A1(\core_pipeline.memory_to_writeback_alu_data[2] ),
    .A2(net255),
    .B1(_04210_),
    .C1(net639),
    .X(_00169_));
 sky130_fd_sc_hd__and3_2 _07794_ (.A(\core_pipeline.pipeline_csr.instret[3] ),
    .B(\core_pipeline.pipeline_csr.instret[2] ),
    .C(_04206_),
    .X(_04211_));
 sky130_fd_sc_hd__a21oi_1 _07795_ (.A1(\core_pipeline.pipeline_csr.instret[2] ),
    .A2(_04206_),
    .B1(\core_pipeline.pipeline_csr.instret[3] ),
    .Y(_04212_));
 sky130_fd_sc_hd__o21ai_1 _07796_ (.A1(_04211_),
    .A2(_04212_),
    .B1(net255),
    .Y(_04213_));
 sky130_fd_sc_hd__o211a_1 _07797_ (.A1(\core_pipeline.memory_to_writeback_alu_data[3] ),
    .A2(net255),
    .B1(_04213_),
    .C1(net639),
    .X(_00170_));
 sky130_fd_sc_hd__xnor2_1 _07798_ (.A(\core_pipeline.pipeline_csr.instret[4] ),
    .B(_04211_),
    .Y(_04214_));
 sky130_fd_sc_hd__nand2_1 _07799_ (.A(net255),
    .B(_04214_),
    .Y(_04215_));
 sky130_fd_sc_hd__o211a_1 _07800_ (.A1(\core_pipeline.memory_to_writeback_alu_data[4] ),
    .A2(net255),
    .B1(_04215_),
    .C1(net639),
    .X(_00171_));
 sky130_fd_sc_hd__and2_1 _07801_ (.A(\core_pipeline.pipeline_csr.instret[5] ),
    .B(\core_pipeline.pipeline_csr.instret[4] ),
    .X(_04216_));
 sky130_fd_sc_hd__and4_2 _07802_ (.A(\core_pipeline.pipeline_csr.instret[3] ),
    .B(\core_pipeline.pipeline_csr.instret[2] ),
    .C(_04206_),
    .D(_04216_),
    .X(_04217_));
 sky130_fd_sc_hd__a21oi_1 _07803_ (.A1(\core_pipeline.pipeline_csr.instret[4] ),
    .A2(_04211_),
    .B1(\core_pipeline.pipeline_csr.instret[5] ),
    .Y(_04218_));
 sky130_fd_sc_hd__o21ai_1 _07804_ (.A1(_04217_),
    .A2(_04218_),
    .B1(net255),
    .Y(_04219_));
 sky130_fd_sc_hd__o211a_1 _07805_ (.A1(\core_pipeline.memory_to_writeback_alu_data[5] ),
    .A2(net255),
    .B1(_04219_),
    .C1(net639),
    .X(_00172_));
 sky130_fd_sc_hd__nand2_1 _07806_ (.A(\core_pipeline.pipeline_csr.instret[6] ),
    .B(_04217_),
    .Y(_04220_));
 sky130_fd_sc_hd__or2_1 _07807_ (.A(\core_pipeline.pipeline_csr.instret[6] ),
    .B(_04217_),
    .X(_04221_));
 sky130_fd_sc_hd__a21bo_1 _07808_ (.A1(_04220_),
    .A2(_04221_),
    .B1_N(net255),
    .X(_04222_));
 sky130_fd_sc_hd__o211a_1 _07809_ (.A1(\core_pipeline.memory_to_writeback_alu_data[6] ),
    .A2(net255),
    .B1(_04222_),
    .C1(net640),
    .X(_00173_));
 sky130_fd_sc_hd__xor2_1 _07810_ (.A(\core_pipeline.pipeline_csr.instret[7] ),
    .B(_04220_),
    .X(_04223_));
 sky130_fd_sc_hd__nand2_1 _07811_ (.A(net255),
    .B(_04223_),
    .Y(_04224_));
 sky130_fd_sc_hd__o211a_1 _07812_ (.A1(\core_pipeline.memory_to_writeback_alu_data[7] ),
    .A2(net255),
    .B1(_04224_),
    .C1(net640),
    .X(_00174_));
 sky130_fd_sc_hd__and4_4 _07813_ (.A(\core_pipeline.pipeline_csr.instret[8] ),
    .B(\core_pipeline.pipeline_csr.instret[7] ),
    .C(\core_pipeline.pipeline_csr.instret[6] ),
    .D(_04217_),
    .X(_04225_));
 sky130_fd_sc_hd__a31o_1 _07814_ (.A1(\core_pipeline.pipeline_csr.instret[7] ),
    .A2(\core_pipeline.pipeline_csr.instret[6] ),
    .A3(_04217_),
    .B1(\core_pipeline.pipeline_csr.instret[8] ),
    .X(_04226_));
 sky130_fd_sc_hd__nand2b_1 _07815_ (.A_N(_04225_),
    .B(_04226_),
    .Y(_04227_));
 sky130_fd_sc_hd__nand2_1 _07816_ (.A(net255),
    .B(_04227_),
    .Y(_04228_));
 sky130_fd_sc_hd__o211a_1 _07817_ (.A1(\core_pipeline.memory_to_writeback_alu_data[8] ),
    .A2(net256),
    .B1(_04228_),
    .C1(net640),
    .X(_00175_));
 sky130_fd_sc_hd__xnor2_1 _07818_ (.A(\core_pipeline.pipeline_csr.instret[9] ),
    .B(_04225_),
    .Y(_04229_));
 sky130_fd_sc_hd__nand2_1 _07819_ (.A(net258),
    .B(_04229_),
    .Y(_04230_));
 sky130_fd_sc_hd__o211a_1 _07820_ (.A1(\core_pipeline.memory_to_writeback_alu_data[9] ),
    .A2(net258),
    .B1(_04230_),
    .C1(net636),
    .X(_00176_));
 sky130_fd_sc_hd__and3_1 _07821_ (.A(\core_pipeline.pipeline_csr.instret[10] ),
    .B(\core_pipeline.pipeline_csr.instret[9] ),
    .C(_04225_),
    .X(_04231_));
 sky130_fd_sc_hd__a21oi_1 _07822_ (.A1(\core_pipeline.pipeline_csr.instret[9] ),
    .A2(_04225_),
    .B1(\core_pipeline.pipeline_csr.instret[10] ),
    .Y(_04232_));
 sky130_fd_sc_hd__o21ai_1 _07823_ (.A1(_04231_),
    .A2(_04232_),
    .B1(net258),
    .Y(_04233_));
 sky130_fd_sc_hd__o211a_1 _07824_ (.A1(\core_pipeline.memory_to_writeback_alu_data[10] ),
    .A2(net258),
    .B1(_04233_),
    .C1(net637),
    .X(_00177_));
 sky130_fd_sc_hd__and4_4 _07825_ (.A(\core_pipeline.pipeline_csr.instret[11] ),
    .B(\core_pipeline.pipeline_csr.instret[10] ),
    .C(\core_pipeline.pipeline_csr.instret[9] ),
    .D(_04225_),
    .X(_04234_));
 sky130_fd_sc_hd__a31oi_1 _07826_ (.A1(\core_pipeline.pipeline_csr.instret[10] ),
    .A2(\core_pipeline.pipeline_csr.instret[9] ),
    .A3(_04225_),
    .B1(\core_pipeline.pipeline_csr.instret[11] ),
    .Y(_04235_));
 sky130_fd_sc_hd__o21ai_1 _07827_ (.A1(_04234_),
    .A2(_04235_),
    .B1(net258),
    .Y(_04236_));
 sky130_fd_sc_hd__o211a_1 _07828_ (.A1(\core_pipeline.memory_to_writeback_alu_data[11] ),
    .A2(net258),
    .B1(_04236_),
    .C1(net637),
    .X(_00178_));
 sky130_fd_sc_hd__xnor2_1 _07829_ (.A(\core_pipeline.pipeline_csr.instret[12] ),
    .B(_04234_),
    .Y(_04237_));
 sky130_fd_sc_hd__nand2_1 _07830_ (.A(net258),
    .B(_04237_),
    .Y(_04238_));
 sky130_fd_sc_hd__o211a_1 _07831_ (.A1(\core_pipeline.memory_to_writeback_alu_data[12] ),
    .A2(net258),
    .B1(_04238_),
    .C1(net637),
    .X(_00179_));
 sky130_fd_sc_hd__and3_1 _07832_ (.A(\core_pipeline.pipeline_csr.instret[13] ),
    .B(\core_pipeline.pipeline_csr.instret[12] ),
    .C(_04234_),
    .X(_04239_));
 sky130_fd_sc_hd__a21oi_1 _07833_ (.A1(\core_pipeline.pipeline_csr.instret[12] ),
    .A2(_04234_),
    .B1(\core_pipeline.pipeline_csr.instret[13] ),
    .Y(_04240_));
 sky130_fd_sc_hd__o21ai_1 _07834_ (.A1(_04239_),
    .A2(_04240_),
    .B1(net258),
    .Y(_04241_));
 sky130_fd_sc_hd__o211a_1 _07835_ (.A1(\core_pipeline.memory_to_writeback_alu_data[13] ),
    .A2(net258),
    .B1(_04241_),
    .C1(net637),
    .X(_00180_));
 sky130_fd_sc_hd__and4_2 _07836_ (.A(\core_pipeline.pipeline_csr.instret[14] ),
    .B(\core_pipeline.pipeline_csr.instret[13] ),
    .C(\core_pipeline.pipeline_csr.instret[12] ),
    .D(_04234_),
    .X(_04242_));
 sky130_fd_sc_hd__nor2_1 _07837_ (.A(\core_pipeline.pipeline_csr.instret[14] ),
    .B(_04239_),
    .Y(_04243_));
 sky130_fd_sc_hd__o21ai_1 _07838_ (.A1(_04242_),
    .A2(_04243_),
    .B1(net258),
    .Y(_04244_));
 sky130_fd_sc_hd__o211a_1 _07839_ (.A1(\core_pipeline.memory_to_writeback_alu_data[14] ),
    .A2(net258),
    .B1(_04244_),
    .C1(net637),
    .X(_00181_));
 sky130_fd_sc_hd__nand2_1 _07840_ (.A(\core_pipeline.pipeline_csr.instret[15] ),
    .B(_04242_),
    .Y(_04245_));
 sky130_fd_sc_hd__or2_1 _07841_ (.A(\core_pipeline.pipeline_csr.instret[15] ),
    .B(_04242_),
    .X(_04246_));
 sky130_fd_sc_hd__a21bo_1 _07842_ (.A1(_04245_),
    .A2(_04246_),
    .B1_N(net258),
    .X(_04247_));
 sky130_fd_sc_hd__o211a_1 _07843_ (.A1(\core_pipeline.memory_to_writeback_alu_data[15] ),
    .A2(net258),
    .B1(_04247_),
    .C1(net643),
    .X(_00182_));
 sky130_fd_sc_hd__xor2_1 _07844_ (.A(\core_pipeline.pipeline_csr.instret[16] ),
    .B(_04245_),
    .X(_04248_));
 sky130_fd_sc_hd__a21oi_1 _07845_ (.A1(_04203_),
    .A2(_04248_),
    .B1(net35),
    .Y(_04249_));
 sky130_fd_sc_hd__o21a_1 _07846_ (.A1(\core_pipeline.memory_to_writeback_alu_data[16] ),
    .A2(net258),
    .B1(_04249_),
    .X(_00183_));
 sky130_fd_sc_hd__and4_2 _07847_ (.A(\core_pipeline.pipeline_csr.instret[17] ),
    .B(\core_pipeline.pipeline_csr.instret[16] ),
    .C(\core_pipeline.pipeline_csr.instret[15] ),
    .D(_04242_),
    .X(_04250_));
 sky130_fd_sc_hd__a31oi_1 _07848_ (.A1(\core_pipeline.pipeline_csr.instret[16] ),
    .A2(\core_pipeline.pipeline_csr.instret[15] ),
    .A3(_04242_),
    .B1(\core_pipeline.pipeline_csr.instret[17] ),
    .Y(_04251_));
 sky130_fd_sc_hd__o21ai_1 _07849_ (.A1(_04250_),
    .A2(_04251_),
    .B1(net258),
    .Y(_04252_));
 sky130_fd_sc_hd__o211a_1 _07850_ (.A1(\core_pipeline.memory_to_writeback_alu_data[17] ),
    .A2(net257),
    .B1(_04252_),
    .C1(net643),
    .X(_00184_));
 sky130_fd_sc_hd__nand2_1 _07851_ (.A(\core_pipeline.pipeline_csr.instret[18] ),
    .B(_04250_),
    .Y(_04253_));
 sky130_fd_sc_hd__or2_1 _07852_ (.A(\core_pipeline.pipeline_csr.instret[18] ),
    .B(_04250_),
    .X(_04254_));
 sky130_fd_sc_hd__a21bo_1 _07853_ (.A1(_04253_),
    .A2(_04254_),
    .B1_N(net257),
    .X(_04255_));
 sky130_fd_sc_hd__o211a_1 _07854_ (.A1(\core_pipeline.memory_to_writeback_alu_data[18] ),
    .A2(net257),
    .B1(_04255_),
    .C1(net645),
    .X(_00185_));
 sky130_fd_sc_hd__xor2_1 _07855_ (.A(\core_pipeline.pipeline_csr.instret[19] ),
    .B(_04253_),
    .X(_04256_));
 sky130_fd_sc_hd__a21oi_1 _07856_ (.A1(net257),
    .A2(_04256_),
    .B1(net35),
    .Y(_04257_));
 sky130_fd_sc_hd__o21a_1 _07857_ (.A1(\core_pipeline.memory_to_writeback_alu_data[19] ),
    .A2(net257),
    .B1(_04257_),
    .X(_00186_));
 sky130_fd_sc_hd__and4_2 _07858_ (.A(\core_pipeline.pipeline_csr.instret[20] ),
    .B(\core_pipeline.pipeline_csr.instret[19] ),
    .C(\core_pipeline.pipeline_csr.instret[18] ),
    .D(_04250_),
    .X(_04258_));
 sky130_fd_sc_hd__a31oi_1 _07859_ (.A1(\core_pipeline.pipeline_csr.instret[19] ),
    .A2(\core_pipeline.pipeline_csr.instret[18] ),
    .A3(_04250_),
    .B1(\core_pipeline.pipeline_csr.instret[20] ),
    .Y(_04259_));
 sky130_fd_sc_hd__o21ai_1 _07860_ (.A1(_04258_),
    .A2(_04259_),
    .B1(net257),
    .Y(_04260_));
 sky130_fd_sc_hd__o211a_1 _07861_ (.A1(\core_pipeline.memory_to_writeback_alu_data[20] ),
    .A2(net257),
    .B1(_04260_),
    .C1(net644),
    .X(_00187_));
 sky130_fd_sc_hd__nand2_1 _07862_ (.A(\core_pipeline.pipeline_csr.instret[21] ),
    .B(_04258_),
    .Y(_04261_));
 sky130_fd_sc_hd__or2_1 _07863_ (.A(\core_pipeline.pipeline_csr.instret[21] ),
    .B(_04258_),
    .X(_04262_));
 sky130_fd_sc_hd__a21bo_1 _07864_ (.A1(_04261_),
    .A2(_04262_),
    .B1_N(net257),
    .X(_04263_));
 sky130_fd_sc_hd__o211a_1 _07865_ (.A1(\core_pipeline.memory_to_writeback_alu_data[21] ),
    .A2(net257),
    .B1(_04263_),
    .C1(net644),
    .X(_00188_));
 sky130_fd_sc_hd__xor2_1 _07866_ (.A(\core_pipeline.pipeline_csr.instret[22] ),
    .B(_04261_),
    .X(_04264_));
 sky130_fd_sc_hd__a21oi_1 _07867_ (.A1(net257),
    .A2(_04264_),
    .B1(net35),
    .Y(_04265_));
 sky130_fd_sc_hd__o21a_1 _07868_ (.A1(\core_pipeline.memory_to_writeback_alu_data[22] ),
    .A2(net257),
    .B1(_04265_),
    .X(_00189_));
 sky130_fd_sc_hd__and4_4 _07869_ (.A(\core_pipeline.pipeline_csr.instret[23] ),
    .B(\core_pipeline.pipeline_csr.instret[22] ),
    .C(\core_pipeline.pipeline_csr.instret[21] ),
    .D(_04258_),
    .X(_04266_));
 sky130_fd_sc_hd__a31oi_1 _07870_ (.A1(\core_pipeline.pipeline_csr.instret[22] ),
    .A2(\core_pipeline.pipeline_csr.instret[21] ),
    .A3(_04258_),
    .B1(\core_pipeline.pipeline_csr.instret[23] ),
    .Y(_04267_));
 sky130_fd_sc_hd__o21ai_1 _07871_ (.A1(_04266_),
    .A2(_04267_),
    .B1(net257),
    .Y(_04268_));
 sky130_fd_sc_hd__o211a_1 _07872_ (.A1(\core_pipeline.memory_to_writeback_alu_data[23] ),
    .A2(net257),
    .B1(_04268_),
    .C1(net644),
    .X(_00190_));
 sky130_fd_sc_hd__xnor2_1 _07873_ (.A(\core_pipeline.pipeline_csr.instret[24] ),
    .B(_04266_),
    .Y(_04269_));
 sky130_fd_sc_hd__nand2_1 _07874_ (.A(net257),
    .B(_04269_),
    .Y(_04270_));
 sky130_fd_sc_hd__o211a_1 _07875_ (.A1(\core_pipeline.memory_to_writeback_alu_data[24] ),
    .A2(net257),
    .B1(_04270_),
    .C1(net644),
    .X(_00191_));
 sky130_fd_sc_hd__and2_1 _07876_ (.A(\core_pipeline.pipeline_csr.instret[25] ),
    .B(\core_pipeline.pipeline_csr.instret[24] ),
    .X(_04271_));
 sky130_fd_sc_hd__nand2_1 _07877_ (.A(_04266_),
    .B(_04271_),
    .Y(_04272_));
 sky130_fd_sc_hd__a21o_1 _07878_ (.A1(\core_pipeline.pipeline_csr.instret[24] ),
    .A2(_04266_),
    .B1(\core_pipeline.pipeline_csr.instret[25] ),
    .X(_04273_));
 sky130_fd_sc_hd__a21bo_1 _07879_ (.A1(_04272_),
    .A2(_04273_),
    .B1_N(net257),
    .X(_04274_));
 sky130_fd_sc_hd__o211a_1 _07880_ (.A1(\core_pipeline.memory_to_writeback_alu_data[25] ),
    .A2(net257),
    .B1(_04274_),
    .C1(net644),
    .X(_00192_));
 sky130_fd_sc_hd__xor2_1 _07881_ (.A(\core_pipeline.pipeline_csr.instret[26] ),
    .B(_04272_),
    .X(_04275_));
 sky130_fd_sc_hd__nand2_1 _07882_ (.A(net256),
    .B(_04275_),
    .Y(_04276_));
 sky130_fd_sc_hd__o211a_1 _07883_ (.A1(\core_pipeline.memory_to_writeback_alu_data[26] ),
    .A2(net256),
    .B1(_04276_),
    .C1(net642),
    .X(_00193_));
 sky130_fd_sc_hd__and4_4 _07884_ (.A(\core_pipeline.pipeline_csr.instret[27] ),
    .B(\core_pipeline.pipeline_csr.instret[26] ),
    .C(_04266_),
    .D(_04271_),
    .X(_04277_));
 sky130_fd_sc_hd__a31o_1 _07885_ (.A1(\core_pipeline.pipeline_csr.instret[26] ),
    .A2(_04266_),
    .A3(_04271_),
    .B1(\core_pipeline.pipeline_csr.instret[27] ),
    .X(_04278_));
 sky130_fd_sc_hd__inv_2 _07886_ (.A(_04278_),
    .Y(_04279_));
 sky130_fd_sc_hd__o21ai_1 _07887_ (.A1(_04277_),
    .A2(_04279_),
    .B1(net256),
    .Y(_04280_));
 sky130_fd_sc_hd__o211a_1 _07888_ (.A1(\core_pipeline.memory_to_writeback_alu_data[27] ),
    .A2(net256),
    .B1(_04280_),
    .C1(net642),
    .X(_00194_));
 sky130_fd_sc_hd__xnor2_1 _07889_ (.A(\core_pipeline.pipeline_csr.instret[28] ),
    .B(_04277_),
    .Y(_04281_));
 sky130_fd_sc_hd__nand2_1 _07890_ (.A(net256),
    .B(_04281_),
    .Y(_04282_));
 sky130_fd_sc_hd__o211a_1 _07891_ (.A1(\core_pipeline.memory_to_writeback_alu_data[28] ),
    .A2(net256),
    .B1(_04282_),
    .C1(net641),
    .X(_00195_));
 sky130_fd_sc_hd__and2_1 _07892_ (.A(\core_pipeline.pipeline_csr.instret[29] ),
    .B(\core_pipeline.pipeline_csr.instret[28] ),
    .X(_04283_));
 sky130_fd_sc_hd__nand2_1 _07893_ (.A(_04277_),
    .B(_04283_),
    .Y(_04284_));
 sky130_fd_sc_hd__a21o_1 _07894_ (.A1(\core_pipeline.pipeline_csr.instret[28] ),
    .A2(_04277_),
    .B1(\core_pipeline.pipeline_csr.instret[29] ),
    .X(_04285_));
 sky130_fd_sc_hd__a21bo_1 _07895_ (.A1(_04284_),
    .A2(_04285_),
    .B1_N(net256),
    .X(_04286_));
 sky130_fd_sc_hd__o211a_1 _07896_ (.A1(\core_pipeline.memory_to_writeback_alu_data[29] ),
    .A2(net256),
    .B1(_04286_),
    .C1(net642),
    .X(_00196_));
 sky130_fd_sc_hd__xor2_1 _07897_ (.A(\core_pipeline.pipeline_csr.instret[30] ),
    .B(_04284_),
    .X(_04287_));
 sky130_fd_sc_hd__nand2_1 _07898_ (.A(net256),
    .B(_04287_),
    .Y(_04288_));
 sky130_fd_sc_hd__o211a_1 _07899_ (.A1(\core_pipeline.memory_to_writeback_alu_data[30] ),
    .A2(net256),
    .B1(_04288_),
    .C1(net641),
    .X(_00197_));
 sky130_fd_sc_hd__and4_2 _07900_ (.A(\core_pipeline.pipeline_csr.instret[31] ),
    .B(\core_pipeline.pipeline_csr.instret[30] ),
    .C(_04277_),
    .D(_04283_),
    .X(_04289_));
 sky130_fd_sc_hd__a31o_1 _07901_ (.A1(\core_pipeline.pipeline_csr.instret[30] ),
    .A2(_04277_),
    .A3(_04283_),
    .B1(\core_pipeline.pipeline_csr.instret[31] ),
    .X(_04290_));
 sky130_fd_sc_hd__nand2b_1 _07902_ (.A_N(_04289_),
    .B(_04290_),
    .Y(_04291_));
 sky130_fd_sc_hd__nand2_1 _07903_ (.A(net256),
    .B(_04291_),
    .Y(_04292_));
 sky130_fd_sc_hd__o211a_1 _07904_ (.A1(\core_pipeline.memory_to_writeback_alu_data[31] ),
    .A2(net256),
    .B1(_04292_),
    .C1(net641),
    .X(_00198_));
 sky130_fd_sc_hd__nand2_1 _07905_ (.A(\core_pipeline.pipeline_csr.instret[32] ),
    .B(_04289_),
    .Y(_04293_));
 sky130_fd_sc_hd__or2_1 _07906_ (.A(\core_pipeline.pipeline_csr.instret[32] ),
    .B(_04289_),
    .X(_04294_));
 sky130_fd_sc_hd__nand2_4 _07907_ (.A(_04111_),
    .B(_04202_),
    .Y(_04295_));
 sky130_fd_sc_hd__a21bo_1 _07908_ (.A1(_04293_),
    .A2(_04294_),
    .B1_N(net223),
    .X(_04296_));
 sky130_fd_sc_hd__o211a_1 _07909_ (.A1(\core_pipeline.memory_to_writeback_alu_data[0] ),
    .A2(net223),
    .B1(_04296_),
    .C1(net641),
    .X(_00199_));
 sky130_fd_sc_hd__xor2_1 _07910_ (.A(\core_pipeline.pipeline_csr.instret[33] ),
    .B(_04293_),
    .X(_04297_));
 sky130_fd_sc_hd__nand2_1 _07911_ (.A(net223),
    .B(_04297_),
    .Y(_04298_));
 sky130_fd_sc_hd__o211a_1 _07912_ (.A1(\core_pipeline.memory_to_writeback_alu_data[1] ),
    .A2(net223),
    .B1(_04298_),
    .C1(net641),
    .X(_00200_));
 sky130_fd_sc_hd__and4_2 _07913_ (.A(\core_pipeline.pipeline_csr.instret[34] ),
    .B(\core_pipeline.pipeline_csr.instret[33] ),
    .C(\core_pipeline.pipeline_csr.instret[32] ),
    .D(_04289_),
    .X(_04299_));
 sky130_fd_sc_hd__a31oi_1 _07914_ (.A1(\core_pipeline.pipeline_csr.instret[33] ),
    .A2(\core_pipeline.pipeline_csr.instret[32] ),
    .A3(_04289_),
    .B1(\core_pipeline.pipeline_csr.instret[34] ),
    .Y(_04300_));
 sky130_fd_sc_hd__o21ai_1 _07915_ (.A1(_04299_),
    .A2(_04300_),
    .B1(net223),
    .Y(_04301_));
 sky130_fd_sc_hd__o211a_1 _07916_ (.A1(\core_pipeline.memory_to_writeback_alu_data[2] ),
    .A2(net223),
    .B1(_04301_),
    .C1(net641),
    .X(_00201_));
 sky130_fd_sc_hd__nand2_1 _07917_ (.A(\core_pipeline.pipeline_csr.instret[35] ),
    .B(_04299_),
    .Y(_04302_));
 sky130_fd_sc_hd__or2_1 _07918_ (.A(\core_pipeline.pipeline_csr.instret[35] ),
    .B(_04299_),
    .X(_04303_));
 sky130_fd_sc_hd__a21bo_1 _07919_ (.A1(_04302_),
    .A2(_04303_),
    .B1_N(net224),
    .X(_04304_));
 sky130_fd_sc_hd__o211a_1 _07920_ (.A1(\core_pipeline.memory_to_writeback_alu_data[3] ),
    .A2(net224),
    .B1(_04304_),
    .C1(net639),
    .X(_00202_));
 sky130_fd_sc_hd__xor2_1 _07921_ (.A(\core_pipeline.pipeline_csr.instret[36] ),
    .B(_04302_),
    .X(_04305_));
 sky130_fd_sc_hd__a21oi_1 _07922_ (.A1(net224),
    .A2(_04305_),
    .B1(net35),
    .Y(_04306_));
 sky130_fd_sc_hd__o21a_1 _07923_ (.A1(\core_pipeline.memory_to_writeback_alu_data[4] ),
    .A2(net224),
    .B1(_04306_),
    .X(_00203_));
 sky130_fd_sc_hd__and4_2 _07924_ (.A(\core_pipeline.pipeline_csr.instret[37] ),
    .B(\core_pipeline.pipeline_csr.instret[36] ),
    .C(\core_pipeline.pipeline_csr.instret[35] ),
    .D(_04299_),
    .X(_04307_));
 sky130_fd_sc_hd__a31oi_1 _07925_ (.A1(\core_pipeline.pipeline_csr.instret[36] ),
    .A2(\core_pipeline.pipeline_csr.instret[35] ),
    .A3(_04299_),
    .B1(\core_pipeline.pipeline_csr.instret[37] ),
    .Y(_04308_));
 sky130_fd_sc_hd__o21ai_1 _07926_ (.A1(_04307_),
    .A2(_04308_),
    .B1(net224),
    .Y(_04309_));
 sky130_fd_sc_hd__o211a_1 _07927_ (.A1(\core_pipeline.memory_to_writeback_alu_data[5] ),
    .A2(net224),
    .B1(_04309_),
    .C1(net639),
    .X(_00204_));
 sky130_fd_sc_hd__nand2_1 _07928_ (.A(\core_pipeline.pipeline_csr.instret[38] ),
    .B(_04307_),
    .Y(_04310_));
 sky130_fd_sc_hd__or2_1 _07929_ (.A(\core_pipeline.pipeline_csr.instret[38] ),
    .B(_04307_),
    .X(_04311_));
 sky130_fd_sc_hd__a21bo_1 _07930_ (.A1(_04310_),
    .A2(_04311_),
    .B1_N(net224),
    .X(_04312_));
 sky130_fd_sc_hd__o211a_1 _07931_ (.A1(\core_pipeline.memory_to_writeback_alu_data[6] ),
    .A2(net224),
    .B1(_04312_),
    .C1(net640),
    .X(_00205_));
 sky130_fd_sc_hd__xor2_1 _07932_ (.A(\core_pipeline.pipeline_csr.instret[39] ),
    .B(_04310_),
    .X(_04313_));
 sky130_fd_sc_hd__a21oi_1 _07933_ (.A1(net224),
    .A2(_04313_),
    .B1(net35),
    .Y(_04314_));
 sky130_fd_sc_hd__o21a_1 _07934_ (.A1(\core_pipeline.memory_to_writeback_alu_data[7] ),
    .A2(net224),
    .B1(_04314_),
    .X(_00206_));
 sky130_fd_sc_hd__and4_2 _07935_ (.A(\core_pipeline.pipeline_csr.instret[40] ),
    .B(\core_pipeline.pipeline_csr.instret[39] ),
    .C(\core_pipeline.pipeline_csr.instret[38] ),
    .D(_04307_),
    .X(_04315_));
 sky130_fd_sc_hd__a31oi_1 _07936_ (.A1(\core_pipeline.pipeline_csr.instret[39] ),
    .A2(\core_pipeline.pipeline_csr.instret[38] ),
    .A3(_04307_),
    .B1(\core_pipeline.pipeline_csr.instret[40] ),
    .Y(_04316_));
 sky130_fd_sc_hd__o21ai_1 _07937_ (.A1(_04315_),
    .A2(_04316_),
    .B1(net224),
    .Y(_04317_));
 sky130_fd_sc_hd__o211a_1 _07938_ (.A1(\core_pipeline.memory_to_writeback_alu_data[8] ),
    .A2(net224),
    .B1(_04317_),
    .C1(net640),
    .X(_00207_));
 sky130_fd_sc_hd__nand2_1 _07939_ (.A(\core_pipeline.pipeline_csr.instret[41] ),
    .B(_04315_),
    .Y(_04318_));
 sky130_fd_sc_hd__or2_1 _07940_ (.A(\core_pipeline.pipeline_csr.instret[41] ),
    .B(_04315_),
    .X(_04319_));
 sky130_fd_sc_hd__a21bo_1 _07941_ (.A1(_04318_),
    .A2(_04319_),
    .B1_N(net226),
    .X(_04320_));
 sky130_fd_sc_hd__o211a_1 _07942_ (.A1(\core_pipeline.memory_to_writeback_alu_data[9] ),
    .A2(net226),
    .B1(_04320_),
    .C1(net643),
    .X(_00208_));
 sky130_fd_sc_hd__xor2_1 _07943_ (.A(\core_pipeline.pipeline_csr.instret[42] ),
    .B(_04318_),
    .X(_04321_));
 sky130_fd_sc_hd__a21oi_1 _07944_ (.A1(net226),
    .A2(_04321_),
    .B1(net35),
    .Y(_04322_));
 sky130_fd_sc_hd__o21a_1 _07945_ (.A1(\core_pipeline.memory_to_writeback_alu_data[10] ),
    .A2(net226),
    .B1(_04322_),
    .X(_00209_));
 sky130_fd_sc_hd__and4_4 _07946_ (.A(\core_pipeline.pipeline_csr.instret[43] ),
    .B(\core_pipeline.pipeline_csr.instret[42] ),
    .C(\core_pipeline.pipeline_csr.instret[41] ),
    .D(_04315_),
    .X(_04323_));
 sky130_fd_sc_hd__a31oi_1 _07947_ (.A1(\core_pipeline.pipeline_csr.instret[42] ),
    .A2(\core_pipeline.pipeline_csr.instret[41] ),
    .A3(_04315_),
    .B1(\core_pipeline.pipeline_csr.instret[43] ),
    .Y(_04324_));
 sky130_fd_sc_hd__o21ai_1 _07948_ (.A1(_04323_),
    .A2(_04324_),
    .B1(net226),
    .Y(_04325_));
 sky130_fd_sc_hd__o211a_1 _07949_ (.A1(\core_pipeline.memory_to_writeback_alu_data[11] ),
    .A2(net226),
    .B1(_04325_),
    .C1(net643),
    .X(_00210_));
 sky130_fd_sc_hd__xnor2_1 _07950_ (.A(\core_pipeline.pipeline_csr.instret[44] ),
    .B(_04323_),
    .Y(_04326_));
 sky130_fd_sc_hd__nand2_1 _07951_ (.A(net226),
    .B(_04326_),
    .Y(_04327_));
 sky130_fd_sc_hd__o211a_1 _07952_ (.A1(\core_pipeline.memory_to_writeback_alu_data[12] ),
    .A2(net226),
    .B1(_04327_),
    .C1(net646),
    .X(_00211_));
 sky130_fd_sc_hd__and2_1 _07953_ (.A(\core_pipeline.pipeline_csr.instret[45] ),
    .B(\core_pipeline.pipeline_csr.instret[44] ),
    .X(_04328_));
 sky130_fd_sc_hd__nand2_1 _07954_ (.A(_04323_),
    .B(_04328_),
    .Y(_04329_));
 sky130_fd_sc_hd__a21o_1 _07955_ (.A1(\core_pipeline.pipeline_csr.instret[44] ),
    .A2(_04323_),
    .B1(\core_pipeline.pipeline_csr.instret[45] ),
    .X(_04330_));
 sky130_fd_sc_hd__a21bo_1 _07956_ (.A1(_04329_),
    .A2(_04330_),
    .B1_N(net226),
    .X(_04331_));
 sky130_fd_sc_hd__o211a_1 _07957_ (.A1(\core_pipeline.memory_to_writeback_alu_data[13] ),
    .A2(net226),
    .B1(_04331_),
    .C1(net646),
    .X(_00212_));
 sky130_fd_sc_hd__xor2_1 _07958_ (.A(\core_pipeline.pipeline_csr.instret[46] ),
    .B(_04329_),
    .X(_04332_));
 sky130_fd_sc_hd__nand2_1 _07959_ (.A(net226),
    .B(_04332_),
    .Y(_04333_));
 sky130_fd_sc_hd__o211a_1 _07960_ (.A1(\core_pipeline.memory_to_writeback_alu_data[14] ),
    .A2(net226),
    .B1(_04333_),
    .C1(net646),
    .X(_00213_));
 sky130_fd_sc_hd__and4_2 _07961_ (.A(\core_pipeline.pipeline_csr.instret[47] ),
    .B(\core_pipeline.pipeline_csr.instret[46] ),
    .C(_04323_),
    .D(_04328_),
    .X(_04334_));
 sky130_fd_sc_hd__a31o_1 _07962_ (.A1(\core_pipeline.pipeline_csr.instret[46] ),
    .A2(_04323_),
    .A3(_04328_),
    .B1(\core_pipeline.pipeline_csr.instret[47] ),
    .X(_04335_));
 sky130_fd_sc_hd__nand2b_1 _07963_ (.A_N(_04334_),
    .B(_04335_),
    .Y(_04336_));
 sky130_fd_sc_hd__nand2_1 _07964_ (.A(net226),
    .B(_04336_),
    .Y(_04337_));
 sky130_fd_sc_hd__o211a_1 _07965_ (.A1(\core_pipeline.memory_to_writeback_alu_data[15] ),
    .A2(net226),
    .B1(_04337_),
    .C1(net646),
    .X(_00214_));
 sky130_fd_sc_hd__nand2_1 _07966_ (.A(\core_pipeline.pipeline_csr.instret[48] ),
    .B(_04334_),
    .Y(_04338_));
 sky130_fd_sc_hd__or2_1 _07967_ (.A(\core_pipeline.pipeline_csr.instret[48] ),
    .B(_04334_),
    .X(_04339_));
 sky130_fd_sc_hd__a21bo_1 _07968_ (.A1(_04338_),
    .A2(_04339_),
    .B1_N(net225),
    .X(_04340_));
 sky130_fd_sc_hd__o211a_1 _07969_ (.A1(\core_pipeline.memory_to_writeback_alu_data[16] ),
    .A2(net225),
    .B1(_04340_),
    .C1(net645),
    .X(_00215_));
 sky130_fd_sc_hd__xor2_1 _07970_ (.A(\core_pipeline.pipeline_csr.instret[49] ),
    .B(_04338_),
    .X(_04341_));
 sky130_fd_sc_hd__nand2_1 _07971_ (.A(net225),
    .B(_04341_),
    .Y(_04342_));
 sky130_fd_sc_hd__o211a_1 _07972_ (.A1(\core_pipeline.memory_to_writeback_alu_data[17] ),
    .A2(net225),
    .B1(_04342_),
    .C1(net645),
    .X(_00216_));
 sky130_fd_sc_hd__and4_2 _07973_ (.A(\core_pipeline.pipeline_csr.instret[50] ),
    .B(\core_pipeline.pipeline_csr.instret[49] ),
    .C(\core_pipeline.pipeline_csr.instret[48] ),
    .D(_04334_),
    .X(_04343_));
 sky130_fd_sc_hd__a31oi_1 _07974_ (.A1(\core_pipeline.pipeline_csr.instret[49] ),
    .A2(\core_pipeline.pipeline_csr.instret[48] ),
    .A3(_04334_),
    .B1(\core_pipeline.pipeline_csr.instret[50] ),
    .Y(_04344_));
 sky130_fd_sc_hd__o21ai_1 _07975_ (.A1(_04343_),
    .A2(_04344_),
    .B1(net225),
    .Y(_04345_));
 sky130_fd_sc_hd__o211a_1 _07976_ (.A1(\core_pipeline.memory_to_writeback_alu_data[18] ),
    .A2(net225),
    .B1(_04345_),
    .C1(net645),
    .X(_00217_));
 sky130_fd_sc_hd__nand2_1 _07977_ (.A(\core_pipeline.pipeline_csr.instret[51] ),
    .B(_04343_),
    .Y(_04346_));
 sky130_fd_sc_hd__or2_1 _07978_ (.A(\core_pipeline.pipeline_csr.instret[51] ),
    .B(_04343_),
    .X(_04347_));
 sky130_fd_sc_hd__a21bo_1 _07979_ (.A1(_04346_),
    .A2(_04347_),
    .B1_N(net225),
    .X(_04348_));
 sky130_fd_sc_hd__o211a_1 _07980_ (.A1(\core_pipeline.memory_to_writeback_alu_data[19] ),
    .A2(net225),
    .B1(_04348_),
    .C1(net645),
    .X(_00218_));
 sky130_fd_sc_hd__xor2_1 _07981_ (.A(\core_pipeline.pipeline_csr.instret[52] ),
    .B(_04346_),
    .X(_04349_));
 sky130_fd_sc_hd__a21oi_1 _07982_ (.A1(net225),
    .A2(_04349_),
    .B1(net35),
    .Y(_04350_));
 sky130_fd_sc_hd__o21a_1 _07983_ (.A1(\core_pipeline.memory_to_writeback_alu_data[20] ),
    .A2(net225),
    .B1(_04350_),
    .X(_00219_));
 sky130_fd_sc_hd__and4_2 _07984_ (.A(\core_pipeline.pipeline_csr.instret[53] ),
    .B(\core_pipeline.pipeline_csr.instret[52] ),
    .C(\core_pipeline.pipeline_csr.instret[51] ),
    .D(_04343_),
    .X(_04351_));
 sky130_fd_sc_hd__a31oi_1 _07985_ (.A1(\core_pipeline.pipeline_csr.instret[52] ),
    .A2(\core_pipeline.pipeline_csr.instret[51] ),
    .A3(_04343_),
    .B1(\core_pipeline.pipeline_csr.instret[53] ),
    .Y(_04352_));
 sky130_fd_sc_hd__o21ai_1 _07986_ (.A1(_04351_),
    .A2(_04352_),
    .B1(net226),
    .Y(_04353_));
 sky130_fd_sc_hd__o211a_1 _07987_ (.A1(\core_pipeline.memory_to_writeback_alu_data[21] ),
    .A2(net225),
    .B1(_04353_),
    .C1(net645),
    .X(_00220_));
 sky130_fd_sc_hd__nand2_1 _07988_ (.A(\core_pipeline.pipeline_csr.instret[54] ),
    .B(_04351_),
    .Y(_04354_));
 sky130_fd_sc_hd__or2_1 _07989_ (.A(\core_pipeline.pipeline_csr.instret[54] ),
    .B(_04351_),
    .X(_04355_));
 sky130_fd_sc_hd__a21bo_1 _07990_ (.A1(_04354_),
    .A2(_04355_),
    .B1_N(net225),
    .X(_04356_));
 sky130_fd_sc_hd__o211a_1 _07991_ (.A1(\core_pipeline.memory_to_writeback_alu_data[22] ),
    .A2(net225),
    .B1(_04356_),
    .C1(net644),
    .X(_00221_));
 sky130_fd_sc_hd__xor2_1 _07992_ (.A(\core_pipeline.pipeline_csr.instret[55] ),
    .B(_04354_),
    .X(_04357_));
 sky130_fd_sc_hd__a21oi_1 _07993_ (.A1(net225),
    .A2(_04357_),
    .B1(net35),
    .Y(_04358_));
 sky130_fd_sc_hd__o21a_1 _07994_ (.A1(\core_pipeline.memory_to_writeback_alu_data[23] ),
    .A2(net225),
    .B1(_04358_),
    .X(_00222_));
 sky130_fd_sc_hd__and4_2 _07995_ (.A(\core_pipeline.pipeline_csr.instret[56] ),
    .B(\core_pipeline.pipeline_csr.instret[55] ),
    .C(\core_pipeline.pipeline_csr.instret[54] ),
    .D(_04351_),
    .X(_04359_));
 sky130_fd_sc_hd__a31oi_1 _07996_ (.A1(\core_pipeline.pipeline_csr.instret[55] ),
    .A2(\core_pipeline.pipeline_csr.instret[54] ),
    .A3(_04351_),
    .B1(\core_pipeline.pipeline_csr.instret[56] ),
    .Y(_04360_));
 sky130_fd_sc_hd__o21ai_1 _07997_ (.A1(_04359_),
    .A2(_04360_),
    .B1(net225),
    .Y(_04361_));
 sky130_fd_sc_hd__o211a_1 _07998_ (.A1(\core_pipeline.memory_to_writeback_alu_data[24] ),
    .A2(net225),
    .B1(_04361_),
    .C1(net644),
    .X(_00223_));
 sky130_fd_sc_hd__nand2_1 _07999_ (.A(\core_pipeline.pipeline_csr.instret[57] ),
    .B(_04359_),
    .Y(_04362_));
 sky130_fd_sc_hd__or2_1 _08000_ (.A(\core_pipeline.pipeline_csr.instret[57] ),
    .B(_04359_),
    .X(_04363_));
 sky130_fd_sc_hd__a21bo_1 _08001_ (.A1(_04362_),
    .A2(_04363_),
    .B1_N(net223),
    .X(_04364_));
 sky130_fd_sc_hd__o211a_1 _08002_ (.A1(\core_pipeline.memory_to_writeback_alu_data[25] ),
    .A2(net223),
    .B1(_04364_),
    .C1(net644),
    .X(_00224_));
 sky130_fd_sc_hd__xor2_1 _08003_ (.A(\core_pipeline.pipeline_csr.instret[58] ),
    .B(_04362_),
    .X(_04365_));
 sky130_fd_sc_hd__a21oi_1 _08004_ (.A1(net223),
    .A2(_04365_),
    .B1(net35),
    .Y(_04366_));
 sky130_fd_sc_hd__o21a_1 _08005_ (.A1(\core_pipeline.memory_to_writeback_alu_data[26] ),
    .A2(net223),
    .B1(_04366_),
    .X(_00225_));
 sky130_fd_sc_hd__and4_2 _08006_ (.A(\core_pipeline.pipeline_csr.instret[59] ),
    .B(\core_pipeline.pipeline_csr.instret[58] ),
    .C(\core_pipeline.pipeline_csr.instret[57] ),
    .D(_04359_),
    .X(_04367_));
 sky130_fd_sc_hd__a31oi_1 _08007_ (.A1(\core_pipeline.pipeline_csr.instret[58] ),
    .A2(\core_pipeline.pipeline_csr.instret[57] ),
    .A3(_04359_),
    .B1(\core_pipeline.pipeline_csr.instret[59] ),
    .Y(_04368_));
 sky130_fd_sc_hd__o21ai_1 _08008_ (.A1(_04367_),
    .A2(_04368_),
    .B1(net224),
    .Y(_04369_));
 sky130_fd_sc_hd__o211a_1 _08009_ (.A1(\core_pipeline.memory_to_writeback_alu_data[27] ),
    .A2(net224),
    .B1(_04369_),
    .C1(net641),
    .X(_00226_));
 sky130_fd_sc_hd__xnor2_1 _08010_ (.A(\core_pipeline.pipeline_csr.instret[60] ),
    .B(_04367_),
    .Y(_04370_));
 sky130_fd_sc_hd__nand2_1 _08011_ (.A(net223),
    .B(_04370_),
    .Y(_04371_));
 sky130_fd_sc_hd__o211a_1 _08012_ (.A1(\core_pipeline.memory_to_writeback_alu_data[28] ),
    .A2(net224),
    .B1(_04371_),
    .C1(net642),
    .X(_00227_));
 sky130_fd_sc_hd__and3_1 _08013_ (.A(\core_pipeline.pipeline_csr.instret[61] ),
    .B(\core_pipeline.pipeline_csr.instret[60] ),
    .C(_04367_),
    .X(_04372_));
 sky130_fd_sc_hd__a21oi_1 _08014_ (.A1(\core_pipeline.pipeline_csr.instret[60] ),
    .A2(_04367_),
    .B1(\core_pipeline.pipeline_csr.instret[61] ),
    .Y(_04373_));
 sky130_fd_sc_hd__o21ai_1 _08015_ (.A1(_04372_),
    .A2(_04373_),
    .B1(net223),
    .Y(_04374_));
 sky130_fd_sc_hd__o211a_1 _08016_ (.A1(\core_pipeline.memory_to_writeback_alu_data[29] ),
    .A2(net223),
    .B1(_04374_),
    .C1(net641),
    .X(_00228_));
 sky130_fd_sc_hd__and4_1 _08017_ (.A(\core_pipeline.pipeline_csr.instret[62] ),
    .B(\core_pipeline.pipeline_csr.instret[61] ),
    .C(\core_pipeline.pipeline_csr.instret[60] ),
    .D(_04367_),
    .X(_04375_));
 sky130_fd_sc_hd__xnor2_1 _08018_ (.A(\core_pipeline.pipeline_csr.instret[62] ),
    .B(_04372_),
    .Y(_04376_));
 sky130_fd_sc_hd__nor2_1 _08019_ (.A(\core_pipeline.memory_to_writeback_alu_data[30] ),
    .B(net223),
    .Y(_04377_));
 sky130_fd_sc_hd__a211oi_1 _08020_ (.A1(net223),
    .A2(_04376_),
    .B1(_04377_),
    .C1(net35),
    .Y(_00229_));
 sky130_fd_sc_hd__xnor2_1 _08021_ (.A(\core_pipeline.pipeline_csr.instret[63] ),
    .B(_04375_),
    .Y(_04378_));
 sky130_fd_sc_hd__nor2_1 _08022_ (.A(\core_pipeline.memory_to_writeback_alu_data[31] ),
    .B(net223),
    .Y(_04379_));
 sky130_fd_sc_hd__a211oi_1 _08023_ (.A1(net223),
    .A2(_04378_),
    .B1(_04379_),
    .C1(net35),
    .Y(_00230_));
 sky130_fd_sc_hd__o22a_1 _08024_ (.A1(\core_pipeline.pipeline_csr.ie ),
    .A2(net400),
    .B1(_03515_),
    .B2(\core_pipeline.pipeline_csr.pie ),
    .X(_04380_));
 sky130_fd_sc_hd__or3_4 _08025_ (.A(\core_pipeline.memory_to_writeback_csr_address[0] ),
    .B(\core_pipeline.memory_to_writeback_csr_address[1] ),
    .C(_04018_),
    .X(_04381_));
 sky130_fd_sc_hd__nor2_1 _08026_ (.A(_03646_),
    .B(_04381_),
    .Y(_04382_));
 sky130_fd_sc_hd__or2_1 _08027_ (.A(_03646_),
    .B(_04381_),
    .X(_04383_));
 sky130_fd_sc_hd__or2_1 _08028_ (.A(_04380_),
    .B(_04382_),
    .X(_04384_));
 sky130_fd_sc_hd__o211a_1 _08029_ (.A1(\core_pipeline.memory_to_writeback_alu_data[7] ),
    .A2(_04383_),
    .B1(_04384_),
    .C1(net638),
    .X(_00231_));
 sky130_fd_sc_hd__nor2_8 _08030_ (.A(_03479_),
    .B(_03513_),
    .Y(_04385_));
 sky130_fd_sc_hd__a221o_1 _08031_ (.A1(\core_pipeline.pipeline_csr.ie ),
    .A2(_03514_),
    .B1(_04385_),
    .B2(\core_pipeline.pipeline_csr.pie ),
    .C1(_04382_),
    .X(_04386_));
 sky130_fd_sc_hd__o211a_1 _08032_ (.A1(\core_pipeline.memory_to_writeback_alu_data[3] ),
    .A2(_04383_),
    .B1(_04386_),
    .C1(net638),
    .X(_00232_));
 sky130_fd_sc_hd__nor2_4 _08033_ (.A(_04017_),
    .B(_04381_),
    .Y(_04387_));
 sky130_fd_sc_hd__mux2_1 _08034_ (.A0(\core_pipeline.pipeline_csr.meie ),
    .A1(\core_pipeline.memory_to_writeback_alu_data[11] ),
    .S(_04387_),
    .X(_00233_));
 sky130_fd_sc_hd__mux2_1 _08035_ (.A0(\core_pipeline.pipeline_csr.msie ),
    .A1(\core_pipeline.memory_to_writeback_alu_data[3] ),
    .S(_04387_),
    .X(_00234_));
 sky130_fd_sc_hd__nand2_1 _08036_ (.A(_03481_),
    .B(_03645_),
    .Y(_04388_));
 sky130_fd_sc_hd__or4_2 _08037_ (.A(\core_pipeline.memory_to_writeback_csr_address[0] ),
    .B(\core_pipeline.memory_to_writeback_csr_address[1] ),
    .C(_04017_),
    .D(_04388_),
    .X(_04389_));
 sky130_fd_sc_hd__mux2_1 _08038_ (.A0(\core_pipeline.memory_to_writeback_alu_data[3] ),
    .A1(\core_pipeline.pipeline_csr.msip ),
    .S(_04389_),
    .X(_00235_));
 sky130_fd_sc_hd__mux2_1 _08039_ (.A0(\core_pipeline.pipeline_csr.mtie ),
    .A1(\core_pipeline.memory_to_writeback_alu_data[7] ),
    .S(_04387_),
    .X(_00236_));
 sky130_fd_sc_hd__or3b_4 _08040_ (.A(_03648_),
    .B(\core_pipeline.memory_to_writeback_csr_address[0] ),
    .C_N(_03645_),
    .X(_04390_));
 sky130_fd_sc_hd__mux2_1 _08041_ (.A0(\core_pipeline.memory_to_writeback_alu_data[0] ),
    .A1(\core_pipeline.pipeline_csr.mscratch[0] ),
    .S(net221),
    .X(_00237_));
 sky130_fd_sc_hd__mux2_1 _08042_ (.A0(\core_pipeline.memory_to_writeback_alu_data[1] ),
    .A1(\core_pipeline.pipeline_csr.mscratch[1] ),
    .S(net221),
    .X(_00238_));
 sky130_fd_sc_hd__mux2_1 _08043_ (.A0(\core_pipeline.memory_to_writeback_alu_data[2] ),
    .A1(\core_pipeline.pipeline_csr.mscratch[2] ),
    .S(net221),
    .X(_00239_));
 sky130_fd_sc_hd__mux2_1 _08044_ (.A0(\core_pipeline.memory_to_writeback_alu_data[3] ),
    .A1(\core_pipeline.pipeline_csr.mscratch[3] ),
    .S(net221),
    .X(_00240_));
 sky130_fd_sc_hd__mux2_1 _08045_ (.A0(\core_pipeline.memory_to_writeback_alu_data[4] ),
    .A1(\core_pipeline.pipeline_csr.mscratch[4] ),
    .S(net221),
    .X(_00241_));
 sky130_fd_sc_hd__mux2_1 _08046_ (.A0(\core_pipeline.memory_to_writeback_alu_data[5] ),
    .A1(\core_pipeline.pipeline_csr.mscratch[5] ),
    .S(net221),
    .X(_00242_));
 sky130_fd_sc_hd__mux2_1 _08047_ (.A0(\core_pipeline.memory_to_writeback_alu_data[6] ),
    .A1(\core_pipeline.pipeline_csr.mscratch[6] ),
    .S(net221),
    .X(_00243_));
 sky130_fd_sc_hd__mux2_1 _08048_ (.A0(\core_pipeline.memory_to_writeback_alu_data[7] ),
    .A1(\core_pipeline.pipeline_csr.mscratch[7] ),
    .S(net221),
    .X(_00244_));
 sky130_fd_sc_hd__mux2_1 _08049_ (.A0(\core_pipeline.memory_to_writeback_alu_data[8] ),
    .A1(\core_pipeline.pipeline_csr.mscratch[8] ),
    .S(net222),
    .X(_00245_));
 sky130_fd_sc_hd__mux2_1 _08050_ (.A0(\core_pipeline.memory_to_writeback_alu_data[9] ),
    .A1(\core_pipeline.pipeline_csr.mscratch[9] ),
    .S(net222),
    .X(_00246_));
 sky130_fd_sc_hd__mux2_1 _08051_ (.A0(\core_pipeline.memory_to_writeback_alu_data[10] ),
    .A1(\core_pipeline.pipeline_csr.mscratch[10] ),
    .S(net222),
    .X(_00247_));
 sky130_fd_sc_hd__mux2_1 _08052_ (.A0(\core_pipeline.memory_to_writeback_alu_data[11] ),
    .A1(\core_pipeline.pipeline_csr.mscratch[11] ),
    .S(net221),
    .X(_00248_));
 sky130_fd_sc_hd__mux2_1 _08053_ (.A0(\core_pipeline.memory_to_writeback_alu_data[12] ),
    .A1(\core_pipeline.pipeline_csr.mscratch[12] ),
    .S(net222),
    .X(_00249_));
 sky130_fd_sc_hd__mux2_1 _08054_ (.A0(\core_pipeline.memory_to_writeback_alu_data[13] ),
    .A1(\core_pipeline.pipeline_csr.mscratch[13] ),
    .S(net222),
    .X(_00250_));
 sky130_fd_sc_hd__mux2_1 _08055_ (.A0(\core_pipeline.memory_to_writeback_alu_data[14] ),
    .A1(\core_pipeline.pipeline_csr.mscratch[14] ),
    .S(net222),
    .X(_00251_));
 sky130_fd_sc_hd__mux2_1 _08056_ (.A0(\core_pipeline.memory_to_writeback_alu_data[15] ),
    .A1(\core_pipeline.pipeline_csr.mscratch[15] ),
    .S(net222),
    .X(_00252_));
 sky130_fd_sc_hd__mux2_1 _08057_ (.A0(\core_pipeline.memory_to_writeback_alu_data[16] ),
    .A1(\core_pipeline.pipeline_csr.mscratch[16] ),
    .S(net222),
    .X(_00253_));
 sky130_fd_sc_hd__mux2_1 _08058_ (.A0(\core_pipeline.memory_to_writeback_alu_data[17] ),
    .A1(\core_pipeline.pipeline_csr.mscratch[17] ),
    .S(net222),
    .X(_00254_));
 sky130_fd_sc_hd__mux2_1 _08059_ (.A0(\core_pipeline.memory_to_writeback_alu_data[18] ),
    .A1(\core_pipeline.pipeline_csr.mscratch[18] ),
    .S(net221),
    .X(_00255_));
 sky130_fd_sc_hd__mux2_1 _08060_ (.A0(\core_pipeline.memory_to_writeback_alu_data[19] ),
    .A1(\core_pipeline.pipeline_csr.mscratch[19] ),
    .S(net221),
    .X(_00256_));
 sky130_fd_sc_hd__mux2_1 _08061_ (.A0(\core_pipeline.memory_to_writeback_alu_data[20] ),
    .A1(\core_pipeline.pipeline_csr.mscratch[20] ),
    .S(net222),
    .X(_00257_));
 sky130_fd_sc_hd__mux2_1 _08062_ (.A0(\core_pipeline.memory_to_writeback_alu_data[21] ),
    .A1(\core_pipeline.pipeline_csr.mscratch[21] ),
    .S(net222),
    .X(_00258_));
 sky130_fd_sc_hd__mux2_1 _08063_ (.A0(\core_pipeline.memory_to_writeback_alu_data[22] ),
    .A1(\core_pipeline.pipeline_csr.mscratch[22] ),
    .S(net222),
    .X(_00259_));
 sky130_fd_sc_hd__mux2_1 _08064_ (.A0(\core_pipeline.memory_to_writeback_alu_data[23] ),
    .A1(\core_pipeline.pipeline_csr.mscratch[23] ),
    .S(net222),
    .X(_00260_));
 sky130_fd_sc_hd__mux2_1 _08065_ (.A0(\core_pipeline.memory_to_writeback_alu_data[24] ),
    .A1(\core_pipeline.pipeline_csr.mscratch[24] ),
    .S(net222),
    .X(_00261_));
 sky130_fd_sc_hd__mux2_1 _08066_ (.A0(\core_pipeline.memory_to_writeback_alu_data[25] ),
    .A1(\core_pipeline.pipeline_csr.mscratch[25] ),
    .S(net222),
    .X(_00262_));
 sky130_fd_sc_hd__mux2_1 _08067_ (.A0(\core_pipeline.memory_to_writeback_alu_data[26] ),
    .A1(\core_pipeline.pipeline_csr.mscratch[26] ),
    .S(net221),
    .X(_00263_));
 sky130_fd_sc_hd__mux2_1 _08068_ (.A0(\core_pipeline.memory_to_writeback_alu_data[27] ),
    .A1(\core_pipeline.pipeline_csr.mscratch[27] ),
    .S(net221),
    .X(_00264_));
 sky130_fd_sc_hd__mux2_1 _08069_ (.A0(\core_pipeline.memory_to_writeback_alu_data[28] ),
    .A1(\core_pipeline.pipeline_csr.mscratch[28] ),
    .S(net221),
    .X(_00265_));
 sky130_fd_sc_hd__mux2_1 _08070_ (.A0(\core_pipeline.memory_to_writeback_alu_data[29] ),
    .A1(\core_pipeline.pipeline_csr.mscratch[29] ),
    .S(net221),
    .X(_00266_));
 sky130_fd_sc_hd__mux2_1 _08071_ (.A0(\core_pipeline.memory_to_writeback_alu_data[30] ),
    .A1(\core_pipeline.pipeline_csr.mscratch[30] ),
    .S(net221),
    .X(_00267_));
 sky130_fd_sc_hd__mux2_1 _08072_ (.A0(\core_pipeline.memory_to_writeback_alu_data[31] ),
    .A1(\core_pipeline.pipeline_csr.mscratch[31] ),
    .S(net221),
    .X(_00268_));
 sky130_fd_sc_hd__mux2_1 _08073_ (.A0(\core_pipeline.memory_to_writeback_ecause[0] ),
    .A1(\core_pipeline.pipeline_csr.mcause[0] ),
    .S(_03477_),
    .X(_04391_));
 sky130_fd_sc_hd__nand2_4 _08074_ (.A(_03645_),
    .B(_04202_),
    .Y(_04392_));
 sky130_fd_sc_hd__or3b_1 _08075_ (.A(_03476_),
    .B(_04391_),
    .C_N(_04392_),
    .X(_04393_));
 sky130_fd_sc_hd__o211a_1 _08076_ (.A1(\core_pipeline.memory_to_writeback_alu_data[0] ),
    .A2(_04392_),
    .B1(_04393_),
    .C1(net639),
    .X(_00269_));
 sky130_fd_sc_hd__mux2_1 _08077_ (.A0(\core_pipeline.memory_to_writeback_ecause[1] ),
    .A1(\core_pipeline.pipeline_csr.mcause[1] ),
    .S(_03477_),
    .X(_04394_));
 sky130_fd_sc_hd__or3b_1 _08078_ (.A(_04394_),
    .B(_03476_),
    .C_N(_04392_),
    .X(_04395_));
 sky130_fd_sc_hd__o211a_1 _08079_ (.A1(\core_pipeline.memory_to_writeback_alu_data[1] ),
    .A2(_04392_),
    .B1(_04395_),
    .C1(net639),
    .X(_00270_));
 sky130_fd_sc_hd__a31o_1 _08080_ (.A1(\core_pipeline.memory_to_writeback_exception ),
    .A2(\core_pipeline.memory_to_writeback_ecause[2] ),
    .A3(_03473_),
    .B1(_03472_),
    .X(_04396_));
 sky130_fd_sc_hd__a21o_1 _08081_ (.A1(_03475_),
    .A2(_04396_),
    .B1(net400),
    .X(_04397_));
 sky130_fd_sc_hd__o21ai_1 _08082_ (.A1(\core_pipeline.pipeline_csr.mcause[2] ),
    .A2(_03479_),
    .B1(_04397_),
    .Y(_04398_));
 sky130_fd_sc_hd__nand2_1 _08083_ (.A(_04392_),
    .B(_04398_),
    .Y(_04399_));
 sky130_fd_sc_hd__o211a_1 _08084_ (.A1(\core_pipeline.memory_to_writeback_alu_data[2] ),
    .A2(_04392_),
    .B1(_04399_),
    .C1(net639),
    .X(_00271_));
 sky130_fd_sc_hd__mux2_1 _08085_ (.A0(\core_pipeline.memory_to_writeback_ecause[3] ),
    .A1(\core_pipeline.pipeline_csr.mcause[3] ),
    .S(_03477_),
    .X(_04400_));
 sky130_fd_sc_hd__nand2_1 _08086_ (.A(_03474_),
    .B(_04400_),
    .Y(_04401_));
 sky130_fd_sc_hd__a31o_1 _08087_ (.A1(_03475_),
    .A2(_04392_),
    .A3(_04401_),
    .B1(net35),
    .X(_04402_));
 sky130_fd_sc_hd__o21ba_1 _08088_ (.A1(\core_pipeline.memory_to_writeback_alu_data[3] ),
    .A2(_04392_),
    .B1_N(_04402_),
    .X(_00272_));
 sky130_fd_sc_hd__a21oi_1 _08089_ (.A1(\core_pipeline.pipeline_csr.minterupt ),
    .A2(_03477_),
    .B1(_03476_),
    .Y(_04403_));
 sky130_fd_sc_hd__a21oi_1 _08090_ (.A1(_04392_),
    .A2(_04403_),
    .B1(net35),
    .Y(_04404_));
 sky130_fd_sc_hd__o21a_1 _08091_ (.A1(\core_pipeline.memory_to_writeback_alu_data[31] ),
    .A2(_04392_),
    .B1(_04404_),
    .X(_00273_));
 sky130_fd_sc_hd__mux2_1 _08092_ (.A0(net8),
    .A1(net17),
    .S(net497),
    .X(_04405_));
 sky130_fd_sc_hd__nand2b_2 _08093_ (.A_N(_04405_),
    .B(net491),
    .Y(_04406_));
 sky130_fd_sc_hd__mux2_1 _08094_ (.A0(net1),
    .A1(net31),
    .S(net494),
    .X(_04407_));
 sky130_fd_sc_hd__or2_1 _08095_ (.A(net490),
    .B(_04407_),
    .X(_04408_));
 sky130_fd_sc_hd__and2_4 _08096_ (.A(net446),
    .B(_03716_),
    .X(_04409_));
 sky130_fd_sc_hd__a32o_1 _08097_ (.A1(_04406_),
    .A2(_04408_),
    .A3(_04409_),
    .B1(net458),
    .B2(\core_pipeline.memory_to_writeback_load_data[0] ),
    .X(_00274_));
 sky130_fd_sc_hd__mux2_1 _08098_ (.A0(net9),
    .A1(net18),
    .S(net496),
    .X(_04410_));
 sky130_fd_sc_hd__mux4_1 _08099_ (.A0(net12),
    .A1(net32),
    .A2(net9),
    .A3(net18),
    .S0(net495),
    .S1(net490),
    .X(_04411_));
 sky130_fd_sc_hd__a22o_1 _08100_ (.A1(\core_pipeline.memory_to_writeback_load_data[1] ),
    .A2(net458),
    .B1(_04409_),
    .B2(_04411_),
    .X(_00275_));
 sky130_fd_sc_hd__mux2_1 _08101_ (.A0(net10),
    .A1(net19),
    .S(net497),
    .X(_04412_));
 sky130_fd_sc_hd__mux4_1 _08102_ (.A0(net23),
    .A1(net2),
    .A2(net10),
    .A3(net19),
    .S0(net494),
    .S1(net492),
    .X(_04413_));
 sky130_fd_sc_hd__a22o_1 _08103_ (.A1(\core_pipeline.memory_to_writeback_load_data[2] ),
    .A2(net458),
    .B1(_04409_),
    .B2(_04413_),
    .X(_00276_));
 sky130_fd_sc_hd__mux2_1 _08104_ (.A0(net11),
    .A1(net20),
    .S(net497),
    .X(_04414_));
 sky130_fd_sc_hd__mux4_1 _08105_ (.A0(net26),
    .A1(net3),
    .A2(net11),
    .A3(net20),
    .S0(net495),
    .S1(net490),
    .X(_04415_));
 sky130_fd_sc_hd__a22o_1 _08106_ (.A1(\core_pipeline.memory_to_writeback_load_data[3] ),
    .A2(net458),
    .B1(_04409_),
    .B2(_04415_),
    .X(_00277_));
 sky130_fd_sc_hd__mux2_1 _08107_ (.A0(net13),
    .A1(net21),
    .S(net496),
    .X(_04416_));
 sky130_fd_sc_hd__mux4_1 _08108_ (.A0(net27),
    .A1(net4),
    .A2(net13),
    .A3(net21),
    .S0(net495),
    .S1(net490),
    .X(_04417_));
 sky130_fd_sc_hd__a22o_1 _08109_ (.A1(\core_pipeline.memory_to_writeback_load_data[4] ),
    .A2(net458),
    .B1(_04409_),
    .B2(_04417_),
    .X(_00278_));
 sky130_fd_sc_hd__mux2_1 _08110_ (.A0(net14),
    .A1(net22),
    .S(net496),
    .X(_04418_));
 sky130_fd_sc_hd__mux4_1 _08111_ (.A0(net28),
    .A1(net5),
    .A2(net14),
    .A3(net22),
    .S0(net495),
    .S1(net490),
    .X(_04419_));
 sky130_fd_sc_hd__a22o_1 _08112_ (.A1(\core_pipeline.memory_to_writeback_load_data[5] ),
    .A2(net458),
    .B1(_04409_),
    .B2(_04419_),
    .X(_00279_));
 sky130_fd_sc_hd__mux2_1 _08113_ (.A0(net15),
    .A1(net24),
    .S(net497),
    .X(_04420_));
 sky130_fd_sc_hd__mux4_1 _08114_ (.A0(net29),
    .A1(net6),
    .A2(net15),
    .A3(net24),
    .S0(net495),
    .S1(net490),
    .X(_04421_));
 sky130_fd_sc_hd__a22o_1 _08115_ (.A1(\core_pipeline.memory_to_writeback_load_data[6] ),
    .A2(net458),
    .B1(_04409_),
    .B2(_04421_),
    .X(_00280_));
 sky130_fd_sc_hd__mux2_1 _08116_ (.A0(net16),
    .A1(net25),
    .S(net496),
    .X(_04422_));
 sky130_fd_sc_hd__mux4_2 _08117_ (.A0(net30),
    .A1(net7),
    .A2(net16),
    .A3(net25),
    .S0(net495),
    .S1(net490),
    .X(_04423_));
 sky130_fd_sc_hd__a22o_1 _08118_ (.A1(\core_pipeline.memory_to_writeback_load_data[7] ),
    .A2(net458),
    .B1(_04409_),
    .B2(_04423_),
    .X(_00281_));
 sky130_fd_sc_hd__a41o_4 _08119_ (.A1(_03315_),
    .A2(_03316_),
    .A3(\core_busio.mem_signed ),
    .A4(_04423_),
    .B1(net458),
    .X(_04424_));
 sky130_fd_sc_hd__mux2_1 _08120_ (.A0(net31),
    .A1(net8),
    .S(net496),
    .X(_04425_));
 sky130_fd_sc_hd__and2_4 _08121_ (.A(_03424_),
    .B(_03716_),
    .X(_04426_));
 sky130_fd_sc_hd__o21ai_1 _08122_ (.A1(net496),
    .A2(_03413_),
    .B1(net491),
    .Y(_04427_));
 sky130_fd_sc_hd__o211a_1 _08123_ (.A1(net491),
    .A2(_04425_),
    .B1(_04426_),
    .C1(_04427_),
    .X(_04428_));
 sky130_fd_sc_hd__o22a_1 _08124_ (.A1(\core_pipeline.memory_to_writeback_load_data[8] ),
    .A2(net451),
    .B1(_04424_),
    .B2(_04428_),
    .X(_00282_));
 sky130_fd_sc_hd__mux2_1 _08125_ (.A0(net32),
    .A1(net9),
    .S(net496),
    .X(_04429_));
 sky130_fd_sc_hd__o21ai_1 _08126_ (.A1(net496),
    .A2(_03414_),
    .B1(net491),
    .Y(_04430_));
 sky130_fd_sc_hd__o211a_1 _08127_ (.A1(net491),
    .A2(_04429_),
    .B1(_04430_),
    .C1(_04426_),
    .X(_04431_));
 sky130_fd_sc_hd__o22a_1 _08128_ (.A1(\core_pipeline.memory_to_writeback_load_data[9] ),
    .A2(net451),
    .B1(_04424_),
    .B2(_04431_),
    .X(_00283_));
 sky130_fd_sc_hd__mux2_1 _08129_ (.A0(net2),
    .A1(net10),
    .S(net497),
    .X(_04432_));
 sky130_fd_sc_hd__o21ai_1 _08130_ (.A1(net497),
    .A2(_03415_),
    .B1(net491),
    .Y(_04433_));
 sky130_fd_sc_hd__o211a_1 _08131_ (.A1(net490),
    .A2(_04432_),
    .B1(_04433_),
    .C1(_04426_),
    .X(_04434_));
 sky130_fd_sc_hd__o22a_1 _08132_ (.A1(\core_pipeline.memory_to_writeback_load_data[10] ),
    .A2(net451),
    .B1(_04424_),
    .B2(_04434_),
    .X(_00284_));
 sky130_fd_sc_hd__mux2_1 _08133_ (.A0(net3),
    .A1(net11),
    .S(net496),
    .X(_04435_));
 sky130_fd_sc_hd__o21ai_1 _08134_ (.A1(net496),
    .A2(_03416_),
    .B1(net490),
    .Y(_04436_));
 sky130_fd_sc_hd__o211a_1 _08135_ (.A1(net491),
    .A2(_04435_),
    .B1(_04436_),
    .C1(_04426_),
    .X(_04437_));
 sky130_fd_sc_hd__o22a_1 _08136_ (.A1(\core_pipeline.memory_to_writeback_load_data[11] ),
    .A2(net446),
    .B1(_04424_),
    .B2(_04437_),
    .X(_00285_));
 sky130_fd_sc_hd__mux2_1 _08137_ (.A0(net4),
    .A1(net13),
    .S(net495),
    .X(_04438_));
 sky130_fd_sc_hd__o21ai_1 _08138_ (.A1(net496),
    .A2(_03417_),
    .B1(net490),
    .Y(_04439_));
 sky130_fd_sc_hd__o211a_1 _08139_ (.A1(net490),
    .A2(_04438_),
    .B1(_04439_),
    .C1(_04426_),
    .X(_04440_));
 sky130_fd_sc_hd__o22a_1 _08140_ (.A1(\core_pipeline.memory_to_writeback_load_data[12] ),
    .A2(net451),
    .B1(_04424_),
    .B2(_04440_),
    .X(_00286_));
 sky130_fd_sc_hd__mux2_1 _08141_ (.A0(net5),
    .A1(net14),
    .S(net495),
    .X(_04441_));
 sky130_fd_sc_hd__o21ai_1 _08142_ (.A1(net496),
    .A2(_03418_),
    .B1(net491),
    .Y(_04442_));
 sky130_fd_sc_hd__o211a_1 _08143_ (.A1(net491),
    .A2(_04441_),
    .B1(_04442_),
    .C1(_04426_),
    .X(_04443_));
 sky130_fd_sc_hd__o22a_1 _08144_ (.A1(\core_pipeline.memory_to_writeback_load_data[13] ),
    .A2(net447),
    .B1(_04424_),
    .B2(_04443_),
    .X(_00287_));
 sky130_fd_sc_hd__mux2_1 _08145_ (.A0(net6),
    .A1(net15),
    .S(net497),
    .X(_04444_));
 sky130_fd_sc_hd__o21ai_1 _08146_ (.A1(net497),
    .A2(_03419_),
    .B1(net490),
    .Y(_04445_));
 sky130_fd_sc_hd__o211a_1 _08147_ (.A1(net491),
    .A2(_04444_),
    .B1(_04445_),
    .C1(_04426_),
    .X(_04446_));
 sky130_fd_sc_hd__o22a_1 _08148_ (.A1(\core_pipeline.memory_to_writeback_load_data[14] ),
    .A2(net451),
    .B1(_04424_),
    .B2(_04446_),
    .X(_00288_));
 sky130_fd_sc_hd__and2b_1 _08149_ (.A_N(net495),
    .B(net25),
    .X(_04447_));
 sky130_fd_sc_hd__mux2_1 _08150_ (.A0(net7),
    .A1(net16),
    .S(net495),
    .X(_04448_));
 sky130_fd_sc_hd__mux2_2 _08151_ (.A0(_04448_),
    .A1(_04447_),
    .S(net490),
    .X(_04449_));
 sky130_fd_sc_hd__a21o_1 _08152_ (.A1(_04426_),
    .A2(_04449_),
    .B1(_04424_),
    .X(_04450_));
 sky130_fd_sc_hd__o21a_1 _08153_ (.A1(\core_pipeline.memory_to_writeback_load_data[15] ),
    .A2(net450),
    .B1(_04450_),
    .X(_00289_));
 sky130_fd_sc_hd__and2_1 _08154_ (.A(_03425_),
    .B(_04405_),
    .X(_04451_));
 sky130_fd_sc_hd__a41o_4 _08155_ (.A1(_03315_),
    .A2(\core_busio.mem_size[0] ),
    .A3(\core_busio.mem_signed ),
    .A4(_04449_),
    .B1(_04424_),
    .X(_04452_));
 sky130_fd_sc_hd__o22a_1 _08156_ (.A1(\core_pipeline.memory_to_writeback_load_data[16] ),
    .A2(net451),
    .B1(_04451_),
    .B2(_04452_),
    .X(_00290_));
 sky130_fd_sc_hd__and2_1 _08157_ (.A(_03425_),
    .B(_04410_),
    .X(_04453_));
 sky130_fd_sc_hd__o22a_1 _08158_ (.A1(\core_pipeline.memory_to_writeback_load_data[17] ),
    .A2(net452),
    .B1(_04452_),
    .B2(_04453_),
    .X(_00291_));
 sky130_fd_sc_hd__and2_1 _08159_ (.A(_03425_),
    .B(_04412_),
    .X(_04454_));
 sky130_fd_sc_hd__o22a_1 _08160_ (.A1(\core_pipeline.memory_to_writeback_load_data[18] ),
    .A2(net451),
    .B1(_04452_),
    .B2(_04454_),
    .X(_00292_));
 sky130_fd_sc_hd__and2_1 _08161_ (.A(_03425_),
    .B(_04414_),
    .X(_04455_));
 sky130_fd_sc_hd__o22a_1 _08162_ (.A1(\core_pipeline.memory_to_writeback_load_data[19] ),
    .A2(net451),
    .B1(_04452_),
    .B2(_04455_),
    .X(_00293_));
 sky130_fd_sc_hd__and2_1 _08163_ (.A(_03425_),
    .B(_04416_),
    .X(_04456_));
 sky130_fd_sc_hd__o22a_1 _08164_ (.A1(\core_pipeline.memory_to_writeback_load_data[20] ),
    .A2(net452),
    .B1(_04452_),
    .B2(_04456_),
    .X(_00294_));
 sky130_fd_sc_hd__and2_1 _08165_ (.A(_03425_),
    .B(_04418_),
    .X(_04457_));
 sky130_fd_sc_hd__o22a_1 _08166_ (.A1(\core_pipeline.memory_to_writeback_load_data[21] ),
    .A2(net452),
    .B1(_04452_),
    .B2(_04457_),
    .X(_00295_));
 sky130_fd_sc_hd__and2_1 _08167_ (.A(_03425_),
    .B(_04420_),
    .X(_04458_));
 sky130_fd_sc_hd__o22a_1 _08168_ (.A1(\core_pipeline.memory_to_writeback_load_data[22] ),
    .A2(net452),
    .B1(_04452_),
    .B2(_04458_),
    .X(_00296_));
 sky130_fd_sc_hd__and2_1 _08169_ (.A(_03425_),
    .B(_04422_),
    .X(_04459_));
 sky130_fd_sc_hd__o22a_1 _08170_ (.A1(\core_pipeline.memory_to_writeback_load_data[23] ),
    .A2(net451),
    .B1(_04452_),
    .B2(_04459_),
    .X(_00297_));
 sky130_fd_sc_hd__and3b_1 _08171_ (.A_N(net496),
    .B(net17),
    .C(_03425_),
    .X(_04460_));
 sky130_fd_sc_hd__o22a_1 _08172_ (.A1(\core_pipeline.memory_to_writeback_load_data[24] ),
    .A2(net451),
    .B1(_04452_),
    .B2(_04460_),
    .X(_00298_));
 sky130_fd_sc_hd__and3b_1 _08173_ (.A_N(net496),
    .B(net18),
    .C(_03425_),
    .X(_04461_));
 sky130_fd_sc_hd__o22a_1 _08174_ (.A1(\core_pipeline.memory_to_writeback_load_data[25] ),
    .A2(net451),
    .B1(_04452_),
    .B2(_04461_),
    .X(_00299_));
 sky130_fd_sc_hd__and3b_1 _08175_ (.A_N(net496),
    .B(net19),
    .C(_03425_),
    .X(_04462_));
 sky130_fd_sc_hd__o22a_1 _08176_ (.A1(\core_pipeline.memory_to_writeback_load_data[26] ),
    .A2(net451),
    .B1(_04452_),
    .B2(_04462_),
    .X(_00300_));
 sky130_fd_sc_hd__and3b_1 _08177_ (.A_N(net496),
    .B(net20),
    .C(_03425_),
    .X(_04463_));
 sky130_fd_sc_hd__o22a_1 _08178_ (.A1(\core_pipeline.memory_to_writeback_load_data[27] ),
    .A2(net452),
    .B1(_04452_),
    .B2(_04463_),
    .X(_00301_));
 sky130_fd_sc_hd__and3b_1 _08179_ (.A_N(net496),
    .B(net21),
    .C(_03425_),
    .X(_04464_));
 sky130_fd_sc_hd__o22a_1 _08180_ (.A1(\core_pipeline.memory_to_writeback_load_data[28] ),
    .A2(net446),
    .B1(_04452_),
    .B2(_04464_),
    .X(_00302_));
 sky130_fd_sc_hd__and3b_1 _08181_ (.A_N(net495),
    .B(net22),
    .C(_03425_),
    .X(_04465_));
 sky130_fd_sc_hd__o22a_1 _08182_ (.A1(\core_pipeline.memory_to_writeback_load_data[29] ),
    .A2(net446),
    .B1(_04452_),
    .B2(_04465_),
    .X(_00303_));
 sky130_fd_sc_hd__and3b_1 _08183_ (.A_N(net495),
    .B(net24),
    .C(_03425_),
    .X(_04466_));
 sky130_fd_sc_hd__o22a_1 _08184_ (.A1(\core_pipeline.memory_to_writeback_load_data[30] ),
    .A2(net446),
    .B1(_04452_),
    .B2(_04466_),
    .X(_00304_));
 sky130_fd_sc_hd__and2_1 _08185_ (.A(_03425_),
    .B(_04447_),
    .X(_04467_));
 sky130_fd_sc_hd__o22a_1 _08186_ (.A1(\core_pipeline.memory_to_writeback_load_data[31] ),
    .A2(net447),
    .B1(_04452_),
    .B2(_04467_),
    .X(_00305_));
 sky130_fd_sc_hd__nand2_4 _08187_ (.A(\core_pipeline.memory_to_writeback_rd_address[3] ),
    .B(_03480_),
    .Y(_04468_));
 sky130_fd_sc_hd__nand4_4 _08188_ (.A(\core_pipeline.memory_to_writeback_rd_address[2] ),
    .B(\core_pipeline.memory_to_writeback_rd_address[3] ),
    .C(\core_pipeline.memory_to_writeback_rd_address[4] ),
    .D(_03480_),
    .Y(_04469_));
 sky130_fd_sc_hd__nor2_8 _08189_ (.A(_03915_),
    .B(_04469_),
    .Y(_04470_));
 sky130_fd_sc_hd__mux2_1 _08190_ (.A0(\core_pipeline.pipeline_registers.registers[31][0] ),
    .A1(net349),
    .S(net253),
    .X(_00306_));
 sky130_fd_sc_hd__mux2_1 _08191_ (.A0(\core_pipeline.pipeline_registers.registers[31][1] ),
    .A1(net346),
    .S(net254),
    .X(_00307_));
 sky130_fd_sc_hd__mux2_1 _08192_ (.A0(\core_pipeline.pipeline_registers.registers[31][2] ),
    .A1(net344),
    .S(net254),
    .X(_00308_));
 sky130_fd_sc_hd__mux2_1 _08193_ (.A0(\core_pipeline.pipeline_registers.registers[31][3] ),
    .A1(net342),
    .S(net253),
    .X(_00309_));
 sky130_fd_sc_hd__mux2_1 _08194_ (.A0(\core_pipeline.pipeline_registers.registers[31][4] ),
    .A1(net341),
    .S(net253),
    .X(_00310_));
 sky130_fd_sc_hd__mux2_1 _08195_ (.A0(\core_pipeline.pipeline_registers.registers[31][5] ),
    .A1(net337),
    .S(net254),
    .X(_00311_));
 sky130_fd_sc_hd__mux2_1 _08196_ (.A0(\core_pipeline.pipeline_registers.registers[31][6] ),
    .A1(net335),
    .S(net254),
    .X(_00312_));
 sky130_fd_sc_hd__mux2_1 _08197_ (.A0(\core_pipeline.pipeline_registers.registers[31][7] ),
    .A1(net333),
    .S(net253),
    .X(_00313_));
 sky130_fd_sc_hd__mux2_1 _08198_ (.A0(\core_pipeline.pipeline_registers.registers[31][8] ),
    .A1(net332),
    .S(net253),
    .X(_00314_));
 sky130_fd_sc_hd__mux2_1 _08199_ (.A0(\core_pipeline.pipeline_registers.registers[31][9] ),
    .A1(net330),
    .S(net253),
    .X(_00315_));
 sky130_fd_sc_hd__mux2_1 _08200_ (.A0(\core_pipeline.pipeline_registers.registers[31][10] ),
    .A1(net328),
    .S(net253),
    .X(_00316_));
 sky130_fd_sc_hd__mux2_1 _08201_ (.A0(\core_pipeline.pipeline_registers.registers[31][11] ),
    .A1(net326),
    .S(net253),
    .X(_00317_));
 sky130_fd_sc_hd__mux2_1 _08202_ (.A0(\core_pipeline.pipeline_registers.registers[31][12] ),
    .A1(net324),
    .S(net253),
    .X(_00318_));
 sky130_fd_sc_hd__mux2_1 _08203_ (.A0(\core_pipeline.pipeline_registers.registers[31][13] ),
    .A1(net322),
    .S(net253),
    .X(_00319_));
 sky130_fd_sc_hd__mux2_1 _08204_ (.A0(\core_pipeline.pipeline_registers.registers[31][14] ),
    .A1(net319),
    .S(net253),
    .X(_00320_));
 sky130_fd_sc_hd__mux2_1 _08205_ (.A0(\core_pipeline.pipeline_registers.registers[31][15] ),
    .A1(net318),
    .S(net253),
    .X(_00321_));
 sky130_fd_sc_hd__mux2_1 _08206_ (.A0(\core_pipeline.pipeline_registers.registers[31][16] ),
    .A1(net316),
    .S(net253),
    .X(_00322_));
 sky130_fd_sc_hd__mux2_1 _08207_ (.A0(\core_pipeline.pipeline_registers.registers[31][17] ),
    .A1(net312),
    .S(net254),
    .X(_00323_));
 sky130_fd_sc_hd__mux2_1 _08208_ (.A0(\core_pipeline.pipeline_registers.registers[31][18] ),
    .A1(net310),
    .S(net254),
    .X(_00324_));
 sky130_fd_sc_hd__mux2_1 _08209_ (.A0(\core_pipeline.pipeline_registers.registers[31][19] ),
    .A1(net309),
    .S(net254),
    .X(_00325_));
 sky130_fd_sc_hd__mux2_1 _08210_ (.A0(\core_pipeline.pipeline_registers.registers[31][20] ),
    .A1(net305),
    .S(net254),
    .X(_00326_));
 sky130_fd_sc_hd__mux2_1 _08211_ (.A0(\core_pipeline.pipeline_registers.registers[31][21] ),
    .A1(net303),
    .S(net254),
    .X(_00327_));
 sky130_fd_sc_hd__mux2_1 _08212_ (.A0(\core_pipeline.pipeline_registers.registers[31][22] ),
    .A1(net301),
    .S(net253),
    .X(_00328_));
 sky130_fd_sc_hd__mux2_1 _08213_ (.A0(\core_pipeline.pipeline_registers.registers[31][23] ),
    .A1(net299),
    .S(net254),
    .X(_00329_));
 sky130_fd_sc_hd__mux2_1 _08214_ (.A0(\core_pipeline.pipeline_registers.registers[31][24] ),
    .A1(net297),
    .S(net253),
    .X(_00330_));
 sky130_fd_sc_hd__mux2_1 _08215_ (.A0(\core_pipeline.pipeline_registers.registers[31][25] ),
    .A1(net296),
    .S(net253),
    .X(_00331_));
 sky130_fd_sc_hd__mux2_1 _08216_ (.A0(\core_pipeline.pipeline_registers.registers[31][26] ),
    .A1(net294),
    .S(net253),
    .X(_00332_));
 sky130_fd_sc_hd__mux2_1 _08217_ (.A0(\core_pipeline.pipeline_registers.registers[31][27] ),
    .A1(net291),
    .S(net254),
    .X(_00333_));
 sky130_fd_sc_hd__mux2_1 _08218_ (.A0(\core_pipeline.pipeline_registers.registers[31][28] ),
    .A1(net289),
    .S(net254),
    .X(_00334_));
 sky130_fd_sc_hd__mux2_1 _08219_ (.A0(\core_pipeline.pipeline_registers.registers[31][29] ),
    .A1(net286),
    .S(net254),
    .X(_00335_));
 sky130_fd_sc_hd__mux2_1 _08220_ (.A0(\core_pipeline.pipeline_registers.registers[31][30] ),
    .A1(net284),
    .S(net254),
    .X(_00336_));
 sky130_fd_sc_hd__mux2_1 _08221_ (.A0(\core_pipeline.pipeline_registers.registers[31][31] ),
    .A1(net282),
    .S(net254),
    .X(_00337_));
 sky130_fd_sc_hd__nor3b_4 _08222_ (.A(\core_pipeline.decode_to_execute_alu_function[2] ),
    .B(\core_pipeline.decode_to_execute_alu_function[1] ),
    .C_N(\core_pipeline.decode_to_execute_alu_function[0] ),
    .Y(_04471_));
 sky130_fd_sc_hd__or3b_4 _08223_ (.A(\core_pipeline.decode_to_execute_alu_function[2] ),
    .B(\core_pipeline.decode_to_execute_alu_function[1] ),
    .C_N(\core_pipeline.decode_to_execute_alu_function[0] ),
    .X(_04472_));
 sky130_fd_sc_hd__and2_1 _08224_ (.A(\core_pipeline.pipeline_execute.ex_alu.result_sll[0] ),
    .B(net435),
    .X(_04473_));
 sky130_fd_sc_hd__nor2_8 _08225_ (.A(net503),
    .B(net501),
    .Y(_04474_));
 sky130_fd_sc_hd__a22o_2 _08226_ (.A1(net501),
    .A2(\core_pipeline.decode_to_execute_csr_data[3] ),
    .B1(\core_pipeline.decode_to_execute_imm_data[3] ),
    .B2(net503),
    .X(_04475_));
 sky130_fd_sc_hd__a21oi_4 _08227_ (.A1(_03886_),
    .A2(net434),
    .B1(_04475_),
    .Y(_04476_));
 sky130_fd_sc_hd__a21o_2 _08228_ (.A1(_03886_),
    .A2(net434),
    .B1(_04475_),
    .X(_04477_));
 sky130_fd_sc_hd__a22o_2 _08229_ (.A1(net501),
    .A2(\core_pipeline.decode_to_execute_csr_data[4] ),
    .B1(\core_pipeline.decode_to_execute_imm_data[4] ),
    .B2(net503),
    .X(_04478_));
 sky130_fd_sc_hd__a21oi_4 _08230_ (.A1(_03869_),
    .A2(net434),
    .B1(_04478_),
    .Y(_04479_));
 sky130_fd_sc_hd__a21o_4 _08231_ (.A1(_03869_),
    .A2(net434),
    .B1(_04478_),
    .X(_04480_));
 sky130_fd_sc_hd__nor2_2 _08232_ (.A(net435),
    .B(net389),
    .Y(_04481_));
 sky130_fd_sc_hd__nand2_1 _08233_ (.A(net437),
    .B(net392),
    .Y(_04482_));
 sky130_fd_sc_hd__a22o_4 _08234_ (.A1(net501),
    .A2(\core_pipeline.decode_to_execute_csr_data[2] ),
    .B1(\core_pipeline.decode_to_execute_imm_data[2] ),
    .B2(net503),
    .X(_04483_));
 sky130_fd_sc_hd__a21oi_4 _08235_ (.A1(_03881_),
    .A2(net434),
    .B1(_04483_),
    .Y(_04484_));
 sky130_fd_sc_hd__a21o_4 _08236_ (.A1(_03881_),
    .A2(net434),
    .B1(_04483_),
    .X(_04485_));
 sky130_fd_sc_hd__and2_2 _08237_ (.A(net503),
    .B(\core_pipeline.decode_to_execute_imm_data[1] ),
    .X(_04486_));
 sky130_fd_sc_hd__a221oi_4 _08238_ (.A1(net501),
    .A2(\core_pipeline.decode_to_execute_csr_data[1] ),
    .B1(_03873_),
    .B2(net434),
    .C1(_04486_),
    .Y(_04487_));
 sky130_fd_sc_hd__a221o_4 _08239_ (.A1(net501),
    .A2(\core_pipeline.decode_to_execute_csr_data[1] ),
    .B1(_03873_),
    .B2(net434),
    .C1(_04486_),
    .X(_04488_));
 sky130_fd_sc_hd__and2_2 _08240_ (.A(net501),
    .B(\core_pipeline.decode_to_execute_csr_data[0] ),
    .X(_04489_));
 sky130_fd_sc_hd__a221oi_4 _08241_ (.A1(\core_pipeline.decode_to_execute_imm_data[0] ),
    .A2(net503),
    .B1(_03877_),
    .B2(net434),
    .C1(_04489_),
    .Y(_04490_));
 sky130_fd_sc_hd__a221o_2 _08242_ (.A1(\core_pipeline.decode_to_execute_imm_data[0] ),
    .A2(net503),
    .B1(_03877_),
    .B2(net434),
    .C1(_04489_),
    .X(_04491_));
 sky130_fd_sc_hd__nor2_2 _08243_ (.A(net379),
    .B(net374),
    .Y(_04492_));
 sky130_fd_sc_hd__nor2_2 _08244_ (.A(net627),
    .B(net629),
    .Y(_04493_));
 sky130_fd_sc_hd__a22o_1 _08245_ (.A1(net630),
    .A2(\core_pipeline.decode_to_execute_next_pc[0] ),
    .B1(\core_pipeline.decode_to_execute_imm_data[0] ),
    .B2(net628),
    .X(_04494_));
 sky130_fd_sc_hd__a21o_4 _08246_ (.A1(_03879_),
    .A2(net432),
    .B1(_04494_),
    .X(_04495_));
 sky130_fd_sc_hd__nand2_2 _08247_ (.A(net377),
    .B(_04495_),
    .Y(_04496_));
 sky130_fd_sc_hd__nor2_2 _08248_ (.A(net379),
    .B(_04496_),
    .Y(_04497_));
 sky130_fd_sc_hd__nor2_8 _08249_ (.A(net395),
    .B(net384),
    .Y(_04498_));
 sky130_fd_sc_hd__nand2_8 _08250_ (.A(net399),
    .B(net388),
    .Y(_04499_));
 sky130_fd_sc_hd__and4_4 _08251_ (.A(net398),
    .B(net387),
    .C(net382),
    .D(net376),
    .X(_04500_));
 sky130_fd_sc_hd__a31o_1 _08252_ (.A1(net280),
    .A2(_04495_),
    .A3(_04500_),
    .B1(_04473_),
    .X(_00338_));
 sky130_fd_sc_hd__a22o_1 _08253_ (.A1(net628),
    .A2(\core_pipeline.decode_to_execute_imm_data[1] ),
    .B1(\core_pipeline.decode_to_execute_next_pc[1] ),
    .B2(net630),
    .X(_04501_));
 sky130_fd_sc_hd__a21o_4 _08254_ (.A1(_03875_),
    .A2(net432),
    .B1(_04501_),
    .X(_04502_));
 sky130_fd_sc_hd__nor2_1 _08255_ (.A(net377),
    .B(_04495_),
    .Y(_04503_));
 sky130_fd_sc_hd__or2_2 _08256_ (.A(net377),
    .B(_04495_),
    .X(_04504_));
 sky130_fd_sc_hd__o21ai_4 _08257_ (.A1(net374),
    .A2(_04502_),
    .B1(_04504_),
    .Y(_04505_));
 sky130_fd_sc_hd__inv_2 _08258_ (.A(_04505_),
    .Y(_04506_));
 sky130_fd_sc_hd__nor2_4 _08259_ (.A(net379),
    .B(_04505_),
    .Y(_04507_));
 sky130_fd_sc_hd__a32o_1 _08260_ (.A1(net280),
    .A2(_04498_),
    .A3(_04507_),
    .B1(net435),
    .B2(\core_pipeline.pipeline_execute.ex_alu.result_sll[1] ),
    .X(_00339_));
 sky130_fd_sc_hd__and2_2 _08261_ (.A(net379),
    .B(_04496_),
    .X(_04508_));
 sky130_fd_sc_hd__nand2_1 _08262_ (.A(net374),
    .B(_04502_),
    .Y(_04509_));
 sky130_fd_sc_hd__a22o_1 _08263_ (.A1(net628),
    .A2(\core_pipeline.decode_to_execute_imm_data[2] ),
    .B1(\core_pipeline.decode_to_execute_pc[2] ),
    .B2(net630),
    .X(_04510_));
 sky130_fd_sc_hd__a21oi_4 _08264_ (.A1(_03882_),
    .A2(net432),
    .B1(_04510_),
    .Y(_04511_));
 sky130_fd_sc_hd__o21a_2 _08265_ (.A1(net374),
    .A2(_04511_),
    .B1(_04509_),
    .X(_04512_));
 sky130_fd_sc_hd__inv_2 _08266_ (.A(_04512_),
    .Y(_04513_));
 sky130_fd_sc_hd__a21oi_4 _08267_ (.A1(net380),
    .A2(_04512_),
    .B1(_04508_),
    .Y(_04514_));
 sky130_fd_sc_hd__a32o_1 _08268_ (.A1(net280),
    .A2(_04498_),
    .A3(_04514_),
    .B1(net435),
    .B2(\core_pipeline.pipeline_execute.ex_alu.result_sll[2] ),
    .X(_00340_));
 sky130_fd_sc_hd__nor2_1 _08269_ (.A(net377),
    .B(_04511_),
    .Y(_04515_));
 sky130_fd_sc_hd__a22o_1 _08270_ (.A1(net628),
    .A2(\core_pipeline.decode_to_execute_imm_data[3] ),
    .B1(\core_pipeline.decode_to_execute_pc[3] ),
    .B2(net630),
    .X(_04516_));
 sky130_fd_sc_hd__a21oi_4 _08271_ (.A1(_03887_),
    .A2(net432),
    .B1(_04516_),
    .Y(_04517_));
 sky130_fd_sc_hd__nor2_1 _08272_ (.A(net374),
    .B(_04517_),
    .Y(_04518_));
 sky130_fd_sc_hd__or2_1 _08273_ (.A(_04515_),
    .B(_04518_),
    .X(_04519_));
 sky130_fd_sc_hd__mux2_4 _08274_ (.A0(_04506_),
    .A1(_04519_),
    .S(net380),
    .X(_04520_));
 sky130_fd_sc_hd__a32o_1 _08275_ (.A1(net280),
    .A2(_04498_),
    .A3(_04520_),
    .B1(net435),
    .B2(\core_pipeline.pipeline_execute.ex_alu.result_sll[3] ),
    .X(_00341_));
 sky130_fd_sc_hd__a22o_1 _08276_ (.A1(net628),
    .A2(\core_pipeline.decode_to_execute_imm_data[4] ),
    .B1(\core_pipeline.decode_to_execute_pc[4] ),
    .B2(net630),
    .X(_04521_));
 sky130_fd_sc_hd__a21o_4 _08277_ (.A1(_03870_),
    .A2(net432),
    .B1(_04521_),
    .X(_04522_));
 sky130_fd_sc_hd__inv_2 _08278_ (.A(_04522_),
    .Y(_04523_));
 sky130_fd_sc_hd__nor2_1 _08279_ (.A(net374),
    .B(_04523_),
    .Y(_04524_));
 sky130_fd_sc_hd__o21bai_2 _08280_ (.A1(net377),
    .A2(_04517_),
    .B1_N(_04524_),
    .Y(_04525_));
 sky130_fd_sc_hd__mux2_1 _08281_ (.A0(_04513_),
    .A1(_04525_),
    .S(net380),
    .X(_04526_));
 sky130_fd_sc_hd__mux2_2 _08282_ (.A0(_04497_),
    .A1(_04526_),
    .S(net388),
    .X(_04527_));
 sky130_fd_sc_hd__a32o_1 _08283_ (.A1(net399),
    .A2(net280),
    .A3(_04527_),
    .B1(net435),
    .B2(\core_pipeline.pipeline_execute.ex_alu.result_sll[4] ),
    .X(_00342_));
 sky130_fd_sc_hd__nor2_1 _08284_ (.A(net377),
    .B(_04523_),
    .Y(_04528_));
 sky130_fd_sc_hd__a22o_1 _08285_ (.A1(net628),
    .A2(\core_pipeline.decode_to_execute_imm_data[5] ),
    .B1(\core_pipeline.decode_to_execute_pc[5] ),
    .B2(net630),
    .X(_04529_));
 sky130_fd_sc_hd__a21o_4 _08286_ (.A1(_03867_),
    .A2(net432),
    .B1(_04529_),
    .X(_04530_));
 sky130_fd_sc_hd__and2_1 _08287_ (.A(net377),
    .B(_04530_),
    .X(_04531_));
 sky130_fd_sc_hd__or2_1 _08288_ (.A(_04528_),
    .B(_04531_),
    .X(_04532_));
 sky130_fd_sc_hd__mux2_1 _08289_ (.A0(_04519_),
    .A1(_04532_),
    .S(net380),
    .X(_04533_));
 sky130_fd_sc_hd__mux2_2 _08290_ (.A0(_04507_),
    .A1(_04533_),
    .S(net388),
    .X(_04534_));
 sky130_fd_sc_hd__a32o_1 _08291_ (.A1(net399),
    .A2(net280),
    .A3(_04534_),
    .B1(net435),
    .B2(\core_pipeline.pipeline_execute.ex_alu.result_sll[5] ),
    .X(_00343_));
 sky130_fd_sc_hd__or2_1 _08292_ (.A(net386),
    .B(_04514_),
    .X(_04535_));
 sky130_fd_sc_hd__and2_1 _08293_ (.A(net374),
    .B(_04530_),
    .X(_04536_));
 sky130_fd_sc_hd__a22o_1 _08294_ (.A1(net627),
    .A2(\core_pipeline.decode_to_execute_imm_data[6] ),
    .B1(\core_pipeline.decode_to_execute_pc[6] ),
    .B2(net629),
    .X(_04537_));
 sky130_fd_sc_hd__a21o_4 _08295_ (.A1(_03860_),
    .A2(net432),
    .B1(_04537_),
    .X(_04538_));
 sky130_fd_sc_hd__a211o_1 _08296_ (.A1(net377),
    .A2(_04538_),
    .B1(_04536_),
    .C1(net379),
    .X(_04539_));
 sky130_fd_sc_hd__o21ai_2 _08297_ (.A1(net380),
    .A2(_04525_),
    .B1(_04539_),
    .Y(_04540_));
 sky130_fd_sc_hd__nand2_1 _08298_ (.A(net386),
    .B(_04540_),
    .Y(_04541_));
 sky130_fd_sc_hd__and3_1 _08299_ (.A(net397),
    .B(_04535_),
    .C(_04541_),
    .X(_04542_));
 sky130_fd_sc_hd__a22o_1 _08300_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_sll[6] ),
    .A2(net435),
    .B1(net280),
    .B2(_04542_),
    .X(_00344_));
 sky130_fd_sc_hd__and2_1 _08301_ (.A(net374),
    .B(_04538_),
    .X(_04543_));
 sky130_fd_sc_hd__a22o_1 _08302_ (.A1(net628),
    .A2(\core_pipeline.decode_to_execute_imm_data[7] ),
    .B1(\core_pipeline.decode_to_execute_pc[7] ),
    .B2(net630),
    .X(_04544_));
 sky130_fd_sc_hd__a21oi_4 _08303_ (.A1(_03863_),
    .A2(net432),
    .B1(_04544_),
    .Y(_04545_));
 sky130_fd_sc_hd__nor2_1 _08304_ (.A(net374),
    .B(_04545_),
    .Y(_04546_));
 sky130_fd_sc_hd__or2_1 _08305_ (.A(_04543_),
    .B(_04546_),
    .X(_04547_));
 sky130_fd_sc_hd__mux2_1 _08306_ (.A0(_04532_),
    .A1(_04547_),
    .S(net380),
    .X(_04548_));
 sky130_fd_sc_hd__or2_1 _08307_ (.A(net384),
    .B(_04548_),
    .X(_04549_));
 sky130_fd_sc_hd__o21ai_1 _08308_ (.A1(net388),
    .A2(_04520_),
    .B1(_04549_),
    .Y(_04550_));
 sky130_fd_sc_hd__nor2_1 _08309_ (.A(net395),
    .B(_04550_),
    .Y(_04551_));
 sky130_fd_sc_hd__a22o_1 _08310_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_sll[7] ),
    .A2(net435),
    .B1(net280),
    .B2(_04551_),
    .X(_00345_));
 sky130_fd_sc_hd__a22o_2 _08311_ (.A1(net627),
    .A2(\core_pipeline.decode_to_execute_imm_data[8] ),
    .B1(\core_pipeline.decode_to_execute_pc[8] ),
    .B2(net629),
    .X(_04552_));
 sky130_fd_sc_hd__a21oi_4 _08312_ (.A1(_03854_),
    .A2(net431),
    .B1(_04552_),
    .Y(_04553_));
 sky130_fd_sc_hd__inv_2 _08313_ (.A(_04553_),
    .Y(_04554_));
 sky130_fd_sc_hd__nor2_1 _08314_ (.A(net372),
    .B(_04553_),
    .Y(_04555_));
 sky130_fd_sc_hd__nor2_1 _08315_ (.A(net377),
    .B(_04545_),
    .Y(_04556_));
 sky130_fd_sc_hd__nor2_1 _08316_ (.A(_04555_),
    .B(_04556_),
    .Y(_04557_));
 sky130_fd_sc_hd__a211o_1 _08317_ (.A1(net377),
    .A2(_04538_),
    .B1(_04536_),
    .C1(net380),
    .X(_04558_));
 sky130_fd_sc_hd__o31a_1 _08318_ (.A1(net379),
    .A2(_04555_),
    .A3(_04556_),
    .B1(_04558_),
    .X(_04559_));
 sky130_fd_sc_hd__mux2_2 _08319_ (.A0(_04526_),
    .A1(_04559_),
    .S(net388),
    .X(_04560_));
 sky130_fd_sc_hd__nor2_2 _08320_ (.A(net396),
    .B(net385),
    .Y(_04561_));
 sky130_fd_sc_hd__a22o_1 _08321_ (.A1(net396),
    .A2(_04560_),
    .B1(_04561_),
    .B2(_04497_),
    .X(_04562_));
 sky130_fd_sc_hd__a22o_1 _08322_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_sll[8] ),
    .A2(net436),
    .B1(net280),
    .B2(_04562_),
    .X(_00346_));
 sky130_fd_sc_hd__nor2_1 _08323_ (.A(net375),
    .B(_04553_),
    .Y(_04563_));
 sky130_fd_sc_hd__a22o_2 _08324_ (.A1(net627),
    .A2(\core_pipeline.decode_to_execute_imm_data[9] ),
    .B1(\core_pipeline.decode_to_execute_pc[9] ),
    .B2(net629),
    .X(_04564_));
 sky130_fd_sc_hd__a21oi_4 _08325_ (.A1(_03849_),
    .A2(net431),
    .B1(_04564_),
    .Y(_04565_));
 sky130_fd_sc_hd__inv_2 _08326_ (.A(_04565_),
    .Y(_04566_));
 sky130_fd_sc_hd__nor2_1 _08327_ (.A(net372),
    .B(_04565_),
    .Y(_04567_));
 sky130_fd_sc_hd__or2_1 _08328_ (.A(_04563_),
    .B(_04567_),
    .X(_04568_));
 sky130_fd_sc_hd__mux2_1 _08329_ (.A0(_04547_),
    .A1(_04568_),
    .S(net380),
    .X(_04569_));
 sky130_fd_sc_hd__mux2_2 _08330_ (.A0(_04533_),
    .A1(_04569_),
    .S(net388),
    .X(_04570_));
 sky130_fd_sc_hd__a22o_1 _08331_ (.A1(_04507_),
    .A2(_04561_),
    .B1(_04570_),
    .B2(net397),
    .X(_04571_));
 sky130_fd_sc_hd__a22o_1 _08332_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_sll[9] ),
    .A2(net435),
    .B1(net280),
    .B2(_04571_),
    .X(_00347_));
 sky130_fd_sc_hd__nor2_1 _08333_ (.A(net375),
    .B(_04565_),
    .Y(_04572_));
 sky130_fd_sc_hd__a22o_1 _08334_ (.A1(net628),
    .A2(\core_pipeline.decode_to_execute_imm_data[10] ),
    .B1(\core_pipeline.decode_to_execute_pc[10] ),
    .B2(net630),
    .X(_04573_));
 sky130_fd_sc_hd__a21o_4 _08335_ (.A1(_03842_),
    .A2(net431),
    .B1(_04573_),
    .X(_04574_));
 sky130_fd_sc_hd__a21oi_1 _08336_ (.A1(net375),
    .A2(_04574_),
    .B1(_04572_),
    .Y(_04575_));
 sky130_fd_sc_hd__mux2_1 _08337_ (.A0(_04557_),
    .A1(_04575_),
    .S(net381),
    .X(_04576_));
 sky130_fd_sc_hd__mux2_1 _08338_ (.A0(_04540_),
    .A1(_04576_),
    .S(net386),
    .X(_04577_));
 sky130_fd_sc_hd__a2bb2o_1 _08339_ (.A1_N(net394),
    .A2_N(_04577_),
    .B1(_04561_),
    .B2(_04514_),
    .X(_04578_));
 sky130_fd_sc_hd__a22o_1 _08340_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_sll[10] ),
    .A2(net436),
    .B1(net280),
    .B2(_04578_),
    .X(_00348_));
 sky130_fd_sc_hd__and2_1 _08341_ (.A(net372),
    .B(_04574_),
    .X(_04579_));
 sky130_fd_sc_hd__a22o_1 _08342_ (.A1(net627),
    .A2(\core_pipeline.decode_to_execute_imm_data[11] ),
    .B1(\core_pipeline.decode_to_execute_pc[11] ),
    .B2(net629),
    .X(_04580_));
 sky130_fd_sc_hd__a21oi_4 _08343_ (.A1(_03845_),
    .A2(net431),
    .B1(_04580_),
    .Y(_04581_));
 sky130_fd_sc_hd__inv_2 _08344_ (.A(_04581_),
    .Y(_04582_));
 sky130_fd_sc_hd__nor2_1 _08345_ (.A(net372),
    .B(_04581_),
    .Y(_04583_));
 sky130_fd_sc_hd__or2_1 _08346_ (.A(_04579_),
    .B(_04583_),
    .X(_04584_));
 sky130_fd_sc_hd__mux2_1 _08347_ (.A0(_04568_),
    .A1(_04584_),
    .S(net380),
    .X(_04585_));
 sky130_fd_sc_hd__mux2_1 _08348_ (.A0(_04548_),
    .A1(_04585_),
    .S(net388),
    .X(_04586_));
 sky130_fd_sc_hd__a22o_2 _08349_ (.A1(_04520_),
    .A2(_04561_),
    .B1(_04586_),
    .B2(net396),
    .X(_04587_));
 sky130_fd_sc_hd__a22o_1 _08350_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_sll[11] ),
    .A2(net436),
    .B1(net280),
    .B2(_04587_),
    .X(_00349_));
 sky130_fd_sc_hd__nor2_1 _08351_ (.A(net375),
    .B(_04581_),
    .Y(_04588_));
 sky130_fd_sc_hd__a22o_1 _08352_ (.A1(net627),
    .A2(\core_pipeline.decode_to_execute_imm_data[12] ),
    .B1(\core_pipeline.decode_to_execute_pc[12] ),
    .B2(net629),
    .X(_04589_));
 sky130_fd_sc_hd__a21oi_4 _08353_ (.A1(_03838_),
    .A2(net431),
    .B1(_04589_),
    .Y(_04590_));
 sky130_fd_sc_hd__nor2_1 _08354_ (.A(net372),
    .B(_04590_),
    .Y(_04591_));
 sky130_fd_sc_hd__nor2_1 _08355_ (.A(_04588_),
    .B(_04591_),
    .Y(_04592_));
 sky130_fd_sc_hd__mux2_1 _08356_ (.A0(_04575_),
    .A1(_04592_),
    .S(net381),
    .X(_04593_));
 sky130_fd_sc_hd__inv_2 _08357_ (.A(_04593_),
    .Y(_04594_));
 sky130_fd_sc_hd__mux2_1 _08358_ (.A0(_04559_),
    .A1(_04594_),
    .S(net386),
    .X(_04595_));
 sky130_fd_sc_hd__mux2_2 _08359_ (.A0(_04527_),
    .A1(_04595_),
    .S(net397),
    .X(_04596_));
 sky130_fd_sc_hd__a22o_1 _08360_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_sll[12] ),
    .A2(net436),
    .B1(net280),
    .B2(_04596_),
    .X(_00350_));
 sky130_fd_sc_hd__nor2_1 _08361_ (.A(net376),
    .B(_04590_),
    .Y(_04597_));
 sky130_fd_sc_hd__a22o_2 _08362_ (.A1(net627),
    .A2(\core_pipeline.decode_to_execute_imm_data[13] ),
    .B1(\core_pipeline.decode_to_execute_pc[13] ),
    .B2(net629),
    .X(_04598_));
 sky130_fd_sc_hd__a21oi_4 _08363_ (.A1(_03832_),
    .A2(net431),
    .B1(_04598_),
    .Y(_04599_));
 sky130_fd_sc_hd__nor2_1 _08364_ (.A(net373),
    .B(_04599_),
    .Y(_04600_));
 sky130_fd_sc_hd__nor2_1 _08365_ (.A(_04597_),
    .B(_04600_),
    .Y(_04601_));
 sky130_fd_sc_hd__inv_2 _08366_ (.A(_04601_),
    .Y(_04602_));
 sky130_fd_sc_hd__mux2_1 _08367_ (.A0(_04584_),
    .A1(_04602_),
    .S(net381),
    .X(_04603_));
 sky130_fd_sc_hd__mux2_1 _08368_ (.A0(_04569_),
    .A1(_04603_),
    .S(net386),
    .X(_04604_));
 sky130_fd_sc_hd__mux2_2 _08369_ (.A0(_04534_),
    .A1(_04604_),
    .S(net396),
    .X(_04605_));
 sky130_fd_sc_hd__a22o_1 _08370_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_sll[13] ),
    .A2(net436),
    .B1(net280),
    .B2(_04605_),
    .X(_00351_));
 sky130_fd_sc_hd__nor2_1 _08371_ (.A(net375),
    .B(_04599_),
    .Y(_04606_));
 sky130_fd_sc_hd__a22o_2 _08372_ (.A1(net627),
    .A2(\core_pipeline.decode_to_execute_imm_data[14] ),
    .B1(\core_pipeline.decode_to_execute_pc[14] ),
    .B2(net629),
    .X(_04607_));
 sky130_fd_sc_hd__a21oi_4 _08373_ (.A1(_03828_),
    .A2(net431),
    .B1(_04607_),
    .Y(_04608_));
 sky130_fd_sc_hd__nor2_1 _08374_ (.A(net372),
    .B(_04608_),
    .Y(_04609_));
 sky130_fd_sc_hd__nor2_1 _08375_ (.A(_04606_),
    .B(_04609_),
    .Y(_04610_));
 sky130_fd_sc_hd__mux2_1 _08376_ (.A0(_04592_),
    .A1(_04610_),
    .S(net382),
    .X(_04611_));
 sky130_fd_sc_hd__mux2_1 _08377_ (.A0(_04576_),
    .A1(_04611_),
    .S(net386),
    .X(_04612_));
 sky130_fd_sc_hd__nor2_1 _08378_ (.A(net394),
    .B(_04612_),
    .Y(_04613_));
 sky130_fd_sc_hd__a31o_1 _08379_ (.A1(net394),
    .A2(_04535_),
    .A3(_04541_),
    .B1(_04613_),
    .X(_04614_));
 sky130_fd_sc_hd__a22o_1 _08380_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_sll[14] ),
    .A2(net436),
    .B1(net280),
    .B2(_04614_),
    .X(_00352_));
 sky130_fd_sc_hd__nand2_1 _08381_ (.A(net385),
    .B(_04585_),
    .Y(_04615_));
 sky130_fd_sc_hd__nor2_1 _08382_ (.A(net375),
    .B(_04608_),
    .Y(_04616_));
 sky130_fd_sc_hd__a22o_1 _08383_ (.A1(net627),
    .A2(\core_pipeline.decode_to_execute_imm_data[15] ),
    .B1(\core_pipeline.decode_to_execute_pc[15] ),
    .B2(net629),
    .X(_04617_));
 sky130_fd_sc_hd__a21o_4 _08384_ (.A1(_03824_),
    .A2(net431),
    .B1(_04617_),
    .X(_04618_));
 sky130_fd_sc_hd__a21oi_1 _08385_ (.A1(net375),
    .A2(_04618_),
    .B1(_04616_),
    .Y(_04619_));
 sky130_fd_sc_hd__mux2_1 _08386_ (.A0(_04601_),
    .A1(_04619_),
    .S(net381),
    .X(_04620_));
 sky130_fd_sc_hd__o21a_1 _08387_ (.A1(net385),
    .A2(_04620_),
    .B1(_04615_),
    .X(_04621_));
 sky130_fd_sc_hd__mux2_2 _08388_ (.A0(_04550_),
    .A1(_04621_),
    .S(net399),
    .X(_04622_));
 sky130_fd_sc_hd__a2bb2o_1 _08389_ (.A1_N(_04622_),
    .A2_N(_04482_),
    .B1(net436),
    .B2(\core_pipeline.pipeline_execute.ex_alu.result_sll[15] ),
    .X(_00353_));
 sky130_fd_sc_hd__or3_2 _08390_ (.A(_03460_),
    .B(_03484_),
    .C(_03636_),
    .X(_04623_));
 sky130_fd_sc_hd__nor2_1 _08391_ (.A(\core_pipeline.fetch_to_decode_instruction[5] ),
    .B(_03444_),
    .Y(_04624_));
 sky130_fd_sc_hd__nand2_1 _08392_ (.A(_03322_),
    .B(_03443_),
    .Y(_04625_));
 sky130_fd_sc_hd__nor2_2 _08393_ (.A(\core_pipeline.fetch_to_decode_instruction[4] ),
    .B(_04625_),
    .Y(_04626_));
 sky130_fd_sc_hd__o31a_2 _08394_ (.A1(_03437_),
    .A2(_04623_),
    .A3(_04626_),
    .B1(net142),
    .X(_04627_));
 sky130_fd_sc_hd__a22o_1 _08395_ (.A1(\core_pipeline.decode_to_execute_rd_address[4] ),
    .A2(net127),
    .B1(_04627_),
    .B2(net658),
    .X(_00354_));
 sky130_fd_sc_hd__a22o_1 _08396_ (.A1(\core_pipeline.decode_to_execute_rd_address[3] ),
    .A2(net127),
    .B1(_04627_),
    .B2(net654),
    .X(_00355_));
 sky130_fd_sc_hd__a22o_1 _08397_ (.A1(\core_pipeline.decode_to_execute_rd_address[2] ),
    .A2(net127),
    .B1(_04627_),
    .B2(\core_pipeline.fetch_to_decode_instruction[9] ),
    .X(_00356_));
 sky130_fd_sc_hd__a22o_1 _08398_ (.A1(\core_pipeline.decode_to_execute_rd_address[1] ),
    .A2(net127),
    .B1(_04627_),
    .B2(\core_pipeline.fetch_to_decode_instruction[8] ),
    .X(_00357_));
 sky130_fd_sc_hd__a22o_1 _08399_ (.A1(\core_pipeline.decode_to_execute_rd_address[0] ),
    .A2(net127),
    .B1(_04627_),
    .B2(net655),
    .X(_00358_));
 sky130_fd_sc_hd__or3_1 _08400_ (.A(net127),
    .B(_03437_),
    .C(_04626_),
    .X(_04628_));
 sky130_fd_sc_hd__o21a_1 _08401_ (.A1(\core_pipeline.decode_to_execute_write_select[1] ),
    .A2(net143),
    .B1(_04628_),
    .X(_00359_));
 sky130_fd_sc_hd__or2_2 _08402_ (.A(net127),
    .B(_03437_),
    .X(_04629_));
 sky130_fd_sc_hd__o22a_1 _08403_ (.A1(\core_pipeline.decode_to_execute_write_select[0] ),
    .A2(net142),
    .B1(_03484_),
    .B2(_04629_),
    .X(_00360_));
 sky130_fd_sc_hd__mux2_1 _08404_ (.A0(\core_pipeline.decode_to_execute_bypass_memory ),
    .A1(_04623_),
    .S(net142),
    .X(_00361_));
 sky130_fd_sc_hd__or4_2 _08405_ (.A(net626),
    .B(net581),
    .C(net575),
    .D(net568),
    .X(_04630_));
 sky130_fd_sc_hd__nor2_2 _08406_ (.A(net602),
    .B(_04630_),
    .Y(_04631_));
 sky130_fd_sc_hd__nand2_1 _08407_ (.A(\core_pipeline.fetch_to_decode_instruction[13] ),
    .B(_04631_),
    .Y(_04632_));
 sky130_fd_sc_hd__a32o_1 _08408_ (.A1(_03448_),
    .A2(_03632_),
    .A3(_04632_),
    .B1(net132),
    .B2(\core_pipeline.decode_to_execute_csr_write ),
    .X(_00362_));
 sky130_fd_sc_hd__a32o_1 _08409_ (.A1(_03448_),
    .A2(_03486_),
    .A3(_03632_),
    .B1(net132),
    .B2(\core_pipeline.decode_to_execute_csr_read ),
    .X(_00363_));
 sky130_fd_sc_hd__nand2_1 _08410_ (.A(\core_pipeline.fetch_to_decode_instruction[14] ),
    .B(\core_pipeline.fetch_to_decode_instruction[12] ),
    .Y(_04633_));
 sky130_fd_sc_hd__a31o_1 _08411_ (.A1(\core_pipeline.fetch_to_decode_instruction[14] ),
    .A2(_03321_),
    .A3(\core_pipeline.fetch_to_decode_instruction[12] ),
    .B1(\core_pipeline.fetch_to_decode_instruction[5] ),
    .X(_04634_));
 sky130_fd_sc_hd__a31o_1 _08412_ (.A1(\core_pipeline.decode_to_csr_read_address[10] ),
    .A2(_03460_),
    .A3(_04634_),
    .B1(net126),
    .X(_04635_));
 sky130_fd_sc_hd__o21a_1 _08413_ (.A1(net632),
    .A2(net142),
    .B1(_04635_),
    .X(_04636_));
 sky130_fd_sc_hd__a31o_1 _08414_ (.A1(\core_pipeline.fetch_to_decode_instruction[13] ),
    .A2(\core_pipeline.fetch_to_decode_instruction[12] ),
    .A3(_03632_),
    .B1(_04636_),
    .X(_00364_));
 sky130_fd_sc_hd__a21o_1 _08415_ (.A1(\core_pipeline.fetch_to_decode_instruction[14] ),
    .A2(_03460_),
    .B1(net126),
    .X(_04637_));
 sky130_fd_sc_hd__o32a_1 _08416_ (.A1(_03451_),
    .A2(_03639_),
    .A3(_04637_),
    .B1(net142),
    .B2(\core_pipeline.decode_to_execute_alu_function[2] ),
    .X(_00365_));
 sky130_fd_sc_hd__a211o_1 _08417_ (.A1(\core_pipeline.fetch_to_decode_instruction[13] ),
    .A2(_03460_),
    .B1(_03639_),
    .C1(_03451_),
    .X(_04638_));
 sky130_fd_sc_hd__mux2_1 _08418_ (.A0(\core_pipeline.decode_to_execute_alu_function[1] ),
    .A1(_04638_),
    .S(net140),
    .X(_00366_));
 sky130_fd_sc_hd__a32o_1 _08419_ (.A1(\core_pipeline.fetch_to_decode_instruction[13] ),
    .A2(\core_pipeline.fetch_to_decode_instruction[12] ),
    .A3(_03632_),
    .B1(net126),
    .B2(\core_pipeline.decode_to_execute_alu_function[0] ),
    .X(_04639_));
 sky130_fd_sc_hd__a31o_1 _08420_ (.A1(\core_pipeline.fetch_to_decode_instruction[12] ),
    .A2(net142),
    .A3(_03460_),
    .B1(_04639_),
    .X(_00367_));
 sky130_fd_sc_hd__nand2_2 _08421_ (.A(_03438_),
    .B(_04625_),
    .Y(_04640_));
 sky130_fd_sc_hd__o21a_4 _08422_ (.A1(_03442_),
    .A2(_04640_),
    .B1(\core_pipeline.decode_to_csr_read_address[11] ),
    .X(_04641_));
 sky130_fd_sc_hd__o311a_1 _08423_ (.A1(_03442_),
    .A2(_03637_),
    .A3(_04640_),
    .B1(net149),
    .C1(\core_pipeline.decode_to_csr_read_address[11] ),
    .X(_04642_));
 sky130_fd_sc_hd__a21o_1 _08424_ (.A1(\core_pipeline.decode_to_execute_imm_data[31] ),
    .A2(net126),
    .B1(_04642_),
    .X(_00368_));
 sky130_fd_sc_hd__and3_4 _08425_ (.A(\core_pipeline.fetch_to_decode_instruction[3] ),
    .B(\core_pipeline.decode_to_csr_read_address[11] ),
    .C(_03437_),
    .X(_04643_));
 sky130_fd_sc_hd__or2_4 _08426_ (.A(net128),
    .B(_04641_),
    .X(_04644_));
 sky130_fd_sc_hd__a211o_1 _08427_ (.A1(\core_pipeline.decode_to_csr_read_address[10] ),
    .A2(_03636_),
    .B1(_04643_),
    .C1(net128),
    .X(_04645_));
 sky130_fd_sc_hd__o22a_1 _08428_ (.A1(\core_pipeline.decode_to_execute_imm_data[30] ),
    .A2(net149),
    .B1(_04641_),
    .B2(_04645_),
    .X(_00369_));
 sky130_fd_sc_hd__a211o_1 _08429_ (.A1(\core_pipeline.decode_to_csr_read_address[9] ),
    .A2(_03636_),
    .B1(_04643_),
    .C1(net128),
    .X(_04646_));
 sky130_fd_sc_hd__o22a_1 _08430_ (.A1(\core_pipeline.decode_to_execute_imm_data[29] ),
    .A2(net150),
    .B1(_04641_),
    .B2(_04646_),
    .X(_00370_));
 sky130_fd_sc_hd__a211o_1 _08431_ (.A1(\core_pipeline.decode_to_csr_read_address[8] ),
    .A2(_03636_),
    .B1(_04643_),
    .C1(net128),
    .X(_04647_));
 sky130_fd_sc_hd__o22a_1 _08432_ (.A1(\core_pipeline.decode_to_execute_imm_data[28] ),
    .A2(net150),
    .B1(_04641_),
    .B2(_04647_),
    .X(_00371_));
 sky130_fd_sc_hd__a211o_1 _08433_ (.A1(\core_pipeline.decode_to_csr_read_address[7] ),
    .A2(_03636_),
    .B1(_04643_),
    .C1(net126),
    .X(_04648_));
 sky130_fd_sc_hd__o22a_1 _08434_ (.A1(\core_pipeline.decode_to_execute_imm_data[27] ),
    .A2(net149),
    .B1(_04641_),
    .B2(_04648_),
    .X(_00372_));
 sky130_fd_sc_hd__a211o_1 _08435_ (.A1(\core_pipeline.decode_to_csr_read_address[6] ),
    .A2(_03636_),
    .B1(_04643_),
    .C1(net128),
    .X(_04649_));
 sky130_fd_sc_hd__o22a_1 _08436_ (.A1(\core_pipeline.decode_to_execute_imm_data[26] ),
    .A2(net149),
    .B1(_04641_),
    .B2(_04649_),
    .X(_00373_));
 sky130_fd_sc_hd__a211o_1 _08437_ (.A1(\core_pipeline.decode_to_csr_read_address[5] ),
    .A2(_03636_),
    .B1(_04643_),
    .C1(net128),
    .X(_04650_));
 sky130_fd_sc_hd__o22a_1 _08438_ (.A1(\core_pipeline.decode_to_execute_imm_data[25] ),
    .A2(net150),
    .B1(_04641_),
    .B2(_04650_),
    .X(_00374_));
 sky130_fd_sc_hd__a211o_1 _08439_ (.A1(net511),
    .A2(_03636_),
    .B1(_04643_),
    .C1(net128),
    .X(_04651_));
 sky130_fd_sc_hd__o22a_1 _08440_ (.A1(\core_pipeline.decode_to_execute_imm_data[24] ),
    .A2(net150),
    .B1(_04641_),
    .B2(_04651_),
    .X(_00375_));
 sky130_fd_sc_hd__a21o_1 _08441_ (.A1(net515),
    .A2(_03636_),
    .B1(_04643_),
    .X(_04652_));
 sky130_fd_sc_hd__o22a_1 _08442_ (.A1(\core_pipeline.decode_to_execute_imm_data[23] ),
    .A2(net150),
    .B1(_04644_),
    .B2(_04652_),
    .X(_00376_));
 sky130_fd_sc_hd__a21o_1 _08443_ (.A1(net521),
    .A2(_03636_),
    .B1(_04643_),
    .X(_04653_));
 sky130_fd_sc_hd__o22a_1 _08444_ (.A1(\core_pipeline.decode_to_execute_imm_data[22] ),
    .A2(net150),
    .B1(_04644_),
    .B2(_04653_),
    .X(_00377_));
 sky130_fd_sc_hd__a211o_1 _08445_ (.A1(net543),
    .A2(_03636_),
    .B1(_04643_),
    .C1(net128),
    .X(_04654_));
 sky130_fd_sc_hd__o22a_1 _08446_ (.A1(\core_pipeline.decode_to_execute_imm_data[21] ),
    .A2(net149),
    .B1(_04641_),
    .B2(_04654_),
    .X(_00378_));
 sky130_fd_sc_hd__a211o_1 _08447_ (.A1(net566),
    .A2(_03636_),
    .B1(_04643_),
    .C1(net128),
    .X(_04655_));
 sky130_fd_sc_hd__o22a_1 _08448_ (.A1(\core_pipeline.decode_to_execute_imm_data[20] ),
    .A2(net150),
    .B1(_04641_),
    .B2(_04655_),
    .X(_00379_));
 sky130_fd_sc_hd__and2_1 _08449_ (.A(net567),
    .B(_03637_),
    .X(_04656_));
 sky130_fd_sc_hd__o22a_1 _08450_ (.A1(\core_pipeline.decode_to_execute_imm_data[19] ),
    .A2(net150),
    .B1(_04644_),
    .B2(_04656_),
    .X(_00380_));
 sky130_fd_sc_hd__and2_1 _08451_ (.A(net572),
    .B(_03637_),
    .X(_04657_));
 sky130_fd_sc_hd__o22a_1 _08452_ (.A1(\core_pipeline.decode_to_execute_imm_data[18] ),
    .A2(net151),
    .B1(_04644_),
    .B2(_04657_),
    .X(_00381_));
 sky130_fd_sc_hd__and2_1 _08453_ (.A(net578),
    .B(_03637_),
    .X(_04658_));
 sky130_fd_sc_hd__o22a_1 _08454_ (.A1(\core_pipeline.decode_to_execute_imm_data[17] ),
    .A2(net150),
    .B1(_04644_),
    .B2(_04658_),
    .X(_00382_));
 sky130_fd_sc_hd__and2_1 _08455_ (.A(\core_pipeline.decode_to_regfile_rs1_address[1] ),
    .B(_03637_),
    .X(_04659_));
 sky130_fd_sc_hd__o22a_1 _08456_ (.A1(\core_pipeline.decode_to_execute_imm_data[16] ),
    .A2(net150),
    .B1(_04644_),
    .B2(_04659_),
    .X(_00383_));
 sky130_fd_sc_hd__and2_1 _08457_ (.A(net614),
    .B(_03637_),
    .X(_04660_));
 sky130_fd_sc_hd__o22a_1 _08458_ (.A1(\core_pipeline.decode_to_execute_imm_data[15] ),
    .A2(net152),
    .B1(_04644_),
    .B2(_04660_),
    .X(_00384_));
 sky130_fd_sc_hd__and2_1 _08459_ (.A(\core_pipeline.fetch_to_decode_instruction[14] ),
    .B(_03637_),
    .X(_04661_));
 sky130_fd_sc_hd__o22a_1 _08460_ (.A1(\core_pipeline.decode_to_execute_imm_data[14] ),
    .A2(net150),
    .B1(_04644_),
    .B2(_04661_),
    .X(_00385_));
 sky130_fd_sc_hd__o21a_1 _08461_ (.A1(\core_pipeline.decode_to_execute_imm_data[13] ),
    .A2(net150),
    .B1(_04644_),
    .X(_04662_));
 sky130_fd_sc_hd__a31o_1 _08462_ (.A1(\core_pipeline.fetch_to_decode_instruction[13] ),
    .A2(net150),
    .A3(_03637_),
    .B1(_04662_),
    .X(_00386_));
 sky130_fd_sc_hd__o21a_1 _08463_ (.A1(\core_pipeline.decode_to_execute_imm_data[12] ),
    .A2(net152),
    .B1(_04644_),
    .X(_04663_));
 sky130_fd_sc_hd__a31o_1 _08464_ (.A1(\core_pipeline.fetch_to_decode_instruction[12] ),
    .A2(net152),
    .A3(_03637_),
    .B1(_04663_),
    .X(_00387_));
 sky130_fd_sc_hd__and2b_2 _08465_ (.A_N(\core_pipeline.fetch_to_decode_instruction[6] ),
    .B(_03442_),
    .X(_04664_));
 sky130_fd_sc_hd__o21a_1 _08466_ (.A1(_04640_),
    .A2(_04664_),
    .B1(\core_pipeline.decode_to_csr_read_address[11] ),
    .X(_04665_));
 sky130_fd_sc_hd__a221o_2 _08467_ (.A1(\core_pipeline.fetch_to_decode_instruction[7] ),
    .A2(_03445_),
    .B1(_03635_),
    .B2(net566),
    .C1(_04665_),
    .X(_04666_));
 sky130_fd_sc_hd__mux2_1 _08468_ (.A0(\core_pipeline.decode_to_execute_imm_data[11] ),
    .A1(_04666_),
    .S(net152),
    .X(_00388_));
 sky130_fd_sc_hd__or2_2 _08469_ (.A(_03437_),
    .B(_04624_),
    .X(_04667_));
 sky130_fd_sc_hd__o21a_4 _08470_ (.A1(_03442_),
    .A2(_04667_),
    .B1(net149),
    .X(_04668_));
 sky130_fd_sc_hd__a22o_1 _08471_ (.A1(\core_pipeline.decode_to_execute_imm_data[10] ),
    .A2(net128),
    .B1(_04668_),
    .B2(\core_pipeline.decode_to_csr_read_address[10] ),
    .X(_00389_));
 sky130_fd_sc_hd__a22o_1 _08472_ (.A1(\core_pipeline.decode_to_execute_imm_data[9] ),
    .A2(net128),
    .B1(_04668_),
    .B2(\core_pipeline.decode_to_csr_read_address[9] ),
    .X(_00390_));
 sky130_fd_sc_hd__a22o_1 _08473_ (.A1(\core_pipeline.decode_to_execute_imm_data[8] ),
    .A2(net128),
    .B1(_04668_),
    .B2(\core_pipeline.decode_to_csr_read_address[8] ),
    .X(_00391_));
 sky130_fd_sc_hd__a22o_1 _08474_ (.A1(\core_pipeline.decode_to_execute_imm_data[7] ),
    .A2(net126),
    .B1(_04668_),
    .B2(\core_pipeline.decode_to_csr_read_address[7] ),
    .X(_00392_));
 sky130_fd_sc_hd__a22o_1 _08475_ (.A1(\core_pipeline.decode_to_execute_imm_data[6] ),
    .A2(net128),
    .B1(_04668_),
    .B2(\core_pipeline.decode_to_csr_read_address[6] ),
    .X(_00393_));
 sky130_fd_sc_hd__a22o_1 _08476_ (.A1(\core_pipeline.decode_to_execute_imm_data[5] ),
    .A2(net126),
    .B1(_04668_),
    .B2(\core_pipeline.decode_to_csr_read_address[5] ),
    .X(_00394_));
 sky130_fd_sc_hd__and3_2 _08477_ (.A(\core_pipeline.fetch_to_decode_instruction[14] ),
    .B(_03448_),
    .C(_03451_),
    .X(_04669_));
 sky130_fd_sc_hd__a22o_1 _08478_ (.A1(\core_pipeline.decode_to_csr_read_address[4] ),
    .A2(_04667_),
    .B1(_04669_),
    .B2(net567),
    .X(_04670_));
 sky130_fd_sc_hd__a211o_1 _08479_ (.A1(\core_pipeline.fetch_to_decode_instruction[11] ),
    .A2(_03442_),
    .B1(_04670_),
    .C1(net126),
    .X(_04671_));
 sky130_fd_sc_hd__o21a_1 _08480_ (.A1(\core_pipeline.decode_to_execute_imm_data[4] ),
    .A2(net152),
    .B1(_04671_),
    .X(_00395_));
 sky130_fd_sc_hd__and2_1 _08481_ (.A(net515),
    .B(_04667_),
    .X(_04672_));
 sky130_fd_sc_hd__a221o_1 _08482_ (.A1(\core_pipeline.fetch_to_decode_instruction[10] ),
    .A2(_03442_),
    .B1(_04669_),
    .B2(net572),
    .C1(_04672_),
    .X(_04673_));
 sky130_fd_sc_hd__mux2_1 _08483_ (.A0(\core_pipeline.decode_to_execute_imm_data[3] ),
    .A1(_04673_),
    .S(net149),
    .X(_00396_));
 sky130_fd_sc_hd__a22o_1 _08484_ (.A1(\core_pipeline.fetch_to_decode_instruction[9] ),
    .A2(_03442_),
    .B1(_04667_),
    .B2(net521),
    .X(_04674_));
 sky130_fd_sc_hd__a21o_1 _08485_ (.A1(net578),
    .A2(_04669_),
    .B1(_04674_),
    .X(_04675_));
 sky130_fd_sc_hd__mux2_1 _08486_ (.A0(\core_pipeline.decode_to_execute_imm_data[2] ),
    .A1(_04675_),
    .S(net149),
    .X(_00397_));
 sky130_fd_sc_hd__and2_1 _08487_ (.A(net543),
    .B(_04667_),
    .X(_04676_));
 sky130_fd_sc_hd__a221o_1 _08488_ (.A1(\core_pipeline.fetch_to_decode_instruction[8] ),
    .A2(_03442_),
    .B1(_04669_),
    .B2(\core_pipeline.decode_to_regfile_rs1_address[1] ),
    .C1(_04676_),
    .X(_04677_));
 sky130_fd_sc_hd__mux2_1 _08489_ (.A0(\core_pipeline.decode_to_execute_imm_data[1] ),
    .A1(_04677_),
    .S(net139),
    .X(_00398_));
 sky130_fd_sc_hd__a22o_1 _08490_ (.A1(net566),
    .A2(_04640_),
    .B1(_04664_),
    .B2(\core_pipeline.fetch_to_decode_instruction[7] ),
    .X(_04678_));
 sky130_fd_sc_hd__a211o_1 _08491_ (.A1(net614),
    .A2(_04669_),
    .B1(_04678_),
    .C1(net126),
    .X(_04679_));
 sky130_fd_sc_hd__o21a_1 _08492_ (.A1(\core_pipeline.decode_to_execute_imm_data[0] ),
    .A2(net152),
    .B1(_04679_),
    .X(_00399_));
 sky130_fd_sc_hd__nor2_8 _08493_ (.A(net522),
    .B(net516),
    .Y(_04680_));
 sky130_fd_sc_hd__nor2_8 _08494_ (.A(net558),
    .B(net535),
    .Y(_04681_));
 sky130_fd_sc_hd__nand2_8 _08495_ (.A(_03328_),
    .B(net430),
    .Y(_04682_));
 sky130_fd_sc_hd__nor2_8 _08496_ (.A(net565),
    .B(_04682_),
    .Y(_04683_));
 sky130_fd_sc_hd__nand2_8 _08497_ (.A(_04680_),
    .B(net427),
    .Y(_04684_));
 sky130_fd_sc_hd__nand2_1 _08498_ (.A(\core_pipeline.decode_to_csr_read_address[9] ),
    .B(\core_pipeline.decode_to_csr_read_address[8] ),
    .Y(_04685_));
 sky130_fd_sc_hd__or3b_4 _08499_ (.A(_04685_),
    .B(\core_pipeline.decode_to_csr_read_address[10] ),
    .C_N(\core_pipeline.decode_to_csr_read_address[11] ),
    .X(_04686_));
 sky130_fd_sc_hd__nand2b_1 _08500_ (.A_N(\core_pipeline.decode_to_csr_read_address[5] ),
    .B(\core_pipeline.decode_to_csr_read_address[7] ),
    .Y(_04687_));
 sky130_fd_sc_hd__nand2_1 _08501_ (.A(net460),
    .B(\core_pipeline.decode_to_csr_read_address[6] ),
    .Y(_04688_));
 sky130_fd_sc_hd__or3_4 _08502_ (.A(_04686_),
    .B(_04687_),
    .C(_04688_),
    .X(_04689_));
 sky130_fd_sc_hd__nor2_4 _08503_ (.A(_04684_),
    .B(_04689_),
    .Y(_04690_));
 sky130_fd_sc_hd__or4_4 _08504_ (.A(net513),
    .B(\core_pipeline.decode_to_csr_read_address[5] ),
    .C(\core_pipeline.decode_to_csr_read_address[7] ),
    .D(\core_pipeline.decode_to_csr_read_address[6] ),
    .X(_04691_));
 sky130_fd_sc_hd__or3_4 _08505_ (.A(\core_pipeline.decode_to_csr_read_address[10] ),
    .B(\core_pipeline.decode_to_csr_read_address[11] ),
    .C(_04685_),
    .X(_04692_));
 sky130_fd_sc_hd__nor2_4 _08506_ (.A(_04691_),
    .B(_04692_),
    .Y(_04693_));
 sky130_fd_sc_hd__nor2_8 _08507_ (.A(net464),
    .B(net516),
    .Y(_04694_));
 sky130_fd_sc_hd__nor2_8 _08508_ (.A(_03327_),
    .B(net542),
    .Y(_04695_));
 sky130_fd_sc_hd__nand2_1 _08509_ (.A(net370),
    .B(net366),
    .Y(_04696_));
 sky130_fd_sc_hd__and3_4 _08510_ (.A(_04693_),
    .B(net369),
    .C(net366),
    .X(_04697_));
 sky130_fd_sc_hd__nor2_2 _08511_ (.A(_03327_),
    .B(_04682_),
    .Y(_04698_));
 sky130_fd_sc_hd__nand2_8 _08512_ (.A(net430),
    .B(net366),
    .Y(_04699_));
 sky130_fd_sc_hd__nor2_8 _08513_ (.A(_04689_),
    .B(_04699_),
    .Y(_04700_));
 sky130_fd_sc_hd__a22o_1 _08514_ (.A1(\core_pipeline.csr_to_fetch_trap_vector[31] ),
    .A2(net271),
    .B1(net269),
    .B2(\core_pipeline.pipeline_csr.mtimecmp[63] ),
    .X(_04701_));
 sky130_fd_sc_hd__nand2_1 _08515_ (.A(\core_pipeline.decode_to_csr_read_address[10] ),
    .B(\core_pipeline.decode_to_csr_read_address[11] ),
    .Y(_04702_));
 sky130_fd_sc_hd__o31a_1 _08516_ (.A1(\core_pipeline.decode_to_csr_read_address[9] ),
    .A2(\core_pipeline.decode_to_csr_read_address[8] ),
    .A3(_04702_),
    .B1(_04686_),
    .X(_04703_));
 sky130_fd_sc_hd__or2_4 _08517_ (.A(_04691_),
    .B(_04703_),
    .X(_04704_));
 sky130_fd_sc_hd__nor2_8 _08518_ (.A(_04682_),
    .B(_04704_),
    .Y(_04705_));
 sky130_fd_sc_hd__and2_4 _08519_ (.A(net537),
    .B(net430),
    .X(_04706_));
 sky130_fd_sc_hd__nand2_4 _08520_ (.A(_03327_),
    .B(net361),
    .Y(_04707_));
 sky130_fd_sc_hd__nor2_8 _08521_ (.A(_04704_),
    .B(_04707_),
    .Y(_04708_));
 sky130_fd_sc_hd__or4_4 _08522_ (.A(\core_pipeline.decode_to_csr_read_address[5] ),
    .B(\core_pipeline.decode_to_csr_read_address[7] ),
    .C(_04688_),
    .D(_04692_),
    .X(_04709_));
 sky130_fd_sc_hd__nor2_4 _08523_ (.A(_04707_),
    .B(_04709_),
    .Y(_04710_));
 sky130_fd_sc_hd__nor2_4 _08524_ (.A(_04699_),
    .B(_04709_),
    .Y(_04711_));
 sky130_fd_sc_hd__a22o_1 _08525_ (.A1(\core_pipeline.pipeline_csr.minterupt ),
    .A2(_04710_),
    .B1(net267),
    .B2(\core_pipeline.csr_to_fetch_mret_vector[31] ),
    .X(_04712_));
 sky130_fd_sc_hd__a221o_1 _08526_ (.A1(\core_pipeline.pipeline_csr.cycle[31] ),
    .A2(net251),
    .B1(net249),
    .B2(\core_pipeline.pipeline_csr.instret[31] ),
    .C1(_04712_),
    .X(_04713_));
 sky130_fd_sc_hd__a211o_1 _08527_ (.A1(\core_pipeline.pipeline_csr.mtimecmp[31] ),
    .A2(net273),
    .B1(_04701_),
    .C1(_04713_),
    .X(_04714_));
 sky130_fd_sc_hd__or3_4 _08528_ (.A(\core_pipeline.decode_to_csr_read_address[6] ),
    .B(_04687_),
    .C(_04703_),
    .X(_04715_));
 sky130_fd_sc_hd__or2_4 _08529_ (.A(net513),
    .B(_04707_),
    .X(_04716_));
 sky130_fd_sc_hd__nor2_8 _08530_ (.A(_04715_),
    .B(_04716_),
    .Y(_04717_));
 sky130_fd_sc_hd__nor3_2 _08531_ (.A(net513),
    .B(_04682_),
    .C(_04715_),
    .Y(_04718_));
 sky130_fd_sc_hd__nor2_8 _08532_ (.A(_04684_),
    .B(_04709_),
    .Y(_04719_));
 sky130_fd_sc_hd__a22o_1 _08533_ (.A1(\core_pipeline.pipeline_csr.cycle[63] ),
    .A2(net246),
    .B1(net265),
    .B2(\core_pipeline.pipeline_csr.mscratch[31] ),
    .X(_04720_));
 sky130_fd_sc_hd__a211o_1 _08534_ (.A1(\core_pipeline.pipeline_csr.instret[63] ),
    .A2(net247),
    .B1(_04720_),
    .C1(net136),
    .X(_04721_));
 sky130_fd_sc_hd__and4_2 _08535_ (.A(net565),
    .B(_03328_),
    .C(_04693_),
    .D(net370),
    .X(_04722_));
 sky130_fd_sc_hd__or3_4 _08536_ (.A(_04686_),
    .B(_04687_),
    .C(_04688_),
    .X(_04723_));
 sky130_fd_sc_hd__nor2_4 _08537_ (.A(_04699_),
    .B(_04723_),
    .Y(_04724_));
 sky130_fd_sc_hd__nor2_4 _08538_ (.A(_04684_),
    .B(_04723_),
    .Y(_04725_));
 sky130_fd_sc_hd__o22a_1 _08539_ (.A1(\core_pipeline.decode_to_execute_csr_data[31] ),
    .A2(net159),
    .B1(_04714_),
    .B2(_04721_),
    .X(_00400_));
 sky130_fd_sc_hd__and2_4 _08540_ (.A(_04693_),
    .B(net276),
    .X(_04726_));
 sky130_fd_sc_hd__a221o_1 _08541_ (.A1(\core_pipeline.csr_to_fetch_mret_vector[30] ),
    .A2(net267),
    .B1(net246),
    .B2(\core_pipeline.pipeline_csr.cycle[62] ),
    .C1(_04726_),
    .X(_04727_));
 sky130_fd_sc_hd__a221o_1 _08542_ (.A1(\core_pipeline.pipeline_csr.cycle[30] ),
    .A2(net251),
    .B1(net249),
    .B2(\core_pipeline.pipeline_csr.instret[30] ),
    .C1(_04727_),
    .X(_04728_));
 sky130_fd_sc_hd__a22o_1 _08543_ (.A1(\core_pipeline.pipeline_csr.mtimecmp[62] ),
    .A2(net269),
    .B1(net265),
    .B2(\core_pipeline.pipeline_csr.mscratch[30] ),
    .X(_04729_));
 sky130_fd_sc_hd__a221o_1 _08544_ (.A1(\core_pipeline.pipeline_csr.mtimecmp[30] ),
    .A2(net273),
    .B1(net271),
    .B2(\core_pipeline.csr_to_fetch_trap_vector[30] ),
    .C1(_04729_),
    .X(_04730_));
 sky130_fd_sc_hd__a211o_1 _08545_ (.A1(\core_pipeline.pipeline_csr.instret[62] ),
    .A2(net247),
    .B1(_04730_),
    .C1(net136),
    .X(_04731_));
 sky130_fd_sc_hd__o22a_1 _08546_ (.A1(\core_pipeline.decode_to_execute_csr_data[30] ),
    .A2(net159),
    .B1(_04728_),
    .B2(_04731_),
    .X(_00401_));
 sky130_fd_sc_hd__a22o_1 _08547_ (.A1(\core_pipeline.pipeline_csr.cycle[29] ),
    .A2(net251),
    .B1(net246),
    .B2(\core_pipeline.pipeline_csr.cycle[61] ),
    .X(_04732_));
 sky130_fd_sc_hd__a221o_1 _08548_ (.A1(\core_pipeline.pipeline_csr.instret[29] ),
    .A2(net249),
    .B1(net247),
    .B2(\core_pipeline.pipeline_csr.instret[61] ),
    .C1(_04732_),
    .X(_04733_));
 sky130_fd_sc_hd__a22o_1 _08549_ (.A1(\core_pipeline.pipeline_csr.mtimecmp[29] ),
    .A2(net273),
    .B1(net271),
    .B2(\core_pipeline.csr_to_fetch_trap_vector[29] ),
    .X(_04734_));
 sky130_fd_sc_hd__a22o_1 _08550_ (.A1(\core_pipeline.csr_to_fetch_mret_vector[29] ),
    .A2(net267),
    .B1(net265),
    .B2(\core_pipeline.pipeline_csr.mscratch[29] ),
    .X(_04735_));
 sky130_fd_sc_hd__a211o_1 _08551_ (.A1(\core_pipeline.pipeline_csr.mtimecmp[61] ),
    .A2(net269),
    .B1(_04734_),
    .C1(_04735_),
    .X(_04736_));
 sky130_fd_sc_hd__or3_1 _08552_ (.A(net136),
    .B(_04733_),
    .C(_04736_),
    .X(_04737_));
 sky130_fd_sc_hd__o21a_1 _08553_ (.A1(\core_pipeline.decode_to_execute_csr_data[29] ),
    .A2(net159),
    .B1(_04737_),
    .X(_00402_));
 sky130_fd_sc_hd__a22o_1 _08554_ (.A1(\core_pipeline.pipeline_csr.cycle[28] ),
    .A2(net251),
    .B1(net265),
    .B2(\core_pipeline.pipeline_csr.mscratch[28] ),
    .X(_04738_));
 sky130_fd_sc_hd__a221o_1 _08555_ (.A1(\core_pipeline.pipeline_csr.instret[28] ),
    .A2(net249),
    .B1(net246),
    .B2(\core_pipeline.pipeline_csr.cycle[60] ),
    .C1(_04738_),
    .X(_04739_));
 sky130_fd_sc_hd__a22o_1 _08556_ (.A1(\core_pipeline.pipeline_csr.mtimecmp[28] ),
    .A2(net273),
    .B1(net271),
    .B2(\core_pipeline.csr_to_fetch_trap_vector[28] ),
    .X(_04740_));
 sky130_fd_sc_hd__a22o_1 _08557_ (.A1(\core_pipeline.csr_to_fetch_mret_vector[28] ),
    .A2(net267),
    .B1(net247),
    .B2(\core_pipeline.pipeline_csr.instret[60] ),
    .X(_04741_));
 sky130_fd_sc_hd__a211o_1 _08558_ (.A1(\core_pipeline.pipeline_csr.mtimecmp[60] ),
    .A2(net269),
    .B1(_04740_),
    .C1(_04741_),
    .X(_04742_));
 sky130_fd_sc_hd__or3_1 _08559_ (.A(net136),
    .B(_04739_),
    .C(_04742_),
    .X(_04743_));
 sky130_fd_sc_hd__o21a_1 _08560_ (.A1(\core_pipeline.decode_to_execute_csr_data[28] ),
    .A2(net159),
    .B1(_04743_),
    .X(_00403_));
 sky130_fd_sc_hd__a22o_1 _08561_ (.A1(\core_pipeline.csr_to_fetch_mret_vector[27] ),
    .A2(net267),
    .B1(net265),
    .B2(\core_pipeline.pipeline_csr.mscratch[27] ),
    .X(_04744_));
 sky130_fd_sc_hd__a221o_1 _08562_ (.A1(\core_pipeline.pipeline_csr.cycle[27] ),
    .A2(net251),
    .B1(net249),
    .B2(\core_pipeline.pipeline_csr.instret[27] ),
    .C1(_04744_),
    .X(_04745_));
 sky130_fd_sc_hd__a22o_1 _08563_ (.A1(\core_pipeline.pipeline_csr.instret[59] ),
    .A2(net247),
    .B1(net246),
    .B2(\core_pipeline.pipeline_csr.cycle[59] ),
    .X(_04746_));
 sky130_fd_sc_hd__a22o_1 _08564_ (.A1(\core_pipeline.pipeline_csr.mtimecmp[27] ),
    .A2(net273),
    .B1(net271),
    .B2(\core_pipeline.csr_to_fetch_trap_vector[27] ),
    .X(_04747_));
 sky130_fd_sc_hd__a211o_1 _08565_ (.A1(\core_pipeline.pipeline_csr.mtimecmp[59] ),
    .A2(net269),
    .B1(_04746_),
    .C1(_04747_),
    .X(_04748_));
 sky130_fd_sc_hd__or3_1 _08566_ (.A(net136),
    .B(_04745_),
    .C(_04748_),
    .X(_04749_));
 sky130_fd_sc_hd__o21a_1 _08567_ (.A1(\core_pipeline.decode_to_execute_csr_data[27] ),
    .A2(net159),
    .B1(_04749_),
    .X(_00404_));
 sky130_fd_sc_hd__a22o_1 _08568_ (.A1(\core_pipeline.pipeline_csr.cycle[26] ),
    .A2(net251),
    .B1(net247),
    .B2(\core_pipeline.pipeline_csr.instret[58] ),
    .X(_04750_));
 sky130_fd_sc_hd__a221o_1 _08569_ (.A1(\core_pipeline.pipeline_csr.instret[26] ),
    .A2(net249),
    .B1(net246),
    .B2(\core_pipeline.pipeline_csr.cycle[58] ),
    .C1(_04750_),
    .X(_04751_));
 sky130_fd_sc_hd__a22o_1 _08570_ (.A1(\core_pipeline.pipeline_csr.mtimecmp[26] ),
    .A2(net273),
    .B1(net271),
    .B2(\core_pipeline.csr_to_fetch_trap_vector[26] ),
    .X(_04752_));
 sky130_fd_sc_hd__a22o_1 _08571_ (.A1(\core_pipeline.csr_to_fetch_mret_vector[26] ),
    .A2(net267),
    .B1(net265),
    .B2(\core_pipeline.pipeline_csr.mscratch[26] ),
    .X(_04753_));
 sky130_fd_sc_hd__a2111o_1 _08572_ (.A1(\core_pipeline.pipeline_csr.mtimecmp[58] ),
    .A2(net269),
    .B1(_04751_),
    .C1(_04752_),
    .D1(_04753_),
    .X(_04754_));
 sky130_fd_sc_hd__mux2_1 _08573_ (.A0(\core_pipeline.decode_to_execute_csr_data[26] ),
    .A1(_04754_),
    .S(net159),
    .X(_00405_));
 sky130_fd_sc_hd__a22o_1 _08574_ (.A1(\core_pipeline.pipeline_csr.cycle[25] ),
    .A2(net251),
    .B1(net249),
    .B2(\core_pipeline.pipeline_csr.instret[25] ),
    .X(_04755_));
 sky130_fd_sc_hd__a221o_1 _08575_ (.A1(\core_pipeline.csr_to_fetch_mret_vector[25] ),
    .A2(net267),
    .B1(net248),
    .B2(\core_pipeline.pipeline_csr.instret[57] ),
    .C1(_04755_),
    .X(_04756_));
 sky130_fd_sc_hd__a22o_1 _08576_ (.A1(\core_pipeline.pipeline_csr.mtimecmp[25] ),
    .A2(net273),
    .B1(net271),
    .B2(\core_pipeline.csr_to_fetch_trap_vector[25] ),
    .X(_04757_));
 sky130_fd_sc_hd__a22o_1 _08577_ (.A1(\core_pipeline.pipeline_csr.cycle[57] ),
    .A2(net246),
    .B1(net266),
    .B2(\core_pipeline.pipeline_csr.mscratch[25] ),
    .X(_04758_));
 sky130_fd_sc_hd__a211o_1 _08578_ (.A1(\core_pipeline.pipeline_csr.mtimecmp[57] ),
    .A2(net269),
    .B1(_04757_),
    .C1(_04758_),
    .X(_04759_));
 sky130_fd_sc_hd__or3_1 _08579_ (.A(net136),
    .B(_04756_),
    .C(_04759_),
    .X(_04760_));
 sky130_fd_sc_hd__o21a_1 _08580_ (.A1(\core_pipeline.decode_to_execute_csr_data[25] ),
    .A2(net162),
    .B1(_04760_),
    .X(_00406_));
 sky130_fd_sc_hd__a22o_1 _08581_ (.A1(\core_pipeline.pipeline_csr.cycle[24] ),
    .A2(net251),
    .B1(net266),
    .B2(\core_pipeline.pipeline_csr.mscratch[24] ),
    .X(_04761_));
 sky130_fd_sc_hd__a221o_1 _08582_ (.A1(\core_pipeline.pipeline_csr.instret[24] ),
    .A2(net249),
    .B1(net245),
    .B2(\core_pipeline.pipeline_csr.cycle[56] ),
    .C1(_04761_),
    .X(_04762_));
 sky130_fd_sc_hd__a22o_1 _08583_ (.A1(\core_pipeline.pipeline_csr.mtimecmp[24] ),
    .A2(net274),
    .B1(net272),
    .B2(\core_pipeline.csr_to_fetch_trap_vector[24] ),
    .X(_04763_));
 sky130_fd_sc_hd__a22o_1 _08584_ (.A1(\core_pipeline.csr_to_fetch_mret_vector[24] ),
    .A2(net268),
    .B1(net247),
    .B2(\core_pipeline.pipeline_csr.instret[56] ),
    .X(_04764_));
 sky130_fd_sc_hd__a2111o_1 _08585_ (.A1(\core_pipeline.pipeline_csr.mtimecmp[56] ),
    .A2(net270),
    .B1(_04762_),
    .C1(_04763_),
    .D1(_04764_),
    .X(_04765_));
 sky130_fd_sc_hd__mux2_1 _08586_ (.A0(\core_pipeline.decode_to_execute_csr_data[24] ),
    .A1(_04765_),
    .S(net162),
    .X(_00407_));
 sky130_fd_sc_hd__a22o_1 _08587_ (.A1(\core_pipeline.pipeline_csr.cycle[23] ),
    .A2(net252),
    .B1(net268),
    .B2(\core_pipeline.csr_to_fetch_mret_vector[23] ),
    .X(_04766_));
 sky130_fd_sc_hd__a221o_1 _08588_ (.A1(\core_pipeline.pipeline_csr.instret[23] ),
    .A2(net250),
    .B1(net266),
    .B2(\core_pipeline.pipeline_csr.mscratch[23] ),
    .C1(_04766_),
    .X(_04767_));
 sky130_fd_sc_hd__a22o_1 _08589_ (.A1(\core_pipeline.pipeline_csr.mtimecmp[23] ),
    .A2(net274),
    .B1(net272),
    .B2(\core_pipeline.csr_to_fetch_trap_vector[23] ),
    .X(_04768_));
 sky130_fd_sc_hd__a22o_1 _08590_ (.A1(\core_pipeline.pipeline_csr.instret[55] ),
    .A2(net247),
    .B1(net245),
    .B2(\core_pipeline.pipeline_csr.cycle[55] ),
    .X(_04769_));
 sky130_fd_sc_hd__a2111o_1 _08591_ (.A1(\core_pipeline.pipeline_csr.mtimecmp[55] ),
    .A2(net270),
    .B1(_04767_),
    .C1(_04768_),
    .D1(_04769_),
    .X(_04770_));
 sky130_fd_sc_hd__mux2_1 _08592_ (.A0(\core_pipeline.decode_to_execute_csr_data[23] ),
    .A1(_04770_),
    .S(net162),
    .X(_00408_));
 sky130_fd_sc_hd__a22o_1 _08593_ (.A1(\core_pipeline.pipeline_csr.cycle[22] ),
    .A2(net252),
    .B1(net265),
    .B2(\core_pipeline.pipeline_csr.mscratch[22] ),
    .X(_04771_));
 sky130_fd_sc_hd__a221o_1 _08594_ (.A1(\core_pipeline.pipeline_csr.instret[22] ),
    .A2(net250),
    .B1(net245),
    .B2(\core_pipeline.pipeline_csr.cycle[54] ),
    .C1(_04771_),
    .X(_04772_));
 sky130_fd_sc_hd__a22o_1 _08595_ (.A1(\core_pipeline.pipeline_csr.mtimecmp[22] ),
    .A2(net273),
    .B1(net271),
    .B2(\core_pipeline.csr_to_fetch_trap_vector[22] ),
    .X(_04773_));
 sky130_fd_sc_hd__a22o_1 _08596_ (.A1(\core_pipeline.csr_to_fetch_mret_vector[22] ),
    .A2(net267),
    .B1(net248),
    .B2(\core_pipeline.pipeline_csr.instret[54] ),
    .X(_04774_));
 sky130_fd_sc_hd__a211o_1 _08597_ (.A1(\core_pipeline.pipeline_csr.mtimecmp[54] ),
    .A2(net269),
    .B1(_04773_),
    .C1(_04774_),
    .X(_04775_));
 sky130_fd_sc_hd__or3_1 _08598_ (.A(net136),
    .B(_04772_),
    .C(_04775_),
    .X(_04776_));
 sky130_fd_sc_hd__o21a_1 _08599_ (.A1(\core_pipeline.decode_to_execute_csr_data[22] ),
    .A2(net162),
    .B1(_04776_),
    .X(_00409_));
 sky130_fd_sc_hd__a22o_1 _08600_ (.A1(\core_pipeline.pipeline_csr.cycle[21] ),
    .A2(net252),
    .B1(net245),
    .B2(\core_pipeline.pipeline_csr.cycle[53] ),
    .X(_04777_));
 sky130_fd_sc_hd__a221o_1 _08601_ (.A1(\core_pipeline.pipeline_csr.instret[21] ),
    .A2(net250),
    .B1(net265),
    .B2(\core_pipeline.pipeline_csr.mscratch[21] ),
    .C1(_04777_),
    .X(_04778_));
 sky130_fd_sc_hd__a22o_1 _08602_ (.A1(\core_pipeline.pipeline_csr.mtimecmp[21] ),
    .A2(net273),
    .B1(net271),
    .B2(\core_pipeline.csr_to_fetch_trap_vector[21] ),
    .X(_04779_));
 sky130_fd_sc_hd__a22o_1 _08603_ (.A1(\core_pipeline.csr_to_fetch_mret_vector[21] ),
    .A2(net268),
    .B1(net248),
    .B2(\core_pipeline.pipeline_csr.instret[53] ),
    .X(_04780_));
 sky130_fd_sc_hd__a211o_1 _08604_ (.A1(\core_pipeline.pipeline_csr.mtimecmp[53] ),
    .A2(net269),
    .B1(_04779_),
    .C1(_04780_),
    .X(_04781_));
 sky130_fd_sc_hd__or3_1 _08605_ (.A(net136),
    .B(_04778_),
    .C(_04781_),
    .X(_04782_));
 sky130_fd_sc_hd__o21a_1 _08606_ (.A1(\core_pipeline.decode_to_execute_csr_data[21] ),
    .A2(net162),
    .B1(_04782_),
    .X(_00410_));
 sky130_fd_sc_hd__a22o_1 _08607_ (.A1(\core_pipeline.pipeline_csr.cycle[20] ),
    .A2(net252),
    .B1(net250),
    .B2(\core_pipeline.pipeline_csr.instret[20] ),
    .X(_04783_));
 sky130_fd_sc_hd__a221o_1 _08608_ (.A1(\core_pipeline.csr_to_fetch_mret_vector[20] ),
    .A2(net268),
    .B1(net248),
    .B2(\core_pipeline.pipeline_csr.instret[52] ),
    .C1(_04783_),
    .X(_04784_));
 sky130_fd_sc_hd__a22o_1 _08609_ (.A1(\core_pipeline.pipeline_csr.mtimecmp[20] ),
    .A2(net273),
    .B1(net271),
    .B2(\core_pipeline.csr_to_fetch_trap_vector[20] ),
    .X(_04785_));
 sky130_fd_sc_hd__a22o_1 _08610_ (.A1(\core_pipeline.pipeline_csr.cycle[52] ),
    .A2(net245),
    .B1(net266),
    .B2(\core_pipeline.pipeline_csr.mscratch[20] ),
    .X(_04786_));
 sky130_fd_sc_hd__a211o_1 _08611_ (.A1(\core_pipeline.pipeline_csr.mtimecmp[52] ),
    .A2(net269),
    .B1(_04785_),
    .C1(_04786_),
    .X(_04787_));
 sky130_fd_sc_hd__or3_2 _08612_ (.A(net136),
    .B(_04784_),
    .C(_04787_),
    .X(_04788_));
 sky130_fd_sc_hd__o21a_1 _08613_ (.A1(\core_pipeline.decode_to_execute_csr_data[20] ),
    .A2(net162),
    .B1(_04788_),
    .X(_00411_));
 sky130_fd_sc_hd__a22o_1 _08614_ (.A1(\core_pipeline.pipeline_csr.instret[19] ),
    .A2(net250),
    .B1(net268),
    .B2(\core_pipeline.csr_to_fetch_mret_vector[19] ),
    .X(_04789_));
 sky130_fd_sc_hd__a221o_1 _08615_ (.A1(\core_pipeline.pipeline_csr.cycle[19] ),
    .A2(net252),
    .B1(net266),
    .B2(\core_pipeline.pipeline_csr.mscratch[19] ),
    .C1(_04789_),
    .X(_04790_));
 sky130_fd_sc_hd__a22o_1 _08616_ (.A1(\core_pipeline.pipeline_csr.instret[51] ),
    .A2(net248),
    .B1(net245),
    .B2(\core_pipeline.pipeline_csr.cycle[51] ),
    .X(_04791_));
 sky130_fd_sc_hd__a22o_1 _08617_ (.A1(\core_pipeline.pipeline_csr.mtimecmp[19] ),
    .A2(net273),
    .B1(net271),
    .B2(\core_pipeline.csr_to_fetch_trap_vector[19] ),
    .X(_04792_));
 sky130_fd_sc_hd__a211o_1 _08618_ (.A1(\core_pipeline.pipeline_csr.mtimecmp[51] ),
    .A2(net269),
    .B1(_04791_),
    .C1(_04792_),
    .X(_04793_));
 sky130_fd_sc_hd__or3_1 _08619_ (.A(net136),
    .B(_04790_),
    .C(_04793_),
    .X(_04794_));
 sky130_fd_sc_hd__o21a_1 _08620_ (.A1(\core_pipeline.decode_to_execute_csr_data[19] ),
    .A2(net162),
    .B1(_04794_),
    .X(_00412_));
 sky130_fd_sc_hd__a22o_1 _08621_ (.A1(\core_pipeline.pipeline_csr.instret[18] ),
    .A2(net250),
    .B1(net266),
    .B2(\core_pipeline.pipeline_csr.mscratch[18] ),
    .X(_04795_));
 sky130_fd_sc_hd__a221o_1 _08622_ (.A1(\core_pipeline.pipeline_csr.cycle[18] ),
    .A2(net252),
    .B1(net268),
    .B2(\core_pipeline.csr_to_fetch_mret_vector[18] ),
    .C1(_04795_),
    .X(_04796_));
 sky130_fd_sc_hd__a22o_1 _08623_ (.A1(\core_pipeline.pipeline_csr.instret[50] ),
    .A2(net248),
    .B1(net245),
    .B2(\core_pipeline.pipeline_csr.cycle[50] ),
    .X(_04797_));
 sky130_fd_sc_hd__a22o_1 _08624_ (.A1(\core_pipeline.csr_to_fetch_trap_vector[18] ),
    .A2(net271),
    .B1(net269),
    .B2(\core_pipeline.pipeline_csr.mtimecmp[50] ),
    .X(_04798_));
 sky130_fd_sc_hd__a2111o_2 _08625_ (.A1(\core_pipeline.pipeline_csr.mtimecmp[18] ),
    .A2(net273),
    .B1(_04796_),
    .C1(_04797_),
    .D1(_04798_),
    .X(_04799_));
 sky130_fd_sc_hd__mux2_1 _08626_ (.A0(\core_pipeline.decode_to_execute_csr_data[18] ),
    .A1(_04799_),
    .S(net162),
    .X(_00413_));
 sky130_fd_sc_hd__a22o_1 _08627_ (.A1(\core_pipeline.pipeline_csr.cycle[17] ),
    .A2(net252),
    .B1(net250),
    .B2(\core_pipeline.pipeline_csr.instret[17] ),
    .X(_04800_));
 sky130_fd_sc_hd__a221o_1 _08628_ (.A1(\core_pipeline.csr_to_fetch_mret_vector[17] ),
    .A2(net268),
    .B1(net248),
    .B2(\core_pipeline.pipeline_csr.instret[49] ),
    .C1(_04800_),
    .X(_04801_));
 sky130_fd_sc_hd__a22o_1 _08629_ (.A1(\core_pipeline.pipeline_csr.mtimecmp[17] ),
    .A2(net274),
    .B1(net271),
    .B2(\core_pipeline.csr_to_fetch_trap_vector[17] ),
    .X(_04802_));
 sky130_fd_sc_hd__a22o_1 _08630_ (.A1(\core_pipeline.pipeline_csr.cycle[49] ),
    .A2(net245),
    .B1(net266),
    .B2(\core_pipeline.pipeline_csr.mscratch[17] ),
    .X(_04803_));
 sky130_fd_sc_hd__a211o_1 _08631_ (.A1(\core_pipeline.pipeline_csr.mtimecmp[49] ),
    .A2(net270),
    .B1(_04802_),
    .C1(_04803_),
    .X(_04804_));
 sky130_fd_sc_hd__or3_1 _08632_ (.A(net136),
    .B(_04801_),
    .C(_04804_),
    .X(_04805_));
 sky130_fd_sc_hd__o21a_1 _08633_ (.A1(\core_pipeline.decode_to_execute_csr_data[17] ),
    .A2(net162),
    .B1(_04805_),
    .X(_00414_));
 sky130_fd_sc_hd__a22o_1 _08634_ (.A1(\core_pipeline.csr_to_fetch_mret_vector[16] ),
    .A2(net268),
    .B1(net266),
    .B2(\core_pipeline.pipeline_csr.mscratch[16] ),
    .X(_04806_));
 sky130_fd_sc_hd__a221o_1 _08635_ (.A1(\core_pipeline.pipeline_csr.cycle[16] ),
    .A2(net252),
    .B1(net250),
    .B2(\core_pipeline.pipeline_csr.instret[16] ),
    .C1(_04806_),
    .X(_04807_));
 sky130_fd_sc_hd__a22o_1 _08636_ (.A1(\core_pipeline.pipeline_csr.instret[48] ),
    .A2(net248),
    .B1(net245),
    .B2(\core_pipeline.pipeline_csr.cycle[48] ),
    .X(_04808_));
 sky130_fd_sc_hd__a22o_1 _08637_ (.A1(\core_pipeline.pipeline_csr.mtimecmp[16] ),
    .A2(net274),
    .B1(net272),
    .B2(\core_pipeline.csr_to_fetch_trap_vector[16] ),
    .X(_04809_));
 sky130_fd_sc_hd__a2111o_4 _08638_ (.A1(\core_pipeline.pipeline_csr.mtimecmp[48] ),
    .A2(net270),
    .B1(_04807_),
    .C1(_04808_),
    .D1(_04809_),
    .X(_04810_));
 sky130_fd_sc_hd__mux2_1 _08639_ (.A0(\core_pipeline.decode_to_execute_csr_data[16] ),
    .A1(_04810_),
    .S(net153),
    .X(_00415_));
 sky130_fd_sc_hd__a22o_1 _08640_ (.A1(\core_pipeline.pipeline_csr.cycle[15] ),
    .A2(net252),
    .B1(net268),
    .B2(\core_pipeline.csr_to_fetch_mret_vector[15] ),
    .X(_04811_));
 sky130_fd_sc_hd__a221o_1 _08641_ (.A1(\core_pipeline.pipeline_csr.instret[15] ),
    .A2(net250),
    .B1(net245),
    .B2(\core_pipeline.pipeline_csr.cycle[47] ),
    .C1(_04811_),
    .X(_04812_));
 sky130_fd_sc_hd__a22o_1 _08642_ (.A1(\core_pipeline.csr_to_fetch_trap_vector[15] ),
    .A2(net272),
    .B1(net270),
    .B2(\core_pipeline.pipeline_csr.mtimecmp[47] ),
    .X(_04813_));
 sky130_fd_sc_hd__a22o_1 _08643_ (.A1(\core_pipeline.pipeline_csr.instret[47] ),
    .A2(net248),
    .B1(net266),
    .B2(\core_pipeline.pipeline_csr.mscratch[15] ),
    .X(_04814_));
 sky130_fd_sc_hd__a211o_1 _08644_ (.A1(\core_pipeline.pipeline_csr.mtimecmp[15] ),
    .A2(net274),
    .B1(_04813_),
    .C1(_04814_),
    .X(_04815_));
 sky130_fd_sc_hd__or3_4 _08645_ (.A(net136),
    .B(_04812_),
    .C(_04815_),
    .X(_04816_));
 sky130_fd_sc_hd__o21a_1 _08646_ (.A1(\core_pipeline.decode_to_execute_csr_data[15] ),
    .A2(net153),
    .B1(_04816_),
    .X(_00416_));
 sky130_fd_sc_hd__a22o_1 _08647_ (.A1(\core_pipeline.pipeline_csr.cycle[14] ),
    .A2(net252),
    .B1(net250),
    .B2(\core_pipeline.pipeline_csr.instret[14] ),
    .X(_04817_));
 sky130_fd_sc_hd__a221o_1 _08648_ (.A1(\core_pipeline.csr_to_fetch_mret_vector[14] ),
    .A2(net268),
    .B1(net248),
    .B2(\core_pipeline.pipeline_csr.instret[46] ),
    .C1(_04817_),
    .X(_04818_));
 sky130_fd_sc_hd__a22o_1 _08649_ (.A1(\core_pipeline.pipeline_csr.mtimecmp[14] ),
    .A2(net274),
    .B1(net272),
    .B2(\core_pipeline.csr_to_fetch_trap_vector[14] ),
    .X(_04819_));
 sky130_fd_sc_hd__a22o_1 _08650_ (.A1(\core_pipeline.pipeline_csr.cycle[46] ),
    .A2(net245),
    .B1(net266),
    .B2(\core_pipeline.pipeline_csr.mscratch[14] ),
    .X(_04820_));
 sky130_fd_sc_hd__a211o_1 _08651_ (.A1(\core_pipeline.pipeline_csr.mtimecmp[46] ),
    .A2(net270),
    .B1(_04819_),
    .C1(_04820_),
    .X(_04821_));
 sky130_fd_sc_hd__or3_4 _08652_ (.A(net137),
    .B(_04818_),
    .C(_04821_),
    .X(_04822_));
 sky130_fd_sc_hd__o21a_1 _08653_ (.A1(\core_pipeline.decode_to_execute_csr_data[14] ),
    .A2(net153),
    .B1(_04822_),
    .X(_00417_));
 sky130_fd_sc_hd__a22o_1 _08654_ (.A1(\core_pipeline.pipeline_csr.cycle[13] ),
    .A2(net252),
    .B1(net250),
    .B2(\core_pipeline.pipeline_csr.instret[13] ),
    .X(_04823_));
 sky130_fd_sc_hd__a221o_1 _08655_ (.A1(\core_pipeline.csr_to_fetch_mret_vector[13] ),
    .A2(net268),
    .B1(net248),
    .B2(\core_pipeline.pipeline_csr.instret[45] ),
    .C1(_04823_),
    .X(_04824_));
 sky130_fd_sc_hd__a22o_1 _08656_ (.A1(\core_pipeline.csr_to_fetch_trap_vector[13] ),
    .A2(net272),
    .B1(net270),
    .B2(\core_pipeline.pipeline_csr.mtimecmp[45] ),
    .X(_04825_));
 sky130_fd_sc_hd__a22o_1 _08657_ (.A1(\core_pipeline.pipeline_csr.cycle[45] ),
    .A2(net245),
    .B1(net266),
    .B2(\core_pipeline.pipeline_csr.mscratch[13] ),
    .X(_04826_));
 sky130_fd_sc_hd__a211o_1 _08658_ (.A1(\core_pipeline.pipeline_csr.mtimecmp[13] ),
    .A2(net274),
    .B1(_04825_),
    .C1(_04826_),
    .X(_04827_));
 sky130_fd_sc_hd__or3_4 _08659_ (.A(net136),
    .B(_04824_),
    .C(_04827_),
    .X(_04828_));
 sky130_fd_sc_hd__o21a_1 _08660_ (.A1(\core_pipeline.decode_to_execute_csr_data[13] ),
    .A2(net153),
    .B1(_04828_),
    .X(_00418_));
 sky130_fd_sc_hd__a22o_1 _08661_ (.A1(\core_pipeline.pipeline_csr.instret[12] ),
    .A2(net250),
    .B1(net248),
    .B2(\core_pipeline.pipeline_csr.instret[44] ),
    .X(_04829_));
 sky130_fd_sc_hd__a221o_1 _08662_ (.A1(\core_pipeline.pipeline_csr.cycle[12] ),
    .A2(net252),
    .B1(net245),
    .B2(\core_pipeline.pipeline_csr.cycle[44] ),
    .C1(_04829_),
    .X(_04830_));
 sky130_fd_sc_hd__a22o_1 _08663_ (.A1(\core_pipeline.pipeline_csr.mtimecmp[12] ),
    .A2(net274),
    .B1(net272),
    .B2(\core_pipeline.csr_to_fetch_trap_vector[12] ),
    .X(_04831_));
 sky130_fd_sc_hd__a22o_1 _08664_ (.A1(\core_pipeline.csr_to_fetch_mret_vector[12] ),
    .A2(net268),
    .B1(net266),
    .B2(\core_pipeline.pipeline_csr.mscratch[12] ),
    .X(_04832_));
 sky130_fd_sc_hd__a2111o_4 _08665_ (.A1(\core_pipeline.pipeline_csr.mtimecmp[44] ),
    .A2(net270),
    .B1(_04830_),
    .C1(_04831_),
    .D1(_04832_),
    .X(_04833_));
 sky130_fd_sc_hd__mux2_1 _08666_ (.A0(\core_pipeline.decode_to_execute_csr_data[12] ),
    .A1(_04833_),
    .S(net153),
    .X(_00419_));
 sky130_fd_sc_hd__and3_2 _08667_ (.A(net427),
    .B(_04693_),
    .C(net370),
    .X(_04834_));
 sky130_fd_sc_hd__and4b_4 _08668_ (.A_N(_04709_),
    .B(_03328_),
    .C(_03327_),
    .D(net370),
    .X(_04835_));
 sky130_fd_sc_hd__a22o_1 _08669_ (.A1(\core_pipeline.pipeline_csr.cycle[11] ),
    .A2(net252),
    .B1(net248),
    .B2(\core_pipeline.pipeline_csr.instret[43] ),
    .X(_04836_));
 sky130_fd_sc_hd__a221o_2 _08670_ (.A1(\core_pipeline.pipeline_csr.instret[11] ),
    .A2(net250),
    .B1(net245),
    .B2(\core_pipeline.pipeline_csr.cycle[43] ),
    .C1(_04836_),
    .X(_04837_));
 sky130_fd_sc_hd__a22o_1 _08671_ (.A1(\core_pipeline.pipeline_csr.mscratch[11] ),
    .A2(net265),
    .B1(_04722_),
    .B2(\core_pipeline.csr_to_fetch_trap_vector[11] ),
    .X(_04838_));
 sky130_fd_sc_hd__a22o_1 _08672_ (.A1(\core_pipeline.csr_to_fetch_mret_vector[11] ),
    .A2(net267),
    .B1(_04835_),
    .B2(net34),
    .X(_04839_));
 sky130_fd_sc_hd__a221o_1 _08673_ (.A1(\core_pipeline.pipeline_csr.mtimecmp[43] ),
    .A2(_04724_),
    .B1(_04725_),
    .B2(\core_pipeline.pipeline_csr.mtimecmp[11] ),
    .C1(_04839_),
    .X(_04840_));
 sky130_fd_sc_hd__a2111o_1 _08674_ (.A1(\core_pipeline.pipeline_csr.meie ),
    .A2(_04834_),
    .B1(_04838_),
    .C1(_04840_),
    .D1(net136),
    .X(_04841_));
 sky130_fd_sc_hd__o22a_1 _08675_ (.A1(\core_pipeline.decode_to_execute_csr_data[11] ),
    .A2(net159),
    .B1(_04837_),
    .B2(_04841_),
    .X(_00420_));
 sky130_fd_sc_hd__a22o_1 _08676_ (.A1(\core_pipeline.pipeline_csr.cycle[10] ),
    .A2(net252),
    .B1(net245),
    .B2(\core_pipeline.pipeline_csr.cycle[42] ),
    .X(_04842_));
 sky130_fd_sc_hd__a221o_1 _08677_ (.A1(\core_pipeline.pipeline_csr.instret[10] ),
    .A2(net250),
    .B1(net248),
    .B2(\core_pipeline.pipeline_csr.instret[42] ),
    .C1(_04842_),
    .X(_04843_));
 sky130_fd_sc_hd__a22o_1 _08678_ (.A1(\core_pipeline.csr_to_fetch_trap_vector[10] ),
    .A2(net272),
    .B1(net270),
    .B2(\core_pipeline.pipeline_csr.mtimecmp[42] ),
    .X(_04844_));
 sky130_fd_sc_hd__a22o_1 _08679_ (.A1(\core_pipeline.csr_to_fetch_mret_vector[10] ),
    .A2(net268),
    .B1(net266),
    .B2(\core_pipeline.pipeline_csr.mscratch[10] ),
    .X(_04845_));
 sky130_fd_sc_hd__a211o_1 _08680_ (.A1(\core_pipeline.pipeline_csr.mtimecmp[10] ),
    .A2(net274),
    .B1(_04844_),
    .C1(_04845_),
    .X(_04846_));
 sky130_fd_sc_hd__or3_4 _08681_ (.A(net137),
    .B(_04843_),
    .C(_04846_),
    .X(_04847_));
 sky130_fd_sc_hd__o21a_1 _08682_ (.A1(\core_pipeline.decode_to_execute_csr_data[10] ),
    .A2(net155),
    .B1(_04847_),
    .X(_00421_));
 sky130_fd_sc_hd__a22o_1 _08683_ (.A1(\core_pipeline.pipeline_csr.instret[9] ),
    .A2(net250),
    .B1(net268),
    .B2(\core_pipeline.csr_to_fetch_mret_vector[9] ),
    .X(_04848_));
 sky130_fd_sc_hd__a221o_1 _08684_ (.A1(\core_pipeline.pipeline_csr.cycle[9] ),
    .A2(net252),
    .B1(net266),
    .B2(\core_pipeline.pipeline_csr.mscratch[9] ),
    .C1(_04848_),
    .X(_04849_));
 sky130_fd_sc_hd__a22o_1 _08685_ (.A1(\core_pipeline.pipeline_csr.instret[41] ),
    .A2(net248),
    .B1(net245),
    .B2(\core_pipeline.pipeline_csr.cycle[41] ),
    .X(_04850_));
 sky130_fd_sc_hd__a22o_1 _08686_ (.A1(\core_pipeline.pipeline_csr.mtimecmp[9] ),
    .A2(net274),
    .B1(net272),
    .B2(\core_pipeline.csr_to_fetch_trap_vector[9] ),
    .X(_04851_));
 sky130_fd_sc_hd__a211o_1 _08687_ (.A1(\core_pipeline.pipeline_csr.mtimecmp[41] ),
    .A2(net270),
    .B1(_04850_),
    .C1(_04851_),
    .X(_04852_));
 sky130_fd_sc_hd__or3_4 _08688_ (.A(net137),
    .B(_04849_),
    .C(_04852_),
    .X(_04853_));
 sky130_fd_sc_hd__o21a_1 _08689_ (.A1(\core_pipeline.decode_to_execute_csr_data[9] ),
    .A2(net155),
    .B1(_04853_),
    .X(_00422_));
 sky130_fd_sc_hd__a22o_1 _08690_ (.A1(\core_pipeline.pipeline_csr.mtimecmp[8] ),
    .A2(net274),
    .B1(net272),
    .B2(\core_pipeline.csr_to_fetch_trap_vector[8] ),
    .X(_04854_));
 sky130_fd_sc_hd__a221o_1 _08691_ (.A1(\core_pipeline.csr_to_fetch_mret_vector[8] ),
    .A2(net268),
    .B1(net245),
    .B2(\core_pipeline.pipeline_csr.cycle[40] ),
    .C1(_04726_),
    .X(_04855_));
 sky130_fd_sc_hd__a221o_1 _08692_ (.A1(\core_pipeline.pipeline_csr.cycle[8] ),
    .A2(net251),
    .B1(net249),
    .B2(\core_pipeline.pipeline_csr.instret[8] ),
    .C1(_04855_),
    .X(_04856_));
 sky130_fd_sc_hd__a221o_1 _08693_ (.A1(\core_pipeline.pipeline_csr.mtimecmp[40] ),
    .A2(net270),
    .B1(net266),
    .B2(\core_pipeline.pipeline_csr.mscratch[8] ),
    .C1(_04854_),
    .X(_04857_));
 sky130_fd_sc_hd__a211o_1 _08694_ (.A1(\core_pipeline.pipeline_csr.instret[40] ),
    .A2(net247),
    .B1(_04857_),
    .C1(net136),
    .X(_04858_));
 sky130_fd_sc_hd__o22a_1 _08695_ (.A1(\core_pipeline.decode_to_execute_csr_data[8] ),
    .A2(net159),
    .B1(_04856_),
    .B2(_04858_),
    .X(_00423_));
 sky130_fd_sc_hd__a22o_1 _08696_ (.A1(\core_pipeline.pipeline_csr.instret[39] ),
    .A2(net247),
    .B1(net246),
    .B2(\core_pipeline.pipeline_csr.cycle[39] ),
    .X(_04859_));
 sky130_fd_sc_hd__and3_1 _08697_ (.A(\core_pipeline.pipeline_csr.pie ),
    .B(_04683_),
    .C(_04693_),
    .X(_04860_));
 sky130_fd_sc_hd__a221o_1 _08698_ (.A1(\core_pipeline.pipeline_csr.cycle[7] ),
    .A2(net251),
    .B1(net249),
    .B2(\core_pipeline.pipeline_csr.instret[7] ),
    .C1(_04859_),
    .X(_04861_));
 sky130_fd_sc_hd__a22o_1 _08699_ (.A1(\core_pipeline.csr_to_fetch_mret_vector[7] ),
    .A2(net267),
    .B1(_04724_),
    .B2(\core_pipeline.pipeline_csr.mtimecmp[39] ),
    .X(_04862_));
 sky130_fd_sc_hd__a221o_1 _08700_ (.A1(\core_pipeline.pipeline_csr.mscratch[7] ),
    .A2(net265),
    .B1(_04725_),
    .B2(\core_pipeline.pipeline_csr.mtimecmp[7] ),
    .C1(_04860_),
    .X(_04863_));
 sky130_fd_sc_hd__a221o_1 _08701_ (.A1(\core_pipeline.pipeline_csr.mtie ),
    .A2(_04834_),
    .B1(_04835_),
    .B2(\core_pipeline.pipeline_csr.mtip ),
    .C1(_04863_),
    .X(_04864_));
 sky130_fd_sc_hd__a2111o_1 _08702_ (.A1(\core_pipeline.csr_to_fetch_trap_vector[7] ),
    .A2(_04722_),
    .B1(_04862_),
    .C1(_04864_),
    .D1(net137),
    .X(_04865_));
 sky130_fd_sc_hd__o22a_1 _08703_ (.A1(\core_pipeline.decode_to_execute_csr_data[7] ),
    .A2(net157),
    .B1(_04861_),
    .B2(_04865_),
    .X(_00424_));
 sky130_fd_sc_hd__a22o_1 _08704_ (.A1(\core_pipeline.pipeline_csr.cycle[6] ),
    .A2(net251),
    .B1(net249),
    .B2(\core_pipeline.pipeline_csr.instret[6] ),
    .X(_04866_));
 sky130_fd_sc_hd__a221o_1 _08705_ (.A1(\core_pipeline.csr_to_fetch_mret_vector[6] ),
    .A2(net267),
    .B1(net247),
    .B2(\core_pipeline.pipeline_csr.instret[38] ),
    .C1(_04866_),
    .X(_04867_));
 sky130_fd_sc_hd__a22o_1 _08706_ (.A1(\core_pipeline.pipeline_csr.mtimecmp[6] ),
    .A2(net273),
    .B1(net271),
    .B2(\core_pipeline.csr_to_fetch_trap_vector[6] ),
    .X(_04868_));
 sky130_fd_sc_hd__a22o_1 _08707_ (.A1(\core_pipeline.pipeline_csr.cycle[38] ),
    .A2(net246),
    .B1(net265),
    .B2(\core_pipeline.pipeline_csr.mscratch[6] ),
    .X(_04869_));
 sky130_fd_sc_hd__a211o_1 _08708_ (.A1(\core_pipeline.pipeline_csr.mtimecmp[38] ),
    .A2(net269),
    .B1(_04868_),
    .C1(_04869_),
    .X(_04870_));
 sky130_fd_sc_hd__or3_4 _08709_ (.A(net136),
    .B(_04867_),
    .C(_04870_),
    .X(_04871_));
 sky130_fd_sc_hd__o21a_1 _08710_ (.A1(\core_pipeline.decode_to_execute_csr_data[6] ),
    .A2(net150),
    .B1(_04871_),
    .X(_00425_));
 sky130_fd_sc_hd__a22o_1 _08711_ (.A1(\core_pipeline.pipeline_csr.instret[5] ),
    .A2(net249),
    .B1(net265),
    .B2(\core_pipeline.pipeline_csr.mscratch[5] ),
    .X(_04872_));
 sky130_fd_sc_hd__a221o_1 _08712_ (.A1(\core_pipeline.pipeline_csr.cycle[5] ),
    .A2(net251),
    .B1(net246),
    .B2(\core_pipeline.pipeline_csr.cycle[37] ),
    .C1(_04872_),
    .X(_04873_));
 sky130_fd_sc_hd__a22o_1 _08713_ (.A1(\core_pipeline.pipeline_csr.mtimecmp[5] ),
    .A2(net273),
    .B1(net271),
    .B2(\core_pipeline.csr_to_fetch_trap_vector[5] ),
    .X(_04874_));
 sky130_fd_sc_hd__a22o_1 _08714_ (.A1(\core_pipeline.csr_to_fetch_mret_vector[5] ),
    .A2(net267),
    .B1(net247),
    .B2(\core_pipeline.pipeline_csr.instret[37] ),
    .X(_04875_));
 sky130_fd_sc_hd__a2111o_2 _08715_ (.A1(\core_pipeline.pipeline_csr.mtimecmp[37] ),
    .A2(net269),
    .B1(_04873_),
    .C1(_04874_),
    .D1(_04875_),
    .X(_04876_));
 sky130_fd_sc_hd__mux2_1 _08716_ (.A0(\core_pipeline.decode_to_execute_csr_data[5] ),
    .A1(_04876_),
    .S(net157),
    .X(_00426_));
 sky130_fd_sc_hd__a22o_1 _08717_ (.A1(\core_pipeline.pipeline_csr.instret[4] ),
    .A2(net249),
    .B1(net265),
    .B2(\core_pipeline.pipeline_csr.mscratch[4] ),
    .X(_04877_));
 sky130_fd_sc_hd__a221o_1 _08718_ (.A1(\core_pipeline.pipeline_csr.cycle[4] ),
    .A2(net251),
    .B1(net267),
    .B2(\core_pipeline.csr_to_fetch_mret_vector[4] ),
    .C1(_04877_),
    .X(_04878_));
 sky130_fd_sc_hd__a22o_1 _08719_ (.A1(\core_pipeline.pipeline_csr.instret[36] ),
    .A2(net247),
    .B1(net246),
    .B2(\core_pipeline.pipeline_csr.cycle[36] ),
    .X(_04879_));
 sky130_fd_sc_hd__a22o_1 _08720_ (.A1(\core_pipeline.csr_to_fetch_trap_vector[4] ),
    .A2(net271),
    .B1(net269),
    .B2(\core_pipeline.pipeline_csr.mtimecmp[36] ),
    .X(_04880_));
 sky130_fd_sc_hd__a211o_1 _08721_ (.A1(\core_pipeline.pipeline_csr.mtimecmp[4] ),
    .A2(net273),
    .B1(_04879_),
    .C1(_04880_),
    .X(_04881_));
 sky130_fd_sc_hd__or3_4 _08722_ (.A(net136),
    .B(_04878_),
    .C(_04881_),
    .X(_04882_));
 sky130_fd_sc_hd__o21a_1 _08723_ (.A1(\core_pipeline.decode_to_execute_csr_data[4] ),
    .A2(net152),
    .B1(_04882_),
    .X(_00427_));
 sky130_fd_sc_hd__and3_1 _08724_ (.A(\core_pipeline.pipeline_csr.ie ),
    .B(_04683_),
    .C(_04693_),
    .X(_04883_));
 sky130_fd_sc_hd__a22o_1 _08725_ (.A1(\core_pipeline.pipeline_csr.mcause[3] ),
    .A2(_04710_),
    .B1(net246),
    .B2(\core_pipeline.pipeline_csr.cycle[35] ),
    .X(_04884_));
 sky130_fd_sc_hd__a221o_1 _08726_ (.A1(\core_pipeline.pipeline_csr.mscratch[3] ),
    .A2(net265),
    .B1(_04722_),
    .B2(\core_pipeline.csr_to_fetch_trap_vector[3] ),
    .C1(_04884_),
    .X(_04885_));
 sky130_fd_sc_hd__a221o_1 _08727_ (.A1(\core_pipeline.pipeline_csr.mtimecmp[35] ),
    .A2(_04724_),
    .B1(_04834_),
    .B2(\core_pipeline.pipeline_csr.msie ),
    .C1(_04883_),
    .X(_04886_));
 sky130_fd_sc_hd__a22o_1 _08728_ (.A1(\core_pipeline.pipeline_csr.instret[3] ),
    .A2(net249),
    .B1(net247),
    .B2(\core_pipeline.pipeline_csr.instret[35] ),
    .X(_04887_));
 sky130_fd_sc_hd__a22o_1 _08729_ (.A1(\core_pipeline.csr_to_fetch_mret_vector[3] ),
    .A2(net267),
    .B1(_04725_),
    .B2(\core_pipeline.pipeline_csr.mtimecmp[3] ),
    .X(_04888_));
 sky130_fd_sc_hd__a211o_1 _08730_ (.A1(\core_pipeline.pipeline_csr.msip ),
    .A2(_04835_),
    .B1(_04888_),
    .C1(net134),
    .X(_04889_));
 sky130_fd_sc_hd__a2111o_1 _08731_ (.A1(\core_pipeline.pipeline_csr.cycle[3] ),
    .A2(net251),
    .B1(_04886_),
    .C1(_04887_),
    .D1(_04889_),
    .X(_04890_));
 sky130_fd_sc_hd__o22a_1 _08732_ (.A1(\core_pipeline.decode_to_execute_csr_data[3] ),
    .A2(net157),
    .B1(_04885_),
    .B2(_04890_),
    .X(_00428_));
 sky130_fd_sc_hd__a22o_1 _08733_ (.A1(\core_pipeline.pipeline_csr.mtimecmp[2] ),
    .A2(net273),
    .B1(net269),
    .B2(\core_pipeline.pipeline_csr.mtimecmp[34] ),
    .X(_04891_));
 sky130_fd_sc_hd__a22o_1 _08734_ (.A1(\core_pipeline.pipeline_csr.instret[2] ),
    .A2(net249),
    .B1(net247),
    .B2(\core_pipeline.pipeline_csr.instret[34] ),
    .X(_04892_));
 sky130_fd_sc_hd__a221o_1 _08735_ (.A1(\core_pipeline.pipeline_csr.cycle[2] ),
    .A2(net251),
    .B1(net267),
    .B2(\core_pipeline.csr_to_fetch_mret_vector[2] ),
    .C1(_04892_),
    .X(_04893_));
 sky130_fd_sc_hd__a211o_1 _08736_ (.A1(\core_pipeline.csr_to_fetch_trap_vector[2] ),
    .A2(net271),
    .B1(_04891_),
    .C1(_04893_),
    .X(_04894_));
 sky130_fd_sc_hd__a22o_1 _08737_ (.A1(\core_pipeline.pipeline_csr.mcause[2] ),
    .A2(_04710_),
    .B1(net246),
    .B2(\core_pipeline.pipeline_csr.cycle[34] ),
    .X(_04895_));
 sky130_fd_sc_hd__a211o_1 _08738_ (.A1(\core_pipeline.pipeline_csr.mscratch[2] ),
    .A2(net265),
    .B1(_04895_),
    .C1(net134),
    .X(_04896_));
 sky130_fd_sc_hd__o22a_1 _08739_ (.A1(\core_pipeline.decode_to_execute_csr_data[2] ),
    .A2(net159),
    .B1(_04894_),
    .B2(_04896_),
    .X(_00429_));
 sky130_fd_sc_hd__a22o_1 _08740_ (.A1(\core_pipeline.pipeline_csr.mscratch[1] ),
    .A2(net265),
    .B1(_04724_),
    .B2(\core_pipeline.pipeline_csr.mtimecmp[33] ),
    .X(_04897_));
 sky130_fd_sc_hd__a221o_1 _08741_ (.A1(\core_pipeline.pipeline_csr.mcause[1] ),
    .A2(_04710_),
    .B1(net247),
    .B2(\core_pipeline.pipeline_csr.instret[33] ),
    .C1(_04897_),
    .X(_04898_));
 sky130_fd_sc_hd__a22o_1 _08742_ (.A1(\core_pipeline.pipeline_csr.cycle[1] ),
    .A2(net251),
    .B1(net249),
    .B2(\core_pipeline.pipeline_csr.instret[1] ),
    .X(_04899_));
 sky130_fd_sc_hd__a22o_1 _08743_ (.A1(\core_pipeline.csr_to_fetch_mret_vector[1] ),
    .A2(net267),
    .B1(_04725_),
    .B2(\core_pipeline.pipeline_csr.mtimecmp[1] ),
    .X(_04900_));
 sky130_fd_sc_hd__a2111o_4 _08744_ (.A1(\core_pipeline.pipeline_csr.cycle[33] ),
    .A2(net246),
    .B1(_04898_),
    .C1(_04899_),
    .D1(_04900_),
    .X(_04901_));
 sky130_fd_sc_hd__mux2_1 _08745_ (.A0(\core_pipeline.decode_to_execute_csr_data[1] ),
    .A1(_04901_),
    .S(net152),
    .X(_00430_));
 sky130_fd_sc_hd__a22o_1 _08746_ (.A1(\core_pipeline.pipeline_csr.cycle[0] ),
    .A2(net251),
    .B1(_04710_),
    .B2(\core_pipeline.pipeline_csr.mcause[0] ),
    .X(_04902_));
 sky130_fd_sc_hd__a221o_2 _08747_ (.A1(\core_pipeline.pipeline_csr.instret[32] ),
    .A2(net247),
    .B1(net246),
    .B2(\core_pipeline.pipeline_csr.cycle[32] ),
    .C1(_04902_),
    .X(_04903_));
 sky130_fd_sc_hd__a22o_1 _08748_ (.A1(\core_pipeline.pipeline_csr.mtimecmp[0] ),
    .A2(net273),
    .B1(net269),
    .B2(\core_pipeline.pipeline_csr.mtimecmp[32] ),
    .X(_04904_));
 sky130_fd_sc_hd__a21o_1 _08749_ (.A1(\core_pipeline.csr_to_fetch_mret_vector[0] ),
    .A2(net267),
    .B1(_04904_),
    .X(_04905_));
 sky130_fd_sc_hd__a221o_1 _08750_ (.A1(\core_pipeline.pipeline_csr.instret[0] ),
    .A2(net249),
    .B1(net265),
    .B2(\core_pipeline.pipeline_csr.mscratch[0] ),
    .C1(_04905_),
    .X(_04906_));
 sky130_fd_sc_hd__or3_4 _08751_ (.A(net132),
    .B(_04903_),
    .C(_04906_),
    .X(_04907_));
 sky130_fd_sc_hd__o21a_1 _08752_ (.A1(\core_pipeline.decode_to_execute_csr_data[0] ),
    .A2(net152),
    .B1(_04907_),
    .X(_00431_));
 sky130_fd_sc_hd__or4_1 _08753_ (.A(\core_pipeline.fetch_to_decode_instruction[6] ),
    .B(\core_pipeline.fetch_to_decode_instruction[5] ),
    .C(\core_pipeline.fetch_to_decode_instruction[4] ),
    .D(_03634_),
    .X(_04908_));
 sky130_fd_sc_hd__nand2_1 _08754_ (.A(_03313_),
    .B(_03445_),
    .Y(_04909_));
 sky130_fd_sc_hd__a22o_1 _08755_ (.A1(_03313_),
    .A2(_03321_),
    .B1(_04908_),
    .B2(_04909_),
    .X(_04910_));
 sky130_fd_sc_hd__nor2_2 _08756_ (.A(\core_pipeline.fetch_to_decode_instruction[14] ),
    .B(_03448_),
    .Y(_04911_));
 sky130_fd_sc_hd__o21ai_1 _08757_ (.A1(_03438_),
    .A2(_04911_),
    .B1(_04910_),
    .Y(_04912_));
 sky130_fd_sc_hd__a21o_1 _08758_ (.A1(\core_pipeline.fetch_to_decode_instruction[13] ),
    .A2(_04626_),
    .B1(_04664_),
    .X(_04913_));
 sky130_fd_sc_hd__a21o_1 _08759_ (.A1(\core_pipeline.fetch_to_decode_instruction[13] ),
    .A2(\core_pipeline.fetch_to_decode_instruction[12] ),
    .B1(\core_pipeline.fetch_to_decode_instruction[14] ),
    .X(_04914_));
 sky130_fd_sc_hd__or4_1 _08760_ (.A(\core_pipeline.decode_to_csr_read_address[5] ),
    .B(\core_pipeline.decode_to_csr_read_address[7] ),
    .C(\core_pipeline.decode_to_csr_read_address[6] ),
    .D(\core_pipeline.decode_to_csr_read_address[11] ),
    .X(_04915_));
 sky130_fd_sc_hd__or3_4 _08761_ (.A(\core_pipeline.decode_to_csr_read_address[9] ),
    .B(\core_pipeline.decode_to_csr_read_address[8] ),
    .C(_04915_),
    .X(_04916_));
 sky130_fd_sc_hd__o221a_1 _08762_ (.A1(\core_pipeline.fetch_to_decode_instruction[14] ),
    .A2(_03448_),
    .B1(_04633_),
    .B2(\core_pipeline.fetch_to_decode_instruction[13] ),
    .C1(\core_pipeline.decode_to_csr_read_address[10] ),
    .X(_04917_));
 sky130_fd_sc_hd__o21a_1 _08763_ (.A1(_04916_),
    .A2(_04917_),
    .B1(_03461_),
    .X(_04918_));
 sky130_fd_sc_hd__a21o_1 _08764_ (.A1(_03313_),
    .A2(\core_pipeline.decode_to_csr_read_address[10] ),
    .B1(_04916_),
    .X(_04919_));
 sky130_fd_sc_hd__and4_1 _08765_ (.A(_03321_),
    .B(\core_pipeline.fetch_to_decode_instruction[12] ),
    .C(\core_pipeline.fetch_to_decode_instruction[4] ),
    .D(_04624_),
    .X(_04920_));
 sky130_fd_sc_hd__a221o_1 _08766_ (.A1(_04913_),
    .A2(_04914_),
    .B1(_04919_),
    .B2(_04920_),
    .C1(_04918_),
    .X(_04921_));
 sky130_fd_sc_hd__nor2_1 _08767_ (.A(net513),
    .B(_04696_),
    .Y(_04922_));
 sky130_fd_sc_hd__o31a_1 _08768_ (.A1(net513),
    .A2(\core_pipeline.decode_to_csr_read_address[9] ),
    .A3(_04696_),
    .B1(_04716_),
    .X(_04923_));
 sky130_fd_sc_hd__and2_1 _08769_ (.A(\core_pipeline.decode_to_csr_read_address[9] ),
    .B(_04696_),
    .X(_04924_));
 sky130_fd_sc_hd__or4b_2 _08770_ (.A(\core_pipeline.fetch_to_decode_instruction[7] ),
    .B(\core_pipeline.fetch_to_decode_instruction[9] ),
    .C(_03485_),
    .D_N(_04631_),
    .X(_04925_));
 sky130_fd_sc_hd__o2111a_1 _08771_ (.A1(_04716_),
    .A2(_04924_),
    .B1(_04911_),
    .C1(\core_pipeline.decode_to_csr_read_address[8] ),
    .D1(_03339_),
    .X(_04926_));
 sky130_fd_sc_hd__or4b_2 _08772_ (.A(_04915_),
    .B(_04923_),
    .C(_04925_),
    .D_N(_04926_),
    .X(_04927_));
 sky130_fd_sc_hd__nor3b_1 _08773_ (.A(_03452_),
    .B(_03637_),
    .C_N(_04908_),
    .Y(_04928_));
 sky130_fd_sc_hd__a31o_1 _08774_ (.A1(_03447_),
    .A2(_03451_),
    .A3(_04927_),
    .B1(_04928_),
    .X(_04929_));
 sky130_fd_sc_hd__o31a_2 _08775_ (.A1(_04912_),
    .A2(_04921_),
    .A3(_04929_),
    .B1(net143),
    .X(_04930_));
 sky130_fd_sc_hd__a21o_1 _08776_ (.A1(\core_pipeline.decode_to_execute_exception ),
    .A2(net133),
    .B1(_04930_),
    .X(_00432_));
 sky130_fd_sc_hd__nand2_1 _08777_ (.A(_03632_),
    .B(_04911_),
    .Y(_04931_));
 sky130_fd_sc_hd__or4_1 _08778_ (.A(net513),
    .B(\core_pipeline.decode_to_csr_read_address[10] ),
    .C(_04682_),
    .D(_04916_),
    .X(_04932_));
 sky130_fd_sc_hd__or3_1 _08779_ (.A(_04925_),
    .B(_04931_),
    .C(_04932_),
    .X(_04933_));
 sky130_fd_sc_hd__a2bb2o_1 _08780_ (.A1_N(net565),
    .A2_N(_04933_),
    .B1(net133),
    .B2(\core_pipeline.decode_to_execute_ecause[3] ),
    .X(_00433_));
 sky130_fd_sc_hd__a21o_1 _08781_ (.A1(\core_pipeline.decode_to_execute_ecause[1] ),
    .A2(net133),
    .B1(_04930_),
    .X(_00434_));
 sky130_fd_sc_hd__a21bo_1 _08782_ (.A1(\core_pipeline.decode_to_execute_ecause[0] ),
    .A2(net133),
    .B1_N(_04933_),
    .X(_00435_));
 sky130_fd_sc_hd__or2_4 _08783_ (.A(\core_pipeline.memory_to_writeback_rd_address[0] ),
    .B(_03914_),
    .X(_04934_));
 sky130_fd_sc_hd__or4_4 _08784_ (.A(\core_pipeline.memory_to_writeback_rd_address[2] ),
    .B(\core_pipeline.memory_to_writeback_rd_address[4] ),
    .C(_04468_),
    .D(_04934_),
    .X(_04935_));
 sky130_fd_sc_hd__mux2_1 _08785_ (.A0(net348),
    .A1(\core_pipeline.pipeline_registers.registers[10][0] ),
    .S(net219),
    .X(_00436_));
 sky130_fd_sc_hd__mux2_1 _08786_ (.A0(net347),
    .A1(\core_pipeline.pipeline_registers.registers[10][1] ),
    .S(net220),
    .X(_00437_));
 sky130_fd_sc_hd__mux2_1 _08787_ (.A0(net344),
    .A1(\core_pipeline.pipeline_registers.registers[10][2] ),
    .S(net220),
    .X(_00438_));
 sky130_fd_sc_hd__mux2_1 _08788_ (.A0(net343),
    .A1(\core_pipeline.pipeline_registers.registers[10][3] ),
    .S(net219),
    .X(_00439_));
 sky130_fd_sc_hd__mux2_1 _08789_ (.A0(net340),
    .A1(\core_pipeline.pipeline_registers.registers[10][4] ),
    .S(net219),
    .X(_00440_));
 sky130_fd_sc_hd__mux2_1 _08790_ (.A0(net337),
    .A1(\core_pipeline.pipeline_registers.registers[10][5] ),
    .S(net220),
    .X(_00441_));
 sky130_fd_sc_hd__mux2_1 _08791_ (.A0(net335),
    .A1(\core_pipeline.pipeline_registers.registers[10][6] ),
    .S(net219),
    .X(_00442_));
 sky130_fd_sc_hd__mux2_1 _08792_ (.A0(net334),
    .A1(\core_pipeline.pipeline_registers.registers[10][7] ),
    .S(net219),
    .X(_00443_));
 sky130_fd_sc_hd__mux2_1 _08793_ (.A0(net332),
    .A1(\core_pipeline.pipeline_registers.registers[10][8] ),
    .S(net219),
    .X(_00444_));
 sky130_fd_sc_hd__mux2_1 _08794_ (.A0(net329),
    .A1(\core_pipeline.pipeline_registers.registers[10][9] ),
    .S(net219),
    .X(_00445_));
 sky130_fd_sc_hd__mux2_1 _08795_ (.A0(net327),
    .A1(\core_pipeline.pipeline_registers.registers[10][10] ),
    .S(net219),
    .X(_00446_));
 sky130_fd_sc_hd__mux2_1 _08796_ (.A0(net325),
    .A1(\core_pipeline.pipeline_registers.registers[10][11] ),
    .S(net219),
    .X(_00447_));
 sky130_fd_sc_hd__mux2_1 _08797_ (.A0(net323),
    .A1(\core_pipeline.pipeline_registers.registers[10][12] ),
    .S(net219),
    .X(_00448_));
 sky130_fd_sc_hd__mux2_1 _08798_ (.A0(net321),
    .A1(\core_pipeline.pipeline_registers.registers[10][13] ),
    .S(net219),
    .X(_00449_));
 sky130_fd_sc_hd__mux2_1 _08799_ (.A0(net319),
    .A1(\core_pipeline.pipeline_registers.registers[10][14] ),
    .S(net219),
    .X(_00450_));
 sky130_fd_sc_hd__mux2_1 _08800_ (.A0(net317),
    .A1(\core_pipeline.pipeline_registers.registers[10][15] ),
    .S(net219),
    .X(_00451_));
 sky130_fd_sc_hd__mux2_1 _08801_ (.A0(net315),
    .A1(\core_pipeline.pipeline_registers.registers[10][16] ),
    .S(net219),
    .X(_00452_));
 sky130_fd_sc_hd__mux2_1 _08802_ (.A0(net312),
    .A1(\core_pipeline.pipeline_registers.registers[10][17] ),
    .S(net220),
    .X(_00453_));
 sky130_fd_sc_hd__mux2_1 _08803_ (.A0(net311),
    .A1(\core_pipeline.pipeline_registers.registers[10][18] ),
    .S(net220),
    .X(_00454_));
 sky130_fd_sc_hd__mux2_1 _08804_ (.A0(net308),
    .A1(\core_pipeline.pipeline_registers.registers[10][19] ),
    .S(net220),
    .X(_00455_));
 sky130_fd_sc_hd__mux2_1 _08805_ (.A0(net306),
    .A1(\core_pipeline.pipeline_registers.registers[10][20] ),
    .S(net220),
    .X(_00456_));
 sky130_fd_sc_hd__mux2_1 _08806_ (.A0(net303),
    .A1(\core_pipeline.pipeline_registers.registers[10][21] ),
    .S(net220),
    .X(_00457_));
 sky130_fd_sc_hd__mux2_1 _08807_ (.A0(net301),
    .A1(\core_pipeline.pipeline_registers.registers[10][22] ),
    .S(net220),
    .X(_00458_));
 sky130_fd_sc_hd__mux2_1 _08808_ (.A0(net300),
    .A1(\core_pipeline.pipeline_registers.registers[10][23] ),
    .S(net220),
    .X(_00459_));
 sky130_fd_sc_hd__mux2_1 _08809_ (.A0(net297),
    .A1(\core_pipeline.pipeline_registers.registers[10][24] ),
    .S(net219),
    .X(_00460_));
 sky130_fd_sc_hd__mux2_1 _08810_ (.A0(net295),
    .A1(\core_pipeline.pipeline_registers.registers[10][25] ),
    .S(net219),
    .X(_00461_));
 sky130_fd_sc_hd__mux2_1 _08811_ (.A0(net293),
    .A1(\core_pipeline.pipeline_registers.registers[10][26] ),
    .S(net219),
    .X(_00462_));
 sky130_fd_sc_hd__mux2_1 _08812_ (.A0(net292),
    .A1(\core_pipeline.pipeline_registers.registers[10][27] ),
    .S(net220),
    .X(_00463_));
 sky130_fd_sc_hd__mux2_1 _08813_ (.A0(net289),
    .A1(\core_pipeline.pipeline_registers.registers[10][28] ),
    .S(net220),
    .X(_00464_));
 sky130_fd_sc_hd__mux2_1 _08814_ (.A0(net286),
    .A1(\core_pipeline.pipeline_registers.registers[10][29] ),
    .S(net220),
    .X(_00465_));
 sky130_fd_sc_hd__mux2_1 _08815_ (.A0(net284),
    .A1(\core_pipeline.pipeline_registers.registers[10][30] ),
    .S(net220),
    .X(_00466_));
 sky130_fd_sc_hd__mux2_1 _08816_ (.A0(net282),
    .A1(\core_pipeline.pipeline_registers.registers[10][31] ),
    .S(net220),
    .X(_00467_));
 sky130_fd_sc_hd__nand2_2 _08817_ (.A(\core_pipeline.memory_to_writeback_rd_address[2] ),
    .B(_03480_),
    .Y(_04936_));
 sky130_fd_sc_hd__o31a_4 _08818_ (.A1(\core_pipeline.memory_to_writeback_rd_address[2] ),
    .A2(\core_pipeline.memory_to_writeback_rd_address[3] ),
    .A3(\core_pipeline.memory_to_writeback_rd_address[4] ),
    .B1(_03480_),
    .X(_04937_));
 sky130_fd_sc_hd__nor2_8 _08819_ (.A(_04934_),
    .B(_04937_),
    .Y(_04938_));
 sky130_fd_sc_hd__mux2_1 _08820_ (.A0(\core_pipeline.pipeline_registers.registers[2][0] ),
    .A1(net348),
    .S(net217),
    .X(_00468_));
 sky130_fd_sc_hd__mux2_1 _08821_ (.A0(\core_pipeline.pipeline_registers.registers[2][1] ),
    .A1(net347),
    .S(net218),
    .X(_00469_));
 sky130_fd_sc_hd__mux2_1 _08822_ (.A0(\core_pipeline.pipeline_registers.registers[2][2] ),
    .A1(net345),
    .S(net218),
    .X(_00470_));
 sky130_fd_sc_hd__mux2_1 _08823_ (.A0(\core_pipeline.pipeline_registers.registers[2][3] ),
    .A1(net343),
    .S(net217),
    .X(_00471_));
 sky130_fd_sc_hd__mux2_1 _08824_ (.A0(\core_pipeline.pipeline_registers.registers[2][4] ),
    .A1(net340),
    .S(net217),
    .X(_00472_));
 sky130_fd_sc_hd__mux2_1 _08825_ (.A0(\core_pipeline.pipeline_registers.registers[2][5] ),
    .A1(net338),
    .S(net218),
    .X(_00473_));
 sky130_fd_sc_hd__mux2_1 _08826_ (.A0(\core_pipeline.pipeline_registers.registers[2][6] ),
    .A1(net335),
    .S(net217),
    .X(_00474_));
 sky130_fd_sc_hd__mux2_1 _08827_ (.A0(\core_pipeline.pipeline_registers.registers[2][7] ),
    .A1(net334),
    .S(net217),
    .X(_00475_));
 sky130_fd_sc_hd__mux2_1 _08828_ (.A0(\core_pipeline.pipeline_registers.registers[2][8] ),
    .A1(net332),
    .S(net217),
    .X(_00476_));
 sky130_fd_sc_hd__mux2_1 _08829_ (.A0(\core_pipeline.pipeline_registers.registers[2][9] ),
    .A1(net329),
    .S(net217),
    .X(_00477_));
 sky130_fd_sc_hd__mux2_1 _08830_ (.A0(\core_pipeline.pipeline_registers.registers[2][10] ),
    .A1(net328),
    .S(net217),
    .X(_00478_));
 sky130_fd_sc_hd__mux2_1 _08831_ (.A0(\core_pipeline.pipeline_registers.registers[2][11] ),
    .A1(net325),
    .S(net217),
    .X(_00479_));
 sky130_fd_sc_hd__mux2_1 _08832_ (.A0(\core_pipeline.pipeline_registers.registers[2][12] ),
    .A1(net324),
    .S(net217),
    .X(_00480_));
 sky130_fd_sc_hd__mux2_1 _08833_ (.A0(\core_pipeline.pipeline_registers.registers[2][13] ),
    .A1(net322),
    .S(net217),
    .X(_00481_));
 sky130_fd_sc_hd__mux2_1 _08834_ (.A0(\core_pipeline.pipeline_registers.registers[2][14] ),
    .A1(net320),
    .S(net217),
    .X(_00482_));
 sky130_fd_sc_hd__mux2_1 _08835_ (.A0(\core_pipeline.pipeline_registers.registers[2][15] ),
    .A1(net317),
    .S(net217),
    .X(_00483_));
 sky130_fd_sc_hd__mux2_1 _08836_ (.A0(\core_pipeline.pipeline_registers.registers[2][16] ),
    .A1(net315),
    .S(net217),
    .X(_00484_));
 sky130_fd_sc_hd__mux2_1 _08837_ (.A0(\core_pipeline.pipeline_registers.registers[2][17] ),
    .A1(net312),
    .S(net218),
    .X(_00485_));
 sky130_fd_sc_hd__mux2_1 _08838_ (.A0(\core_pipeline.pipeline_registers.registers[2][18] ),
    .A1(net310),
    .S(net218),
    .X(_00486_));
 sky130_fd_sc_hd__mux2_1 _08839_ (.A0(\core_pipeline.pipeline_registers.registers[2][19] ),
    .A1(net308),
    .S(net218),
    .X(_00487_));
 sky130_fd_sc_hd__mux2_1 _08840_ (.A0(\core_pipeline.pipeline_registers.registers[2][20] ),
    .A1(net305),
    .S(net218),
    .X(_00488_));
 sky130_fd_sc_hd__mux2_1 _08841_ (.A0(\core_pipeline.pipeline_registers.registers[2][21] ),
    .A1(net303),
    .S(net218),
    .X(_00489_));
 sky130_fd_sc_hd__mux2_1 _08842_ (.A0(\core_pipeline.pipeline_registers.registers[2][22] ),
    .A1(net301),
    .S(net218),
    .X(_00490_));
 sky130_fd_sc_hd__mux2_1 _08843_ (.A0(\core_pipeline.pipeline_registers.registers[2][23] ),
    .A1(net300),
    .S(net218),
    .X(_00491_));
 sky130_fd_sc_hd__mux2_1 _08844_ (.A0(\core_pipeline.pipeline_registers.registers[2][24] ),
    .A1(net298),
    .S(net217),
    .X(_00492_));
 sky130_fd_sc_hd__mux2_1 _08845_ (.A0(\core_pipeline.pipeline_registers.registers[2][25] ),
    .A1(net295),
    .S(net217),
    .X(_00493_));
 sky130_fd_sc_hd__mux2_1 _08846_ (.A0(\core_pipeline.pipeline_registers.registers[2][26] ),
    .A1(net293),
    .S(net217),
    .X(_00494_));
 sky130_fd_sc_hd__mux2_1 _08847_ (.A0(\core_pipeline.pipeline_registers.registers[2][27] ),
    .A1(net292),
    .S(net218),
    .X(_00495_));
 sky130_fd_sc_hd__mux2_1 _08848_ (.A0(\core_pipeline.pipeline_registers.registers[2][28] ),
    .A1(net289),
    .S(net218),
    .X(_00496_));
 sky130_fd_sc_hd__mux2_1 _08849_ (.A0(\core_pipeline.pipeline_registers.registers[2][29] ),
    .A1(net288),
    .S(net218),
    .X(_00497_));
 sky130_fd_sc_hd__mux2_1 _08850_ (.A0(\core_pipeline.pipeline_registers.registers[2][30] ),
    .A1(net284),
    .S(net218),
    .X(_00498_));
 sky130_fd_sc_hd__mux2_1 _08851_ (.A0(\core_pipeline.pipeline_registers.registers[2][31] ),
    .A1(net283),
    .S(net218),
    .X(_00499_));
 sky130_fd_sc_hd__nand2_8 _08852_ (.A(_03913_),
    .B(_03914_),
    .Y(_04939_));
 sky130_fd_sc_hd__nor2_8 _08853_ (.A(_04469_),
    .B(_04939_),
    .Y(_04940_));
 sky130_fd_sc_hd__mux2_1 _08854_ (.A0(\core_pipeline.pipeline_registers.registers[28][0] ),
    .A1(net349),
    .S(net215),
    .X(_00500_));
 sky130_fd_sc_hd__mux2_1 _08855_ (.A0(\core_pipeline.pipeline_registers.registers[28][1] ),
    .A1(net346),
    .S(net216),
    .X(_00501_));
 sky130_fd_sc_hd__mux2_1 _08856_ (.A0(\core_pipeline.pipeline_registers.registers[28][2] ),
    .A1(net344),
    .S(net216),
    .X(_00502_));
 sky130_fd_sc_hd__mux2_1 _08857_ (.A0(\core_pipeline.pipeline_registers.registers[28][3] ),
    .A1(net342),
    .S(net215),
    .X(_00503_));
 sky130_fd_sc_hd__mux2_1 _08858_ (.A0(\core_pipeline.pipeline_registers.registers[28][4] ),
    .A1(net341),
    .S(net215),
    .X(_00504_));
 sky130_fd_sc_hd__mux2_1 _08859_ (.A0(\core_pipeline.pipeline_registers.registers[28][5] ),
    .A1(net338),
    .S(net216),
    .X(_00505_));
 sky130_fd_sc_hd__mux2_1 _08860_ (.A0(\core_pipeline.pipeline_registers.registers[28][6] ),
    .A1(net335),
    .S(net216),
    .X(_00506_));
 sky130_fd_sc_hd__mux2_1 _08861_ (.A0(\core_pipeline.pipeline_registers.registers[28][7] ),
    .A1(net333),
    .S(net215),
    .X(_00507_));
 sky130_fd_sc_hd__mux2_1 _08862_ (.A0(\core_pipeline.pipeline_registers.registers[28][8] ),
    .A1(net331),
    .S(net215),
    .X(_00508_));
 sky130_fd_sc_hd__mux2_1 _08863_ (.A0(\core_pipeline.pipeline_registers.registers[28][9] ),
    .A1(net330),
    .S(net215),
    .X(_00509_));
 sky130_fd_sc_hd__mux2_1 _08864_ (.A0(\core_pipeline.pipeline_registers.registers[28][10] ),
    .A1(net328),
    .S(net215),
    .X(_00510_));
 sky130_fd_sc_hd__mux2_1 _08865_ (.A0(\core_pipeline.pipeline_registers.registers[28][11] ),
    .A1(net326),
    .S(net215),
    .X(_00511_));
 sky130_fd_sc_hd__mux2_1 _08866_ (.A0(\core_pipeline.pipeline_registers.registers[28][12] ),
    .A1(net324),
    .S(net215),
    .X(_00512_));
 sky130_fd_sc_hd__mux2_1 _08867_ (.A0(\core_pipeline.pipeline_registers.registers[28][13] ),
    .A1(net322),
    .S(net215),
    .X(_00513_));
 sky130_fd_sc_hd__mux2_1 _08868_ (.A0(\core_pipeline.pipeline_registers.registers[28][14] ),
    .A1(net319),
    .S(net215),
    .X(_00514_));
 sky130_fd_sc_hd__mux2_1 _08869_ (.A0(\core_pipeline.pipeline_registers.registers[28][15] ),
    .A1(net318),
    .S(net215),
    .X(_00515_));
 sky130_fd_sc_hd__mux2_1 _08870_ (.A0(\core_pipeline.pipeline_registers.registers[28][16] ),
    .A1(net315),
    .S(net215),
    .X(_00516_));
 sky130_fd_sc_hd__mux2_1 _08871_ (.A0(\core_pipeline.pipeline_registers.registers[28][17] ),
    .A1(net312),
    .S(net216),
    .X(_00517_));
 sky130_fd_sc_hd__mux2_1 _08872_ (.A0(\core_pipeline.pipeline_registers.registers[28][18] ),
    .A1(net310),
    .S(net216),
    .X(_00518_));
 sky130_fd_sc_hd__mux2_1 _08873_ (.A0(\core_pipeline.pipeline_registers.registers[28][19] ),
    .A1(net309),
    .S(net216),
    .X(_00519_));
 sky130_fd_sc_hd__mux2_1 _08874_ (.A0(\core_pipeline.pipeline_registers.registers[28][20] ),
    .A1(net305),
    .S(net216),
    .X(_00520_));
 sky130_fd_sc_hd__mux2_1 _08875_ (.A0(\core_pipeline.pipeline_registers.registers[28][21] ),
    .A1(net303),
    .S(net216),
    .X(_00521_));
 sky130_fd_sc_hd__mux2_1 _08876_ (.A0(\core_pipeline.pipeline_registers.registers[28][22] ),
    .A1(net302),
    .S(net215),
    .X(_00522_));
 sky130_fd_sc_hd__mux2_1 _08877_ (.A0(\core_pipeline.pipeline_registers.registers[28][23] ),
    .A1(net300),
    .S(net216),
    .X(_00523_));
 sky130_fd_sc_hd__mux2_1 _08878_ (.A0(\core_pipeline.pipeline_registers.registers[28][24] ),
    .A1(net298),
    .S(net215),
    .X(_00524_));
 sky130_fd_sc_hd__mux2_1 _08879_ (.A0(\core_pipeline.pipeline_registers.registers[28][25] ),
    .A1(net296),
    .S(net215),
    .X(_00525_));
 sky130_fd_sc_hd__mux2_1 _08880_ (.A0(\core_pipeline.pipeline_registers.registers[28][26] ),
    .A1(net294),
    .S(net215),
    .X(_00526_));
 sky130_fd_sc_hd__mux2_1 _08881_ (.A0(\core_pipeline.pipeline_registers.registers[28][27] ),
    .A1(net291),
    .S(net216),
    .X(_00527_));
 sky130_fd_sc_hd__mux2_1 _08882_ (.A0(\core_pipeline.pipeline_registers.registers[28][28] ),
    .A1(net290),
    .S(net216),
    .X(_00528_));
 sky130_fd_sc_hd__mux2_1 _08883_ (.A0(\core_pipeline.pipeline_registers.registers[28][29] ),
    .A1(net286),
    .S(net216),
    .X(_00529_));
 sky130_fd_sc_hd__mux2_1 _08884_ (.A0(\core_pipeline.pipeline_registers.registers[28][30] ),
    .A1(net284),
    .S(net216),
    .X(_00530_));
 sky130_fd_sc_hd__mux2_1 _08885_ (.A0(\core_pipeline.pipeline_registers.registers[28][31] ),
    .A1(net282),
    .S(net216),
    .X(_00531_));
 sky130_fd_sc_hd__mux4_1 _08886_ (.A0(\core_pipeline.pipeline_registers.registers[8][0] ),
    .A1(\core_pipeline.pipeline_registers.registers[9][0] ),
    .A2(\core_pipeline.pipeline_registers.registers[10][0] ),
    .A3(\core_pipeline.pipeline_registers.registers[11][0] ),
    .S0(net544),
    .S1(net525),
    .X(_04941_));
 sky130_fd_sc_hd__or2_1 _08887_ (.A(net519),
    .B(_04941_),
    .X(_04942_));
 sky130_fd_sc_hd__mux4_1 _08888_ (.A0(\core_pipeline.pipeline_registers.registers[12][0] ),
    .A1(\core_pipeline.pipeline_registers.registers[13][0] ),
    .A2(\core_pipeline.pipeline_registers.registers[14][0] ),
    .A3(\core_pipeline.pipeline_registers.registers[15][0] ),
    .S0(net544),
    .S1(net525),
    .X(_04943_));
 sky130_fd_sc_hd__o211a_1 _08889_ (.A1(net462),
    .A2(_04943_),
    .B1(_04942_),
    .C1(net514),
    .X(_04944_));
 sky130_fd_sc_hd__mux4_1 _08890_ (.A0(\core_pipeline.pipeline_registers.registers[0][0] ),
    .A1(\core_pipeline.pipeline_registers.registers[1][0] ),
    .A2(\core_pipeline.pipeline_registers.registers[2][0] ),
    .A3(\core_pipeline.pipeline_registers.registers[3][0] ),
    .S0(net544),
    .S1(net525),
    .X(_04945_));
 sky130_fd_sc_hd__mux4_1 _08891_ (.A0(\core_pipeline.pipeline_registers.registers[4][0] ),
    .A1(\core_pipeline.pipeline_registers.registers[5][0] ),
    .A2(\core_pipeline.pipeline_registers.registers[6][0] ),
    .A3(\core_pipeline.pipeline_registers.registers[7][0] ),
    .S0(net545),
    .S1(net528),
    .X(_04946_));
 sky130_fd_sc_hd__a221o_1 _08892_ (.A1(net428),
    .A2(_04945_),
    .B1(_04946_),
    .B2(net367),
    .C1(_04944_),
    .X(_04947_));
 sky130_fd_sc_hd__mux2_1 _08893_ (.A0(\core_pipeline.pipeline_registers.registers[26][0] ),
    .A1(\core_pipeline.pipeline_registers.registers[27][0] ),
    .S(net548),
    .X(_04948_));
 sky130_fd_sc_hd__a221o_1 _08894_ (.A1(\core_pipeline.pipeline_registers.registers[24][0] ),
    .A2(net424),
    .B1(net363),
    .B2(\core_pipeline.pipeline_registers.registers[25][0] ),
    .C1(net519),
    .X(_04949_));
 sky130_fd_sc_hd__a21o_1 _08895_ (.A1(net529),
    .A2(_04948_),
    .B1(_04949_),
    .X(_04950_));
 sky130_fd_sc_hd__mux2_1 _08896_ (.A0(\core_pipeline.pipeline_registers.registers[30][0] ),
    .A1(\core_pipeline.pipeline_registers.registers[31][0] ),
    .S(net548),
    .X(_04951_));
 sky130_fd_sc_hd__a221o_1 _08897_ (.A1(\core_pipeline.pipeline_registers.registers[28][0] ),
    .A2(net424),
    .B1(net363),
    .B2(\core_pipeline.pipeline_registers.registers[29][0] ),
    .C1(net462),
    .X(_04952_));
 sky130_fd_sc_hd__a21o_1 _08898_ (.A1(net529),
    .A2(_04951_),
    .B1(_04952_),
    .X(_04953_));
 sky130_fd_sc_hd__mux4_1 _08899_ (.A0(\core_pipeline.pipeline_registers.registers[16][0] ),
    .A1(\core_pipeline.pipeline_registers.registers[17][0] ),
    .A2(\core_pipeline.pipeline_registers.registers[18][0] ),
    .A3(\core_pipeline.pipeline_registers.registers[19][0] ),
    .S0(net545),
    .S1(net528),
    .X(_04954_));
 sky130_fd_sc_hd__mux4_1 _08900_ (.A0(\core_pipeline.pipeline_registers.registers[20][0] ),
    .A1(\core_pipeline.pipeline_registers.registers[21][0] ),
    .A2(\core_pipeline.pipeline_registers.registers[22][0] ),
    .A3(\core_pipeline.pipeline_registers.registers[23][0] ),
    .S0(net545),
    .S1(net528),
    .X(_04955_));
 sky130_fd_sc_hd__a22o_1 _08901_ (.A1(net428),
    .A2(_04954_),
    .B1(_04955_),
    .B2(net367),
    .X(_04956_));
 sky130_fd_sc_hd__a31o_1 _08902_ (.A1(net514),
    .A2(_04950_),
    .A3(_04953_),
    .B1(net461),
    .X(_04957_));
 sky130_fd_sc_hd__o22a_2 _08903_ (.A1(net511),
    .A2(_04947_),
    .B1(_04956_),
    .B2(_04957_),
    .X(_04958_));
 sky130_fd_sc_hd__mux2_1 _08904_ (.A0(\core_pipeline.decode_to_execute_rs2_data[0] ),
    .A1(_04958_),
    .S(net140),
    .X(_00532_));
 sky130_fd_sc_hd__mux4_1 _08905_ (.A0(\core_pipeline.pipeline_registers.registers[8][1] ),
    .A1(\core_pipeline.pipeline_registers.registers[9][1] ),
    .A2(\core_pipeline.pipeline_registers.registers[10][1] ),
    .A3(\core_pipeline.pipeline_registers.registers[11][1] ),
    .S0(net563),
    .S1(net540),
    .X(_04959_));
 sky130_fd_sc_hd__or2_1 _08906_ (.A(net524),
    .B(_04959_),
    .X(_04960_));
 sky130_fd_sc_hd__mux4_1 _08907_ (.A0(\core_pipeline.pipeline_registers.registers[12][1] ),
    .A1(\core_pipeline.pipeline_registers.registers[13][1] ),
    .A2(\core_pipeline.pipeline_registers.registers[14][1] ),
    .A3(\core_pipeline.pipeline_registers.registers[15][1] ),
    .S0(net563),
    .S1(net540),
    .X(_04961_));
 sky130_fd_sc_hd__o211a_1 _08908_ (.A1(net465),
    .A2(_04961_),
    .B1(_04960_),
    .C1(net517),
    .X(_04962_));
 sky130_fd_sc_hd__mux4_1 _08909_ (.A0(\core_pipeline.pipeline_registers.registers[4][1] ),
    .A1(\core_pipeline.pipeline_registers.registers[5][1] ),
    .A2(\core_pipeline.pipeline_registers.registers[6][1] ),
    .A3(\core_pipeline.pipeline_registers.registers[7][1] ),
    .S0(net563),
    .S1(net540),
    .X(_04963_));
 sky130_fd_sc_hd__mux2_1 _08910_ (.A0(\core_pipeline.pipeline_registers.registers[2][1] ),
    .A1(\core_pipeline.pipeline_registers.registers[3][1] ),
    .S(net565),
    .X(_04964_));
 sky130_fd_sc_hd__a31o_1 _08911_ (.A1(net542),
    .A2(net430),
    .A3(_04964_),
    .B1(net512),
    .X(_04965_));
 sky130_fd_sc_hd__a221o_1 _08912_ (.A1(\core_pipeline.pipeline_registers.registers[0][1] ),
    .A2(net279),
    .B1(net276),
    .B2(\core_pipeline.pipeline_registers.registers[1][1] ),
    .C1(_04965_),
    .X(_04966_));
 sky130_fd_sc_hd__a211o_1 _08913_ (.A1(net369),
    .A2(_04963_),
    .B1(_04966_),
    .C1(_04962_),
    .X(_04967_));
 sky130_fd_sc_hd__mux2_1 _08914_ (.A0(\core_pipeline.pipeline_registers.registers[30][1] ),
    .A1(\core_pipeline.pipeline_registers.registers[31][1] ),
    .S(net563),
    .X(_04968_));
 sky130_fd_sc_hd__a221o_1 _08915_ (.A1(\core_pipeline.pipeline_registers.registers[28][1] ),
    .A2(net427),
    .B1(_04695_),
    .B2(\core_pipeline.pipeline_registers.registers[29][1] ),
    .C1(net465),
    .X(_04969_));
 sky130_fd_sc_hd__a21o_1 _08916_ (.A1(net540),
    .A2(_04968_),
    .B1(_04969_),
    .X(_04970_));
 sky130_fd_sc_hd__mux2_1 _08917_ (.A0(\core_pipeline.pipeline_registers.registers[26][1] ),
    .A1(\core_pipeline.pipeline_registers.registers[27][1] ),
    .S(net561),
    .X(_04971_));
 sky130_fd_sc_hd__a221o_1 _08918_ (.A1(\core_pipeline.pipeline_registers.registers[24][1] ),
    .A2(net427),
    .B1(_04695_),
    .B2(\core_pipeline.pipeline_registers.registers[25][1] ),
    .C1(net522),
    .X(_04972_));
 sky130_fd_sc_hd__a21o_1 _08919_ (.A1(net538),
    .A2(_04971_),
    .B1(_04972_),
    .X(_04973_));
 sky130_fd_sc_hd__and3_1 _08920_ (.A(net517),
    .B(_04970_),
    .C(_04973_),
    .X(_04974_));
 sky130_fd_sc_hd__mux4_1 _08921_ (.A0(\core_pipeline.pipeline_registers.registers[20][1] ),
    .A1(\core_pipeline.pipeline_registers.registers[21][1] ),
    .A2(\core_pipeline.pipeline_registers.registers[22][1] ),
    .A3(\core_pipeline.pipeline_registers.registers[23][1] ),
    .S0(net565),
    .S1(net542),
    .X(_04975_));
 sky130_fd_sc_hd__mux2_1 _08922_ (.A0(\core_pipeline.pipeline_registers.registers[18][1] ),
    .A1(\core_pipeline.pipeline_registers.registers[19][1] ),
    .S(net561),
    .X(_04976_));
 sky130_fd_sc_hd__a31o_1 _08923_ (.A1(net540),
    .A2(net430),
    .A3(_04976_),
    .B1(net460),
    .X(_04977_));
 sky130_fd_sc_hd__a221o_1 _08924_ (.A1(\core_pipeline.pipeline_registers.registers[16][1] ),
    .A2(net278),
    .B1(net276),
    .B2(\core_pipeline.pipeline_registers.registers[17][1] ),
    .C1(_04977_),
    .X(_04978_));
 sky130_fd_sc_hd__a211o_1 _08925_ (.A1(_04694_),
    .A2(_04975_),
    .B1(_04978_),
    .C1(_04974_),
    .X(_04979_));
 sky130_fd_sc_hd__and3_2 _08926_ (.A(net146),
    .B(_04967_),
    .C(_04979_),
    .X(_04980_));
 sky130_fd_sc_hd__a21o_1 _08927_ (.A1(\core_pipeline.decode_to_execute_rs2_data[1] ),
    .A2(net125),
    .B1(_04980_),
    .X(_00533_));
 sky130_fd_sc_hd__mux4_1 _08928_ (.A0(\core_pipeline.pipeline_registers.registers[8][2] ),
    .A1(\core_pipeline.pipeline_registers.registers[9][2] ),
    .A2(\core_pipeline.pipeline_registers.registers[10][2] ),
    .A3(\core_pipeline.pipeline_registers.registers[11][2] ),
    .S0(net559),
    .S1(net537),
    .X(_04981_));
 sky130_fd_sc_hd__or2_1 _08929_ (.A(net523),
    .B(_04981_),
    .X(_04982_));
 sky130_fd_sc_hd__mux4_1 _08930_ (.A0(\core_pipeline.pipeline_registers.registers[12][2] ),
    .A1(\core_pipeline.pipeline_registers.registers[13][2] ),
    .A2(\core_pipeline.pipeline_registers.registers[14][2] ),
    .A3(\core_pipeline.pipeline_registers.registers[15][2] ),
    .S0(net559),
    .S1(net537),
    .X(_04983_));
 sky130_fd_sc_hd__o211a_1 _08931_ (.A1(net465),
    .A2(_04983_),
    .B1(_04982_),
    .C1(net518),
    .X(_04984_));
 sky130_fd_sc_hd__mux4_1 _08932_ (.A0(\core_pipeline.pipeline_registers.registers[4][2] ),
    .A1(\core_pipeline.pipeline_registers.registers[5][2] ),
    .A2(\core_pipeline.pipeline_registers.registers[6][2] ),
    .A3(\core_pipeline.pipeline_registers.registers[7][2] ),
    .S0(net559),
    .S1(net537),
    .X(_04985_));
 sky130_fd_sc_hd__mux2_1 _08933_ (.A0(\core_pipeline.pipeline_registers.registers[2][2] ),
    .A1(\core_pipeline.pipeline_registers.registers[3][2] ),
    .S(net559),
    .X(_04986_));
 sky130_fd_sc_hd__a22o_1 _08934_ (.A1(\core_pipeline.pipeline_registers.registers[1][2] ),
    .A2(net276),
    .B1(net361),
    .B2(_04986_),
    .X(_04987_));
 sky130_fd_sc_hd__a211o_1 _08935_ (.A1(\core_pipeline.pipeline_registers.registers[0][2] ),
    .A2(net278),
    .B1(_04987_),
    .C1(net512),
    .X(_04988_));
 sky130_fd_sc_hd__a211o_1 _08936_ (.A1(net369),
    .A2(_04985_),
    .B1(_04988_),
    .C1(_04984_),
    .X(_04989_));
 sky130_fd_sc_hd__mux2_1 _08937_ (.A0(\core_pipeline.pipeline_registers.registers[30][2] ),
    .A1(\core_pipeline.pipeline_registers.registers[31][2] ),
    .S(net559),
    .X(_04990_));
 sky130_fd_sc_hd__a221o_1 _08938_ (.A1(\core_pipeline.pipeline_registers.registers[28][2] ),
    .A2(net427),
    .B1(net365),
    .B2(\core_pipeline.pipeline_registers.registers[29][2] ),
    .C1(net464),
    .X(_04991_));
 sky130_fd_sc_hd__a21o_1 _08939_ (.A1(net537),
    .A2(_04990_),
    .B1(_04991_),
    .X(_04992_));
 sky130_fd_sc_hd__mux2_1 _08940_ (.A0(\core_pipeline.pipeline_registers.registers[26][2] ),
    .A1(\core_pipeline.pipeline_registers.registers[27][2] ),
    .S(net559),
    .X(_04993_));
 sky130_fd_sc_hd__a221o_1 _08941_ (.A1(\core_pipeline.pipeline_registers.registers[24][2] ),
    .A2(net427),
    .B1(net366),
    .B2(\core_pipeline.pipeline_registers.registers[25][2] ),
    .C1(net523),
    .X(_04994_));
 sky130_fd_sc_hd__a21o_1 _08942_ (.A1(net534),
    .A2(_04993_),
    .B1(_04994_),
    .X(_04995_));
 sky130_fd_sc_hd__and3_1 _08943_ (.A(net516),
    .B(_04992_),
    .C(_04995_),
    .X(_04996_));
 sky130_fd_sc_hd__mux4_1 _08944_ (.A0(\core_pipeline.pipeline_registers.registers[20][2] ),
    .A1(\core_pipeline.pipeline_registers.registers[21][2] ),
    .A2(\core_pipeline.pipeline_registers.registers[22][2] ),
    .A3(\core_pipeline.pipeline_registers.registers[23][2] ),
    .S0(net556),
    .S1(net536),
    .X(_04997_));
 sky130_fd_sc_hd__mux2_1 _08945_ (.A0(\core_pipeline.pipeline_registers.registers[18][2] ),
    .A1(\core_pipeline.pipeline_registers.registers[19][2] ),
    .S(net556),
    .X(_04998_));
 sky130_fd_sc_hd__a22o_1 _08946_ (.A1(\core_pipeline.pipeline_registers.registers[16][2] ),
    .A2(net278),
    .B1(net361),
    .B2(_04998_),
    .X(_04999_));
 sky130_fd_sc_hd__a211o_1 _08947_ (.A1(\core_pipeline.pipeline_registers.registers[17][2] ),
    .A2(net276),
    .B1(_04999_),
    .C1(net460),
    .X(_05000_));
 sky130_fd_sc_hd__a211o_1 _08948_ (.A1(net370),
    .A2(_04997_),
    .B1(_05000_),
    .C1(_04996_),
    .X(_05001_));
 sky130_fd_sc_hd__and3_2 _08949_ (.A(net145),
    .B(_04989_),
    .C(_05001_),
    .X(_05002_));
 sky130_fd_sc_hd__a21o_1 _08950_ (.A1(\core_pipeline.decode_to_execute_rs2_data[2] ),
    .A2(net130),
    .B1(_05002_),
    .X(_00534_));
 sky130_fd_sc_hd__mux4_1 _08951_ (.A0(\core_pipeline.pipeline_registers.registers[8][3] ),
    .A1(\core_pipeline.pipeline_registers.registers[9][3] ),
    .A2(\core_pipeline.pipeline_registers.registers[10][3] ),
    .A3(\core_pipeline.pipeline_registers.registers[11][3] ),
    .S0(net548),
    .S1(net529),
    .X(_05003_));
 sky130_fd_sc_hd__or2_1 _08952_ (.A(net520),
    .B(_05003_),
    .X(_05004_));
 sky130_fd_sc_hd__mux4_1 _08953_ (.A0(\core_pipeline.pipeline_registers.registers[12][3] ),
    .A1(\core_pipeline.pipeline_registers.registers[13][3] ),
    .A2(\core_pipeline.pipeline_registers.registers[14][3] ),
    .A3(\core_pipeline.pipeline_registers.registers[15][3] ),
    .S0(net548),
    .S1(net529),
    .X(_05005_));
 sky130_fd_sc_hd__o211a_1 _08954_ (.A1(net462),
    .A2(_05005_),
    .B1(_05004_),
    .C1(net514),
    .X(_05006_));
 sky130_fd_sc_hd__mux4_1 _08955_ (.A0(\core_pipeline.pipeline_registers.registers[4][3] ),
    .A1(\core_pipeline.pipeline_registers.registers[5][3] ),
    .A2(\core_pipeline.pipeline_registers.registers[6][3] ),
    .A3(\core_pipeline.pipeline_registers.registers[7][3] ),
    .S0(net548),
    .S1(net529),
    .X(_05007_));
 sky130_fd_sc_hd__mux2_1 _08956_ (.A0(\core_pipeline.pipeline_registers.registers[2][3] ),
    .A1(\core_pipeline.pipeline_registers.registers[3][3] ),
    .S(net548),
    .X(_05008_));
 sky130_fd_sc_hd__a22o_1 _08957_ (.A1(\core_pipeline.pipeline_registers.registers[1][3] ),
    .A2(net277),
    .B1(net361),
    .B2(_05008_),
    .X(_05009_));
 sky130_fd_sc_hd__a211o_1 _08958_ (.A1(\core_pipeline.pipeline_registers.registers[0][3] ),
    .A2(net279),
    .B1(_05009_),
    .C1(net511),
    .X(_05010_));
 sky130_fd_sc_hd__a211o_1 _08959_ (.A1(net368),
    .A2(_05007_),
    .B1(_05010_),
    .C1(_05006_),
    .X(_05011_));
 sky130_fd_sc_hd__mux2_1 _08960_ (.A0(\core_pipeline.pipeline_registers.registers[30][3] ),
    .A1(\core_pipeline.pipeline_registers.registers[31][3] ),
    .S(net549),
    .X(_05012_));
 sky130_fd_sc_hd__a221o_1 _08961_ (.A1(\core_pipeline.pipeline_registers.registers[28][3] ),
    .A2(net424),
    .B1(net363),
    .B2(\core_pipeline.pipeline_registers.registers[29][3] ),
    .C1(net462),
    .X(_05013_));
 sky130_fd_sc_hd__a21o_1 _08962_ (.A1(net531),
    .A2(_05012_),
    .B1(_05013_),
    .X(_05014_));
 sky130_fd_sc_hd__mux2_1 _08963_ (.A0(\core_pipeline.pipeline_registers.registers[26][3] ),
    .A1(\core_pipeline.pipeline_registers.registers[27][3] ),
    .S(net549),
    .X(_05015_));
 sky130_fd_sc_hd__a221o_1 _08964_ (.A1(\core_pipeline.pipeline_registers.registers[24][3] ),
    .A2(net424),
    .B1(net363),
    .B2(\core_pipeline.pipeline_registers.registers[25][3] ),
    .C1(net519),
    .X(_05016_));
 sky130_fd_sc_hd__a21o_1 _08965_ (.A1(net531),
    .A2(_05015_),
    .B1(_05016_),
    .X(_05017_));
 sky130_fd_sc_hd__mux4_1 _08966_ (.A0(\core_pipeline.pipeline_registers.registers[16][3] ),
    .A1(\core_pipeline.pipeline_registers.registers[17][3] ),
    .A2(\core_pipeline.pipeline_registers.registers[18][3] ),
    .A3(\core_pipeline.pipeline_registers.registers[19][3] ),
    .S0(net551),
    .S1(net531),
    .X(_05018_));
 sky130_fd_sc_hd__mux4_1 _08967_ (.A0(\core_pipeline.pipeline_registers.registers[20][3] ),
    .A1(\core_pipeline.pipeline_registers.registers[21][3] ),
    .A2(\core_pipeline.pipeline_registers.registers[22][3] ),
    .A3(\core_pipeline.pipeline_registers.registers[23][3] ),
    .S0(net551),
    .S1(net531),
    .X(_05019_));
 sky130_fd_sc_hd__a22o_1 _08968_ (.A1(net429),
    .A2(_05018_),
    .B1(_05019_),
    .B2(net368),
    .X(_05020_));
 sky130_fd_sc_hd__a31o_1 _08969_ (.A1(net514),
    .A2(_05014_),
    .A3(_05017_),
    .B1(net461),
    .X(_05021_));
 sky130_fd_sc_hd__o21a_2 _08970_ (.A1(_05020_),
    .A2(_05021_),
    .B1(_05011_),
    .X(_05022_));
 sky130_fd_sc_hd__mux2_1 _08971_ (.A0(\core_pipeline.decode_to_execute_rs2_data[3] ),
    .A1(_05022_),
    .S(net141),
    .X(_00535_));
 sky130_fd_sc_hd__mux4_1 _08972_ (.A0(\core_pipeline.pipeline_registers.registers[12][4] ),
    .A1(\core_pipeline.pipeline_registers.registers[13][4] ),
    .A2(\core_pipeline.pipeline_registers.registers[14][4] ),
    .A3(\core_pipeline.pipeline_registers.registers[15][4] ),
    .S0(net544),
    .S1(net525),
    .X(_05023_));
 sky130_fd_sc_hd__mux4_1 _08973_ (.A0(\core_pipeline.pipeline_registers.registers[8][4] ),
    .A1(\core_pipeline.pipeline_registers.registers[9][4] ),
    .A2(\core_pipeline.pipeline_registers.registers[10][4] ),
    .A3(\core_pipeline.pipeline_registers.registers[11][4] ),
    .S0(net544),
    .S1(net525),
    .X(_05024_));
 sky130_fd_sc_hd__or2_1 _08974_ (.A(net519),
    .B(_05024_),
    .X(_05025_));
 sky130_fd_sc_hd__o211a_1 _08975_ (.A1(net462),
    .A2(_05023_),
    .B1(_05025_),
    .C1(net514),
    .X(_05026_));
 sky130_fd_sc_hd__mux4_1 _08976_ (.A0(\core_pipeline.pipeline_registers.registers[4][4] ),
    .A1(\core_pipeline.pipeline_registers.registers[5][4] ),
    .A2(\core_pipeline.pipeline_registers.registers[6][4] ),
    .A3(\core_pipeline.pipeline_registers.registers[7][4] ),
    .S0(net544),
    .S1(net525),
    .X(_05027_));
 sky130_fd_sc_hd__mux4_1 _08977_ (.A0(\core_pipeline.pipeline_registers.registers[0][4] ),
    .A1(\core_pipeline.pipeline_registers.registers[1][4] ),
    .A2(\core_pipeline.pipeline_registers.registers[2][4] ),
    .A3(\core_pipeline.pipeline_registers.registers[3][4] ),
    .S0(net544),
    .S1(net525),
    .X(_05028_));
 sky130_fd_sc_hd__a221o_1 _08978_ (.A1(net367),
    .A2(_05027_),
    .B1(_05028_),
    .B2(net428),
    .C1(net511),
    .X(_05029_));
 sky130_fd_sc_hd__mux2_1 _08979_ (.A0(\core_pipeline.pipeline_registers.registers[30][4] ),
    .A1(\core_pipeline.pipeline_registers.registers[31][4] ),
    .S(net548),
    .X(_05030_));
 sky130_fd_sc_hd__a221o_1 _08980_ (.A1(\core_pipeline.pipeline_registers.registers[28][4] ),
    .A2(net424),
    .B1(net363),
    .B2(\core_pipeline.pipeline_registers.registers[29][4] ),
    .C1(net462),
    .X(_05031_));
 sky130_fd_sc_hd__a21o_1 _08981_ (.A1(net528),
    .A2(_05030_),
    .B1(_05031_),
    .X(_05032_));
 sky130_fd_sc_hd__mux2_1 _08982_ (.A0(\core_pipeline.pipeline_registers.registers[26][4] ),
    .A1(\core_pipeline.pipeline_registers.registers[27][4] ),
    .S(net545),
    .X(_05033_));
 sky130_fd_sc_hd__a221o_1 _08983_ (.A1(\core_pipeline.pipeline_registers.registers[24][4] ),
    .A2(net424),
    .B1(net363),
    .B2(\core_pipeline.pipeline_registers.registers[25][4] ),
    .C1(net519),
    .X(_05034_));
 sky130_fd_sc_hd__a21o_1 _08984_ (.A1(net528),
    .A2(_05033_),
    .B1(_05034_),
    .X(_05035_));
 sky130_fd_sc_hd__and3_1 _08985_ (.A(net514),
    .B(_05032_),
    .C(_05035_),
    .X(_05036_));
 sky130_fd_sc_hd__mux4_1 _08986_ (.A0(\core_pipeline.pipeline_registers.registers[20][4] ),
    .A1(\core_pipeline.pipeline_registers.registers[21][4] ),
    .A2(\core_pipeline.pipeline_registers.registers[22][4] ),
    .A3(\core_pipeline.pipeline_registers.registers[23][4] ),
    .S0(net545),
    .S1(net528),
    .X(_05037_));
 sky130_fd_sc_hd__mux2_1 _08987_ (.A0(\core_pipeline.pipeline_registers.registers[18][4] ),
    .A1(\core_pipeline.pipeline_registers.registers[19][4] ),
    .S(net545),
    .X(_05038_));
 sky130_fd_sc_hd__a31o_1 _08988_ (.A1(net528),
    .A2(net428),
    .A3(_05038_),
    .B1(net461),
    .X(_05039_));
 sky130_fd_sc_hd__a221o_1 _08989_ (.A1(\core_pipeline.pipeline_registers.registers[16][4] ),
    .A2(net279),
    .B1(net277),
    .B2(\core_pipeline.pipeline_registers.registers[17][4] ),
    .C1(_05039_),
    .X(_05040_));
 sky130_fd_sc_hd__a21o_1 _08990_ (.A1(net367),
    .A2(_05037_),
    .B1(_05040_),
    .X(_05041_));
 sky130_fd_sc_hd__o22a_2 _08991_ (.A1(_05026_),
    .A2(_05029_),
    .B1(_05036_),
    .B2(_05041_),
    .X(_05042_));
 sky130_fd_sc_hd__mux2_1 _08992_ (.A0(\core_pipeline.decode_to_execute_rs2_data[4] ),
    .A1(_05042_),
    .S(net139),
    .X(_00536_));
 sky130_fd_sc_hd__mux4_1 _08993_ (.A0(\core_pipeline.pipeline_registers.registers[8][5] ),
    .A1(\core_pipeline.pipeline_registers.registers[9][5] ),
    .A2(\core_pipeline.pipeline_registers.registers[10][5] ),
    .A3(\core_pipeline.pipeline_registers.registers[11][5] ),
    .S0(net556),
    .S1(net534),
    .X(_05043_));
 sky130_fd_sc_hd__or2_1 _08994_ (.A(net522),
    .B(_05043_),
    .X(_05044_));
 sky130_fd_sc_hd__mux4_1 _08995_ (.A0(\core_pipeline.pipeline_registers.registers[12][5] ),
    .A1(\core_pipeline.pipeline_registers.registers[13][5] ),
    .A2(\core_pipeline.pipeline_registers.registers[14][5] ),
    .A3(\core_pipeline.pipeline_registers.registers[15][5] ),
    .S0(net556),
    .S1(net536),
    .X(_05045_));
 sky130_fd_sc_hd__o211a_1 _08996_ (.A1(net464),
    .A2(_05045_),
    .B1(_05044_),
    .C1(net516),
    .X(_05046_));
 sky130_fd_sc_hd__mux4_1 _08997_ (.A0(\core_pipeline.pipeline_registers.registers[4][5] ),
    .A1(\core_pipeline.pipeline_registers.registers[5][5] ),
    .A2(\core_pipeline.pipeline_registers.registers[6][5] ),
    .A3(\core_pipeline.pipeline_registers.registers[7][5] ),
    .S0(net556),
    .S1(net534),
    .X(_05047_));
 sky130_fd_sc_hd__mux2_1 _08998_ (.A0(\core_pipeline.pipeline_registers.registers[2][5] ),
    .A1(\core_pipeline.pipeline_registers.registers[3][5] ),
    .S(net556),
    .X(_05048_));
 sky130_fd_sc_hd__a22o_1 _08999_ (.A1(\core_pipeline.pipeline_registers.registers[1][5] ),
    .A2(net276),
    .B1(net361),
    .B2(_05048_),
    .X(_05049_));
 sky130_fd_sc_hd__a211o_1 _09000_ (.A1(\core_pipeline.pipeline_registers.registers[0][5] ),
    .A2(net278),
    .B1(_05049_),
    .C1(net512),
    .X(_05050_));
 sky130_fd_sc_hd__a211o_1 _09001_ (.A1(net370),
    .A2(_05047_),
    .B1(_05050_),
    .C1(_05046_),
    .X(_05051_));
 sky130_fd_sc_hd__mux2_1 _09002_ (.A0(\core_pipeline.pipeline_registers.registers[30][5] ),
    .A1(\core_pipeline.pipeline_registers.registers[31][5] ),
    .S(net556),
    .X(_05052_));
 sky130_fd_sc_hd__a221o_1 _09003_ (.A1(\core_pipeline.pipeline_registers.registers[28][5] ),
    .A2(net426),
    .B1(net365),
    .B2(\core_pipeline.pipeline_registers.registers[29][5] ),
    .C1(net464),
    .X(_05053_));
 sky130_fd_sc_hd__a21o_1 _09004_ (.A1(net534),
    .A2(_05052_),
    .B1(_05053_),
    .X(_05054_));
 sky130_fd_sc_hd__mux2_1 _09005_ (.A0(\core_pipeline.pipeline_registers.registers[26][5] ),
    .A1(\core_pipeline.pipeline_registers.registers[27][5] ),
    .S(net556),
    .X(_05055_));
 sky130_fd_sc_hd__a221o_1 _09006_ (.A1(\core_pipeline.pipeline_registers.registers[24][5] ),
    .A2(net426),
    .B1(net365),
    .B2(\core_pipeline.pipeline_registers.registers[25][5] ),
    .C1(net522),
    .X(_05056_));
 sky130_fd_sc_hd__a21o_1 _09007_ (.A1(net536),
    .A2(_05055_),
    .B1(_05056_),
    .X(_05057_));
 sky130_fd_sc_hd__and3_1 _09008_ (.A(net516),
    .B(_05054_),
    .C(_05057_),
    .X(_05058_));
 sky130_fd_sc_hd__mux4_1 _09009_ (.A0(\core_pipeline.pipeline_registers.registers[20][5] ),
    .A1(\core_pipeline.pipeline_registers.registers[21][5] ),
    .A2(\core_pipeline.pipeline_registers.registers[22][5] ),
    .A3(\core_pipeline.pipeline_registers.registers[23][5] ),
    .S0(net556),
    .S1(net536),
    .X(_05059_));
 sky130_fd_sc_hd__mux2_1 _09010_ (.A0(\core_pipeline.pipeline_registers.registers[18][5] ),
    .A1(\core_pipeline.pipeline_registers.registers[19][5] ),
    .S(net555),
    .X(_05060_));
 sky130_fd_sc_hd__a22o_1 _09011_ (.A1(\core_pipeline.pipeline_registers.registers[16][5] ),
    .A2(net278),
    .B1(net362),
    .B2(_05060_),
    .X(_05061_));
 sky130_fd_sc_hd__a211o_1 _09012_ (.A1(\core_pipeline.pipeline_registers.registers[17][5] ),
    .A2(net276),
    .B1(_05061_),
    .C1(net460),
    .X(_05062_));
 sky130_fd_sc_hd__a211o_1 _09013_ (.A1(net370),
    .A2(_05059_),
    .B1(_05062_),
    .C1(_05058_),
    .X(_05063_));
 sky130_fd_sc_hd__and3_4 _09014_ (.A(net145),
    .B(_05051_),
    .C(_05063_),
    .X(_05064_));
 sky130_fd_sc_hd__a21o_1 _09015_ (.A1(\core_pipeline.decode_to_execute_rs2_data[5] ),
    .A2(net130),
    .B1(_05064_),
    .X(_00537_));
 sky130_fd_sc_hd__mux4_1 _09016_ (.A0(\core_pipeline.pipeline_registers.registers[8][6] ),
    .A1(\core_pipeline.pipeline_registers.registers[9][6] ),
    .A2(\core_pipeline.pipeline_registers.registers[10][6] ),
    .A3(\core_pipeline.pipeline_registers.registers[11][6] ),
    .S0(net555),
    .S1(net534),
    .X(_05065_));
 sky130_fd_sc_hd__or2_1 _09017_ (.A(net522),
    .B(_05065_),
    .X(_05066_));
 sky130_fd_sc_hd__mux4_1 _09018_ (.A0(\core_pipeline.pipeline_registers.registers[12][6] ),
    .A1(\core_pipeline.pipeline_registers.registers[13][6] ),
    .A2(\core_pipeline.pipeline_registers.registers[14][6] ),
    .A3(\core_pipeline.pipeline_registers.registers[15][6] ),
    .S0(net549),
    .S1(net529),
    .X(_05067_));
 sky130_fd_sc_hd__o211a_1 _09019_ (.A1(net464),
    .A2(_05067_),
    .B1(_05066_),
    .C1(net516),
    .X(_05068_));
 sky130_fd_sc_hd__mux4_1 _09020_ (.A0(\core_pipeline.pipeline_registers.registers[4][6] ),
    .A1(\core_pipeline.pipeline_registers.registers[5][6] ),
    .A2(\core_pipeline.pipeline_registers.registers[6][6] ),
    .A3(\core_pipeline.pipeline_registers.registers[7][6] ),
    .S0(net549),
    .S1(net529),
    .X(_05069_));
 sky130_fd_sc_hd__mux2_1 _09021_ (.A0(\core_pipeline.pipeline_registers.registers[2][6] ),
    .A1(\core_pipeline.pipeline_registers.registers[3][6] ),
    .S(net549),
    .X(_05070_));
 sky130_fd_sc_hd__a22o_1 _09022_ (.A1(\core_pipeline.pipeline_registers.registers[1][6] ),
    .A2(net277),
    .B1(net361),
    .B2(_05070_),
    .X(_05071_));
 sky130_fd_sc_hd__a211o_1 _09023_ (.A1(\core_pipeline.pipeline_registers.registers[0][6] ),
    .A2(net279),
    .B1(_05071_),
    .C1(net511),
    .X(_05072_));
 sky130_fd_sc_hd__a211o_1 _09024_ (.A1(net368),
    .A2(_05069_),
    .B1(_05072_),
    .C1(_05068_),
    .X(_05073_));
 sky130_fd_sc_hd__mux2_1 _09025_ (.A0(\core_pipeline.pipeline_registers.registers[26][6] ),
    .A1(\core_pipeline.pipeline_registers.registers[27][6] ),
    .S(net555),
    .X(_05074_));
 sky130_fd_sc_hd__a221o_1 _09026_ (.A1(\core_pipeline.pipeline_registers.registers[24][6] ),
    .A2(net424),
    .B1(net363),
    .B2(\core_pipeline.pipeline_registers.registers[25][6] ),
    .C1(net522),
    .X(_05075_));
 sky130_fd_sc_hd__a21o_1 _09027_ (.A1(net534),
    .A2(_05074_),
    .B1(_05075_),
    .X(_05076_));
 sky130_fd_sc_hd__mux2_1 _09028_ (.A0(\core_pipeline.pipeline_registers.registers[30][6] ),
    .A1(\core_pipeline.pipeline_registers.registers[31][6] ),
    .S(net555),
    .X(_05077_));
 sky130_fd_sc_hd__a221o_1 _09029_ (.A1(\core_pipeline.pipeline_registers.registers[28][6] ),
    .A2(net426),
    .B1(net365),
    .B2(\core_pipeline.pipeline_registers.registers[29][6] ),
    .C1(net464),
    .X(_05078_));
 sky130_fd_sc_hd__a21o_1 _09030_ (.A1(net534),
    .A2(_05077_),
    .B1(_05078_),
    .X(_05079_));
 sky130_fd_sc_hd__mux4_1 _09031_ (.A0(\core_pipeline.pipeline_registers.registers[16][6] ),
    .A1(\core_pipeline.pipeline_registers.registers[17][6] ),
    .A2(\core_pipeline.pipeline_registers.registers[18][6] ),
    .A3(\core_pipeline.pipeline_registers.registers[19][6] ),
    .S0(net555),
    .S1(net534),
    .X(_05080_));
 sky130_fd_sc_hd__mux4_1 _09032_ (.A0(\core_pipeline.pipeline_registers.registers[20][6] ),
    .A1(\core_pipeline.pipeline_registers.registers[21][6] ),
    .A2(\core_pipeline.pipeline_registers.registers[22][6] ),
    .A3(\core_pipeline.pipeline_registers.registers[23][6] ),
    .S0(net555),
    .S1(net534),
    .X(_05081_));
 sky130_fd_sc_hd__a22o_1 _09033_ (.A1(net430),
    .A2(_05080_),
    .B1(_05081_),
    .B2(net370),
    .X(_05082_));
 sky130_fd_sc_hd__a31o_1 _09034_ (.A1(net516),
    .A2(_05076_),
    .A3(_05079_),
    .B1(net460),
    .X(_05083_));
 sky130_fd_sc_hd__o211a_2 _09035_ (.A1(_05082_),
    .A2(_05083_),
    .B1(net144),
    .C1(_05073_),
    .X(_05084_));
 sky130_fd_sc_hd__a21o_1 _09036_ (.A1(\core_pipeline.decode_to_execute_rs2_data[6] ),
    .A2(net125),
    .B1(_05084_),
    .X(_00538_));
 sky130_fd_sc_hd__mux4_1 _09037_ (.A0(\core_pipeline.pipeline_registers.registers[8][7] ),
    .A1(\core_pipeline.pipeline_registers.registers[9][7] ),
    .A2(\core_pipeline.pipeline_registers.registers[10][7] ),
    .A3(\core_pipeline.pipeline_registers.registers[11][7] ),
    .S0(net544),
    .S1(net525),
    .X(_05085_));
 sky130_fd_sc_hd__or2_1 _09038_ (.A(net519),
    .B(_05085_),
    .X(_05086_));
 sky130_fd_sc_hd__mux4_1 _09039_ (.A0(\core_pipeline.pipeline_registers.registers[12][7] ),
    .A1(\core_pipeline.pipeline_registers.registers[13][7] ),
    .A2(\core_pipeline.pipeline_registers.registers[14][7] ),
    .A3(\core_pipeline.pipeline_registers.registers[15][7] ),
    .S0(net544),
    .S1(net525),
    .X(_05087_));
 sky130_fd_sc_hd__o211a_1 _09040_ (.A1(net462),
    .A2(_05087_),
    .B1(_05086_),
    .C1(net514),
    .X(_05088_));
 sky130_fd_sc_hd__mux4_2 _09041_ (.A0(\core_pipeline.pipeline_registers.registers[0][7] ),
    .A1(\core_pipeline.pipeline_registers.registers[1][7] ),
    .A2(\core_pipeline.pipeline_registers.registers[2][7] ),
    .A3(\core_pipeline.pipeline_registers.registers[3][7] ),
    .S0(net544),
    .S1(net525),
    .X(_05089_));
 sky130_fd_sc_hd__mux4_2 _09042_ (.A0(\core_pipeline.pipeline_registers.registers[4][7] ),
    .A1(\core_pipeline.pipeline_registers.registers[5][7] ),
    .A2(\core_pipeline.pipeline_registers.registers[6][7] ),
    .A3(\core_pipeline.pipeline_registers.registers[7][7] ),
    .S0(net544),
    .S1(net525),
    .X(_05090_));
 sky130_fd_sc_hd__a221o_4 _09043_ (.A1(net428),
    .A2(_05089_),
    .B1(_05090_),
    .B2(net367),
    .C1(_05088_),
    .X(_05091_));
 sky130_fd_sc_hd__mux2_1 _09044_ (.A0(\core_pipeline.pipeline_registers.registers[26][7] ),
    .A1(\core_pipeline.pipeline_registers.registers[27][7] ),
    .S(net551),
    .X(_05092_));
 sky130_fd_sc_hd__a221o_1 _09045_ (.A1(\core_pipeline.pipeline_registers.registers[24][7] ),
    .A2(net425),
    .B1(net364),
    .B2(\core_pipeline.pipeline_registers.registers[25][7] ),
    .C1(net520),
    .X(_05093_));
 sky130_fd_sc_hd__a21o_1 _09046_ (.A1(net530),
    .A2(_05092_),
    .B1(_05093_),
    .X(_05094_));
 sky130_fd_sc_hd__mux2_1 _09047_ (.A0(\core_pipeline.pipeline_registers.registers[30][7] ),
    .A1(\core_pipeline.pipeline_registers.registers[31][7] ),
    .S(net551),
    .X(_05095_));
 sky130_fd_sc_hd__a221o_1 _09048_ (.A1(\core_pipeline.pipeline_registers.registers[28][7] ),
    .A2(net425),
    .B1(net364),
    .B2(\core_pipeline.pipeline_registers.registers[29][7] ),
    .C1(net462),
    .X(_05096_));
 sky130_fd_sc_hd__a21o_1 _09049_ (.A1(net530),
    .A2(_05095_),
    .B1(_05096_),
    .X(_05097_));
 sky130_fd_sc_hd__mux4_1 _09050_ (.A0(\core_pipeline.pipeline_registers.registers[16][7] ),
    .A1(\core_pipeline.pipeline_registers.registers[17][7] ),
    .A2(\core_pipeline.pipeline_registers.registers[18][7] ),
    .A3(\core_pipeline.pipeline_registers.registers[19][7] ),
    .S0(net550),
    .S1(net530),
    .X(_05098_));
 sky130_fd_sc_hd__mux4_1 _09051_ (.A0(\core_pipeline.pipeline_registers.registers[20][7] ),
    .A1(\core_pipeline.pipeline_registers.registers[21][7] ),
    .A2(\core_pipeline.pipeline_registers.registers[22][7] ),
    .A3(\core_pipeline.pipeline_registers.registers[23][7] ),
    .S0(net550),
    .S1(net530),
    .X(_05099_));
 sky130_fd_sc_hd__a22o_1 _09052_ (.A1(net429),
    .A2(_05098_),
    .B1(_05099_),
    .B2(net368),
    .X(_05100_));
 sky130_fd_sc_hd__a31o_1 _09053_ (.A1(net514),
    .A2(_05094_),
    .A3(_05097_),
    .B1(net461),
    .X(_05101_));
 sky130_fd_sc_hd__o22a_2 _09054_ (.A1(net511),
    .A2(_05091_),
    .B1(_05100_),
    .B2(_05101_),
    .X(_05102_));
 sky130_fd_sc_hd__mux2_1 _09055_ (.A0(\core_pipeline.decode_to_execute_rs2_data[7] ),
    .A1(_05102_),
    .S(net142),
    .X(_00539_));
 sky130_fd_sc_hd__mux2_1 _09056_ (.A0(\core_pipeline.pipeline_registers.registers[30][8] ),
    .A1(\core_pipeline.pipeline_registers.registers[31][8] ),
    .S(net548),
    .X(_05103_));
 sky130_fd_sc_hd__a221o_1 _09057_ (.A1(\core_pipeline.pipeline_registers.registers[28][8] ),
    .A2(net424),
    .B1(net364),
    .B2(\core_pipeline.pipeline_registers.registers[29][8] ),
    .C1(net462),
    .X(_05104_));
 sky130_fd_sc_hd__a21o_1 _09058_ (.A1(net531),
    .A2(_05103_),
    .B1(_05104_),
    .X(_05105_));
 sky130_fd_sc_hd__mux2_1 _09059_ (.A0(\core_pipeline.pipeline_registers.registers[26][8] ),
    .A1(\core_pipeline.pipeline_registers.registers[27][8] ),
    .S(net548),
    .X(_05106_));
 sky130_fd_sc_hd__a221o_1 _09060_ (.A1(\core_pipeline.pipeline_registers.registers[24][8] ),
    .A2(net425),
    .B1(net364),
    .B2(\core_pipeline.pipeline_registers.registers[25][8] ),
    .C1(net520),
    .X(_05107_));
 sky130_fd_sc_hd__a21o_1 _09061_ (.A1(net529),
    .A2(_05106_),
    .B1(_05107_),
    .X(_05108_));
 sky130_fd_sc_hd__and3_1 _09062_ (.A(net515),
    .B(_05105_),
    .C(_05108_),
    .X(_05109_));
 sky130_fd_sc_hd__mux4_1 _09063_ (.A0(\core_pipeline.pipeline_registers.registers[20][8] ),
    .A1(\core_pipeline.pipeline_registers.registers[21][8] ),
    .A2(\core_pipeline.pipeline_registers.registers[22][8] ),
    .A3(\core_pipeline.pipeline_registers.registers[23][8] ),
    .S0(net548),
    .S1(net529),
    .X(_05110_));
 sky130_fd_sc_hd__mux2_1 _09064_ (.A0(\core_pipeline.pipeline_registers.registers[18][8] ),
    .A1(\core_pipeline.pipeline_registers.registers[19][8] ),
    .S(net548),
    .X(_05111_));
 sky130_fd_sc_hd__a22o_1 _09065_ (.A1(\core_pipeline.pipeline_registers.registers[17][8] ),
    .A2(net277),
    .B1(net361),
    .B2(_05111_),
    .X(_05112_));
 sky130_fd_sc_hd__a211o_1 _09066_ (.A1(\core_pipeline.pipeline_registers.registers[16][8] ),
    .A2(net279),
    .B1(_05112_),
    .C1(net461),
    .X(_05113_));
 sky130_fd_sc_hd__a211o_1 _09067_ (.A1(net368),
    .A2(_05110_),
    .B1(_05113_),
    .C1(_05109_),
    .X(_05114_));
 sky130_fd_sc_hd__mux4_1 _09068_ (.A0(\core_pipeline.pipeline_registers.registers[12][8] ),
    .A1(\core_pipeline.pipeline_registers.registers[13][8] ),
    .A2(\core_pipeline.pipeline_registers.registers[14][8] ),
    .A3(\core_pipeline.pipeline_registers.registers[15][8] ),
    .S0(net549),
    .S1(net529),
    .X(_05115_));
 sky130_fd_sc_hd__mux4_1 _09069_ (.A0(\core_pipeline.pipeline_registers.registers[8][8] ),
    .A1(\core_pipeline.pipeline_registers.registers[9][8] ),
    .A2(\core_pipeline.pipeline_registers.registers[10][8] ),
    .A3(\core_pipeline.pipeline_registers.registers[11][8] ),
    .S0(net549),
    .S1(net529),
    .X(_05116_));
 sky130_fd_sc_hd__or2_1 _09070_ (.A(net520),
    .B(_05116_),
    .X(_05117_));
 sky130_fd_sc_hd__o211a_1 _09071_ (.A1(net462),
    .A2(_05115_),
    .B1(_05117_),
    .C1(net514),
    .X(_05118_));
 sky130_fd_sc_hd__mux4_1 _09072_ (.A0(\core_pipeline.pipeline_registers.registers[4][8] ),
    .A1(\core_pipeline.pipeline_registers.registers[5][8] ),
    .A2(\core_pipeline.pipeline_registers.registers[6][8] ),
    .A3(\core_pipeline.pipeline_registers.registers[7][8] ),
    .S0(net549),
    .S1(net531),
    .X(_05119_));
 sky130_fd_sc_hd__mux2_1 _09073_ (.A0(\core_pipeline.pipeline_registers.registers[2][8] ),
    .A1(\core_pipeline.pipeline_registers.registers[3][8] ),
    .S(net549),
    .X(_05120_));
 sky130_fd_sc_hd__a221o_1 _09074_ (.A1(\core_pipeline.pipeline_registers.registers[0][8] ),
    .A2(net279),
    .B1(net277),
    .B2(\core_pipeline.pipeline_registers.registers[1][8] ),
    .C1(net511),
    .X(_05121_));
 sky130_fd_sc_hd__a21o_1 _09075_ (.A1(net368),
    .A2(_05119_),
    .B1(_05121_),
    .X(_05122_));
 sky130_fd_sc_hd__a211o_1 _09076_ (.A1(net361),
    .A2(_05120_),
    .B1(_05122_),
    .C1(_05118_),
    .X(_05123_));
 sky130_fd_sc_hd__and3_2 _09077_ (.A(net144),
    .B(_05114_),
    .C(_05123_),
    .X(_05124_));
 sky130_fd_sc_hd__a21o_1 _09078_ (.A1(\core_pipeline.decode_to_execute_rs2_data[8] ),
    .A2(net124),
    .B1(_05124_),
    .X(_00540_));
 sky130_fd_sc_hd__mux4_1 _09079_ (.A0(\core_pipeline.pipeline_registers.registers[8][9] ),
    .A1(\core_pipeline.pipeline_registers.registers[9][9] ),
    .A2(\core_pipeline.pipeline_registers.registers[10][9] ),
    .A3(\core_pipeline.pipeline_registers.registers[11][9] ),
    .S0(net546),
    .S1(net526),
    .X(_05125_));
 sky130_fd_sc_hd__or2_1 _09080_ (.A(net519),
    .B(_05125_),
    .X(_05126_));
 sky130_fd_sc_hd__mux4_1 _09081_ (.A0(\core_pipeline.pipeline_registers.registers[12][9] ),
    .A1(\core_pipeline.pipeline_registers.registers[13][9] ),
    .A2(\core_pipeline.pipeline_registers.registers[14][9] ),
    .A3(\core_pipeline.pipeline_registers.registers[15][9] ),
    .S0(net546),
    .S1(net526),
    .X(_05127_));
 sky130_fd_sc_hd__o211a_1 _09082_ (.A1(net463),
    .A2(_05127_),
    .B1(_05126_),
    .C1(net514),
    .X(_05128_));
 sky130_fd_sc_hd__mux4_1 _09083_ (.A0(\core_pipeline.pipeline_registers.registers[0][9] ),
    .A1(\core_pipeline.pipeline_registers.registers[1][9] ),
    .A2(\core_pipeline.pipeline_registers.registers[2][9] ),
    .A3(\core_pipeline.pipeline_registers.registers[3][9] ),
    .S0(net546),
    .S1(net526),
    .X(_05129_));
 sky130_fd_sc_hd__mux4_1 _09084_ (.A0(\core_pipeline.pipeline_registers.registers[4][9] ),
    .A1(\core_pipeline.pipeline_registers.registers[5][9] ),
    .A2(\core_pipeline.pipeline_registers.registers[6][9] ),
    .A3(\core_pipeline.pipeline_registers.registers[7][9] ),
    .S0(net546),
    .S1(net526),
    .X(_05130_));
 sky130_fd_sc_hd__a221o_2 _09085_ (.A1(net428),
    .A2(_05129_),
    .B1(_05130_),
    .B2(net367),
    .C1(_05128_),
    .X(_05131_));
 sky130_fd_sc_hd__mux2_1 _09086_ (.A0(\core_pipeline.pipeline_registers.registers[26][9] ),
    .A1(\core_pipeline.pipeline_registers.registers[27][9] ),
    .S(net546),
    .X(_05132_));
 sky130_fd_sc_hd__a221o_1 _09087_ (.A1(\core_pipeline.pipeline_registers.registers[24][9] ),
    .A2(net424),
    .B1(net363),
    .B2(\core_pipeline.pipeline_registers.registers[25][9] ),
    .C1(net519),
    .X(_05133_));
 sky130_fd_sc_hd__a21o_1 _09088_ (.A1(net527),
    .A2(_05132_),
    .B1(_05133_),
    .X(_05134_));
 sky130_fd_sc_hd__mux2_1 _09089_ (.A0(\core_pipeline.pipeline_registers.registers[30][9] ),
    .A1(\core_pipeline.pipeline_registers.registers[31][9] ),
    .S(net550),
    .X(_05135_));
 sky130_fd_sc_hd__a221o_1 _09090_ (.A1(\core_pipeline.pipeline_registers.registers[28][9] ),
    .A2(net424),
    .B1(net363),
    .B2(\core_pipeline.pipeline_registers.registers[29][9] ),
    .C1(net463),
    .X(_05136_));
 sky130_fd_sc_hd__a21o_1 _09091_ (.A1(net526),
    .A2(_05135_),
    .B1(_05136_),
    .X(_05137_));
 sky130_fd_sc_hd__mux4_1 _09092_ (.A0(\core_pipeline.pipeline_registers.registers[16][9] ),
    .A1(\core_pipeline.pipeline_registers.registers[17][9] ),
    .A2(\core_pipeline.pipeline_registers.registers[18][9] ),
    .A3(\core_pipeline.pipeline_registers.registers[19][9] ),
    .S0(net546),
    .S1(net526),
    .X(_05138_));
 sky130_fd_sc_hd__mux4_1 _09093_ (.A0(\core_pipeline.pipeline_registers.registers[20][9] ),
    .A1(\core_pipeline.pipeline_registers.registers[21][9] ),
    .A2(\core_pipeline.pipeline_registers.registers[22][9] ),
    .A3(\core_pipeline.pipeline_registers.registers[23][9] ),
    .S0(net547),
    .S1(net527),
    .X(_05139_));
 sky130_fd_sc_hd__a22o_1 _09094_ (.A1(net428),
    .A2(_05138_),
    .B1(_05139_),
    .B2(net367),
    .X(_05140_));
 sky130_fd_sc_hd__a31o_1 _09095_ (.A1(net514),
    .A2(_05134_),
    .A3(_05137_),
    .B1(net461),
    .X(_05141_));
 sky130_fd_sc_hd__o22a_1 _09096_ (.A1(net511),
    .A2(_05131_),
    .B1(_05140_),
    .B2(_05141_),
    .X(_05142_));
 sky130_fd_sc_hd__mux2_1 _09097_ (.A0(\core_pipeline.decode_to_execute_rs2_data[9] ),
    .A1(_05142_),
    .S(net139),
    .X(_00541_));
 sky130_fd_sc_hd__mux4_1 _09098_ (.A0(\core_pipeline.pipeline_registers.registers[8][10] ),
    .A1(\core_pipeline.pipeline_registers.registers[9][10] ),
    .A2(\core_pipeline.pipeline_registers.registers[10][10] ),
    .A3(\core_pipeline.pipeline_registers.registers[11][10] ),
    .S0(net552),
    .S1(net532),
    .X(_05143_));
 sky130_fd_sc_hd__or2_1 _09099_ (.A(net521),
    .B(_05143_),
    .X(_05144_));
 sky130_fd_sc_hd__mux4_1 _09100_ (.A0(\core_pipeline.pipeline_registers.registers[12][10] ),
    .A1(\core_pipeline.pipeline_registers.registers[13][10] ),
    .A2(\core_pipeline.pipeline_registers.registers[14][10] ),
    .A3(\core_pipeline.pipeline_registers.registers[15][10] ),
    .S0(net552),
    .S1(net532),
    .X(_05145_));
 sky130_fd_sc_hd__o211a_1 _09101_ (.A1(net463),
    .A2(_05145_),
    .B1(_05144_),
    .C1(net515),
    .X(_05146_));
 sky130_fd_sc_hd__mux4_2 _09102_ (.A0(\core_pipeline.pipeline_registers.registers[0][10] ),
    .A1(\core_pipeline.pipeline_registers.registers[1][10] ),
    .A2(\core_pipeline.pipeline_registers.registers[2][10] ),
    .A3(\core_pipeline.pipeline_registers.registers[3][10] ),
    .S0(net554),
    .S1(net533),
    .X(_05147_));
 sky130_fd_sc_hd__mux4_2 _09103_ (.A0(\core_pipeline.pipeline_registers.registers[4][10] ),
    .A1(\core_pipeline.pipeline_registers.registers[5][10] ),
    .A2(\core_pipeline.pipeline_registers.registers[6][10] ),
    .A3(\core_pipeline.pipeline_registers.registers[7][10] ),
    .S0(net552),
    .S1(net533),
    .X(_05148_));
 sky130_fd_sc_hd__a221o_2 _09104_ (.A1(net428),
    .A2(_05147_),
    .B1(_05148_),
    .B2(net367),
    .C1(_05146_),
    .X(_05149_));
 sky130_fd_sc_hd__mux2_1 _09105_ (.A0(\core_pipeline.pipeline_registers.registers[30][10] ),
    .A1(\core_pipeline.pipeline_registers.registers[31][10] ),
    .S(net547),
    .X(_05150_));
 sky130_fd_sc_hd__a221o_1 _09106_ (.A1(\core_pipeline.pipeline_registers.registers[28][10] ),
    .A2(net425),
    .B1(net364),
    .B2(\core_pipeline.pipeline_registers.registers[29][10] ),
    .C1(net463),
    .X(_05151_));
 sky130_fd_sc_hd__a21o_1 _09107_ (.A1(net527),
    .A2(_05150_),
    .B1(_05151_),
    .X(_05152_));
 sky130_fd_sc_hd__mux2_1 _09108_ (.A0(\core_pipeline.pipeline_registers.registers[26][10] ),
    .A1(\core_pipeline.pipeline_registers.registers[27][10] ),
    .S(net547),
    .X(_05153_));
 sky130_fd_sc_hd__a221o_1 _09109_ (.A1(\core_pipeline.pipeline_registers.registers[24][10] ),
    .A2(net425),
    .B1(net364),
    .B2(\core_pipeline.pipeline_registers.registers[25][10] ),
    .C1(net519),
    .X(_05154_));
 sky130_fd_sc_hd__a21o_1 _09110_ (.A1(net527),
    .A2(_05153_),
    .B1(_05154_),
    .X(_05155_));
 sky130_fd_sc_hd__mux4_1 _09111_ (.A0(\core_pipeline.pipeline_registers.registers[16][10] ),
    .A1(\core_pipeline.pipeline_registers.registers[17][10] ),
    .A2(\core_pipeline.pipeline_registers.registers[18][10] ),
    .A3(\core_pipeline.pipeline_registers.registers[19][10] ),
    .S0(net546),
    .S1(net526),
    .X(_05156_));
 sky130_fd_sc_hd__mux4_1 _09112_ (.A0(\core_pipeline.pipeline_registers.registers[20][10] ),
    .A1(\core_pipeline.pipeline_registers.registers[21][10] ),
    .A2(\core_pipeline.pipeline_registers.registers[22][10] ),
    .A3(\core_pipeline.pipeline_registers.registers[23][10] ),
    .S0(net546),
    .S1(net526),
    .X(_05157_));
 sky130_fd_sc_hd__a22o_1 _09113_ (.A1(net428),
    .A2(_05156_),
    .B1(_05157_),
    .B2(net367),
    .X(_05158_));
 sky130_fd_sc_hd__a31o_1 _09114_ (.A1(net515),
    .A2(_05152_),
    .A3(_05155_),
    .B1(net461),
    .X(_05159_));
 sky130_fd_sc_hd__o22a_2 _09115_ (.A1(net511),
    .A2(_05149_),
    .B1(_05158_),
    .B2(_05159_),
    .X(_05160_));
 sky130_fd_sc_hd__mux2_1 _09116_ (.A0(\core_pipeline.decode_to_execute_rs2_data[10] ),
    .A1(_05160_),
    .S(net140),
    .X(_00542_));
 sky130_fd_sc_hd__mux4_1 _09117_ (.A0(\core_pipeline.pipeline_registers.registers[12][11] ),
    .A1(\core_pipeline.pipeline_registers.registers[13][11] ),
    .A2(\core_pipeline.pipeline_registers.registers[14][11] ),
    .A3(\core_pipeline.pipeline_registers.registers[15][11] ),
    .S0(net544),
    .S1(net525),
    .X(_05161_));
 sky130_fd_sc_hd__mux4_1 _09118_ (.A0(\core_pipeline.pipeline_registers.registers[8][11] ),
    .A1(\core_pipeline.pipeline_registers.registers[9][11] ),
    .A2(\core_pipeline.pipeline_registers.registers[10][11] ),
    .A3(\core_pipeline.pipeline_registers.registers[11][11] ),
    .S0(net544),
    .S1(net526),
    .X(_05162_));
 sky130_fd_sc_hd__or2_1 _09119_ (.A(net519),
    .B(_05162_),
    .X(_05163_));
 sky130_fd_sc_hd__o211a_1 _09120_ (.A1(net462),
    .A2(_05161_),
    .B1(_05163_),
    .C1(net514),
    .X(_05164_));
 sky130_fd_sc_hd__mux4_1 _09121_ (.A0(\core_pipeline.pipeline_registers.registers[0][11] ),
    .A1(\core_pipeline.pipeline_registers.registers[1][11] ),
    .A2(\core_pipeline.pipeline_registers.registers[2][11] ),
    .A3(\core_pipeline.pipeline_registers.registers[3][11] ),
    .S0(net546),
    .S1(net526),
    .X(_05165_));
 sky130_fd_sc_hd__mux4_1 _09122_ (.A0(\core_pipeline.pipeline_registers.registers[4][11] ),
    .A1(\core_pipeline.pipeline_registers.registers[5][11] ),
    .A2(\core_pipeline.pipeline_registers.registers[6][11] ),
    .A3(\core_pipeline.pipeline_registers.registers[7][11] ),
    .S0(net546),
    .S1(net526),
    .X(_05166_));
 sky130_fd_sc_hd__a221o_1 _09123_ (.A1(net428),
    .A2(_05165_),
    .B1(_05166_),
    .B2(net367),
    .C1(net511),
    .X(_05167_));
 sky130_fd_sc_hd__mux2_1 _09124_ (.A0(\core_pipeline.pipeline_registers.registers[30][11] ),
    .A1(\core_pipeline.pipeline_registers.registers[31][11] ),
    .S(net548),
    .X(_05168_));
 sky130_fd_sc_hd__a221o_1 _09125_ (.A1(\core_pipeline.pipeline_registers.registers[28][11] ),
    .A2(net424),
    .B1(net363),
    .B2(\core_pipeline.pipeline_registers.registers[29][11] ),
    .C1(net462),
    .X(_05169_));
 sky130_fd_sc_hd__a21o_1 _09126_ (.A1(net529),
    .A2(_05168_),
    .B1(_05169_),
    .X(_05170_));
 sky130_fd_sc_hd__mux2_1 _09127_ (.A0(\core_pipeline.pipeline_registers.registers[26][11] ),
    .A1(\core_pipeline.pipeline_registers.registers[27][11] ),
    .S(net548),
    .X(_05171_));
 sky130_fd_sc_hd__a221o_1 _09128_ (.A1(\core_pipeline.pipeline_registers.registers[24][11] ),
    .A2(net424),
    .B1(net363),
    .B2(\core_pipeline.pipeline_registers.registers[25][11] ),
    .C1(net519),
    .X(_05172_));
 sky130_fd_sc_hd__a21o_1 _09129_ (.A1(net529),
    .A2(_05171_),
    .B1(_05172_),
    .X(_05173_));
 sky130_fd_sc_hd__and3_1 _09130_ (.A(net514),
    .B(_05170_),
    .C(_05173_),
    .X(_05174_));
 sky130_fd_sc_hd__mux4_1 _09131_ (.A0(\core_pipeline.pipeline_registers.registers[20][11] ),
    .A1(\core_pipeline.pipeline_registers.registers[21][11] ),
    .A2(\core_pipeline.pipeline_registers.registers[22][11] ),
    .A3(\core_pipeline.pipeline_registers.registers[23][11] ),
    .S0(net544),
    .S1(net525),
    .X(_05175_));
 sky130_fd_sc_hd__mux2_1 _09132_ (.A0(\core_pipeline.pipeline_registers.registers[18][11] ),
    .A1(\core_pipeline.pipeline_registers.registers[19][11] ),
    .S(net545),
    .X(_05176_));
 sky130_fd_sc_hd__a31o_1 _09133_ (.A1(net526),
    .A2(net428),
    .A3(_05176_),
    .B1(net461),
    .X(_05177_));
 sky130_fd_sc_hd__a221o_1 _09134_ (.A1(\core_pipeline.pipeline_registers.registers[16][11] ),
    .A2(net279),
    .B1(net277),
    .B2(\core_pipeline.pipeline_registers.registers[17][11] ),
    .C1(_05177_),
    .X(_05178_));
 sky130_fd_sc_hd__a21o_1 _09135_ (.A1(net367),
    .A2(_05175_),
    .B1(_05178_),
    .X(_05179_));
 sky130_fd_sc_hd__o22a_2 _09136_ (.A1(_05164_),
    .A2(_05167_),
    .B1(_05174_),
    .B2(_05179_),
    .X(_05180_));
 sky130_fd_sc_hd__mux2_1 _09137_ (.A0(\core_pipeline.decode_to_execute_rs2_data[11] ),
    .A1(_05180_),
    .S(net139),
    .X(_00543_));
 sky130_fd_sc_hd__mux4_1 _09138_ (.A0(\core_pipeline.pipeline_registers.registers[8][12] ),
    .A1(\core_pipeline.pipeline_registers.registers[9][12] ),
    .A2(\core_pipeline.pipeline_registers.registers[10][12] ),
    .A3(\core_pipeline.pipeline_registers.registers[11][12] ),
    .S0(net547),
    .S1(net527),
    .X(_05181_));
 sky130_fd_sc_hd__or2_1 _09139_ (.A(net519),
    .B(_05181_),
    .X(_05182_));
 sky130_fd_sc_hd__mux4_1 _09140_ (.A0(\core_pipeline.pipeline_registers.registers[12][12] ),
    .A1(\core_pipeline.pipeline_registers.registers[13][12] ),
    .A2(\core_pipeline.pipeline_registers.registers[14][12] ),
    .A3(\core_pipeline.pipeline_registers.registers[15][12] ),
    .S0(net545),
    .S1(net527),
    .X(_05183_));
 sky130_fd_sc_hd__o211a_1 _09141_ (.A1(net462),
    .A2(_05183_),
    .B1(_05182_),
    .C1(net514),
    .X(_05184_));
 sky130_fd_sc_hd__mux4_1 _09142_ (.A0(\core_pipeline.pipeline_registers.registers[4][12] ),
    .A1(\core_pipeline.pipeline_registers.registers[5][12] ),
    .A2(\core_pipeline.pipeline_registers.registers[6][12] ),
    .A3(\core_pipeline.pipeline_registers.registers[7][12] ),
    .S0(net550),
    .S1(net530),
    .X(_05185_));
 sky130_fd_sc_hd__mux2_1 _09143_ (.A0(\core_pipeline.pipeline_registers.registers[2][12] ),
    .A1(\core_pipeline.pipeline_registers.registers[3][12] ),
    .S(net550),
    .X(_05186_));
 sky130_fd_sc_hd__a22o_1 _09144_ (.A1(\core_pipeline.pipeline_registers.registers[0][12] ),
    .A2(net279),
    .B1(net361),
    .B2(_05186_),
    .X(_05187_));
 sky130_fd_sc_hd__a211o_1 _09145_ (.A1(\core_pipeline.pipeline_registers.registers[1][12] ),
    .A2(net277),
    .B1(_05187_),
    .C1(net511),
    .X(_05188_));
 sky130_fd_sc_hd__a211o_1 _09146_ (.A1(net368),
    .A2(_05185_),
    .B1(_05188_),
    .C1(_05184_),
    .X(_05189_));
 sky130_fd_sc_hd__mux2_1 _09147_ (.A0(\core_pipeline.pipeline_registers.registers[26][12] ),
    .A1(\core_pipeline.pipeline_registers.registers[27][12] ),
    .S(net550),
    .X(_05190_));
 sky130_fd_sc_hd__a221o_1 _09148_ (.A1(\core_pipeline.pipeline_registers.registers[24][12] ),
    .A2(net424),
    .B1(net363),
    .B2(\core_pipeline.pipeline_registers.registers[25][12] ),
    .C1(net520),
    .X(_05191_));
 sky130_fd_sc_hd__a21o_1 _09149_ (.A1(net530),
    .A2(_05190_),
    .B1(_05191_),
    .X(_05192_));
 sky130_fd_sc_hd__mux2_1 _09150_ (.A0(\core_pipeline.pipeline_registers.registers[30][12] ),
    .A1(\core_pipeline.pipeline_registers.registers[31][12] ),
    .S(net550),
    .X(_05193_));
 sky130_fd_sc_hd__a221o_1 _09151_ (.A1(\core_pipeline.pipeline_registers.registers[28][12] ),
    .A2(net425),
    .B1(net364),
    .B2(\core_pipeline.pipeline_registers.registers[29][12] ),
    .C1(net463),
    .X(_05194_));
 sky130_fd_sc_hd__a21o_1 _09152_ (.A1(net530),
    .A2(_05193_),
    .B1(_05194_),
    .X(_05195_));
 sky130_fd_sc_hd__mux4_1 _09153_ (.A0(\core_pipeline.pipeline_registers.registers[16][12] ),
    .A1(\core_pipeline.pipeline_registers.registers[17][12] ),
    .A2(\core_pipeline.pipeline_registers.registers[18][12] ),
    .A3(\core_pipeline.pipeline_registers.registers[19][12] ),
    .S0(net550),
    .S1(net530),
    .X(_05196_));
 sky130_fd_sc_hd__mux4_1 _09154_ (.A0(\core_pipeline.pipeline_registers.registers[20][12] ),
    .A1(\core_pipeline.pipeline_registers.registers[21][12] ),
    .A2(\core_pipeline.pipeline_registers.registers[22][12] ),
    .A3(\core_pipeline.pipeline_registers.registers[23][12] ),
    .S0(net550),
    .S1(net530),
    .X(_05197_));
 sky130_fd_sc_hd__a22o_1 _09155_ (.A1(net429),
    .A2(_05196_),
    .B1(_05197_),
    .B2(net368),
    .X(_05198_));
 sky130_fd_sc_hd__a31o_1 _09156_ (.A1(net515),
    .A2(_05192_),
    .A3(_05195_),
    .B1(net461),
    .X(_05199_));
 sky130_fd_sc_hd__o211a_1 _09157_ (.A1(_05198_),
    .A2(_05199_),
    .B1(net144),
    .C1(_05189_),
    .X(_05200_));
 sky130_fd_sc_hd__a21o_1 _09158_ (.A1(\core_pipeline.decode_to_execute_rs2_data[12] ),
    .A2(net121),
    .B1(_05200_),
    .X(_00544_));
 sky130_fd_sc_hd__mux4_1 _09159_ (.A0(\core_pipeline.pipeline_registers.registers[12][13] ),
    .A1(\core_pipeline.pipeline_registers.registers[13][13] ),
    .A2(\core_pipeline.pipeline_registers.registers[14][13] ),
    .A3(\core_pipeline.pipeline_registers.registers[15][13] ),
    .S0(net552),
    .S1(net532),
    .X(_05201_));
 sky130_fd_sc_hd__mux4_1 _09160_ (.A0(\core_pipeline.pipeline_registers.registers[8][13] ),
    .A1(\core_pipeline.pipeline_registers.registers[9][13] ),
    .A2(\core_pipeline.pipeline_registers.registers[10][13] ),
    .A3(\core_pipeline.pipeline_registers.registers[11][13] ),
    .S0(net546),
    .S1(net526),
    .X(_05202_));
 sky130_fd_sc_hd__or2_1 _09161_ (.A(net519),
    .B(_05202_),
    .X(_05203_));
 sky130_fd_sc_hd__o211a_1 _09162_ (.A1(net463),
    .A2(_05201_),
    .B1(_05203_),
    .C1(net515),
    .X(_05204_));
 sky130_fd_sc_hd__mux4_1 _09163_ (.A0(\core_pipeline.pipeline_registers.registers[0][13] ),
    .A1(\core_pipeline.pipeline_registers.registers[1][13] ),
    .A2(\core_pipeline.pipeline_registers.registers[2][13] ),
    .A3(\core_pipeline.pipeline_registers.registers[3][13] ),
    .S0(net552),
    .S1(net533),
    .X(_05205_));
 sky130_fd_sc_hd__mux4_1 _09164_ (.A0(\core_pipeline.pipeline_registers.registers[4][13] ),
    .A1(\core_pipeline.pipeline_registers.registers[5][13] ),
    .A2(\core_pipeline.pipeline_registers.registers[6][13] ),
    .A3(\core_pipeline.pipeline_registers.registers[7][13] ),
    .S0(net552),
    .S1(net532),
    .X(_05206_));
 sky130_fd_sc_hd__a221o_1 _09165_ (.A1(net429),
    .A2(_05205_),
    .B1(_05206_),
    .B2(net368),
    .C1(\core_pipeline.decode_to_csr_read_address[4] ),
    .X(_05207_));
 sky130_fd_sc_hd__mux2_1 _09166_ (.A0(\core_pipeline.pipeline_registers.registers[30][13] ),
    .A1(\core_pipeline.pipeline_registers.registers[31][13] ),
    .S(net553),
    .X(_05208_));
 sky130_fd_sc_hd__a221o_1 _09167_ (.A1(\core_pipeline.pipeline_registers.registers[28][13] ),
    .A2(net425),
    .B1(net364),
    .B2(\core_pipeline.pipeline_registers.registers[29][13] ),
    .C1(net463),
    .X(_05209_));
 sky130_fd_sc_hd__a21o_1 _09168_ (.A1(net532),
    .A2(_05208_),
    .B1(_05209_),
    .X(_05210_));
 sky130_fd_sc_hd__mux2_1 _09169_ (.A0(\core_pipeline.pipeline_registers.registers[26][13] ),
    .A1(\core_pipeline.pipeline_registers.registers[27][13] ),
    .S(net553),
    .X(_05211_));
 sky130_fd_sc_hd__a221o_1 _09170_ (.A1(\core_pipeline.pipeline_registers.registers[24][13] ),
    .A2(net425),
    .B1(net364),
    .B2(\core_pipeline.pipeline_registers.registers[25][13] ),
    .C1(net521),
    .X(_05212_));
 sky130_fd_sc_hd__a21o_1 _09171_ (.A1(net533),
    .A2(_05211_),
    .B1(_05212_),
    .X(_05213_));
 sky130_fd_sc_hd__and3_1 _09172_ (.A(net515),
    .B(_05210_),
    .C(_05213_),
    .X(_05214_));
 sky130_fd_sc_hd__mux4_1 _09173_ (.A0(\core_pipeline.pipeline_registers.registers[20][13] ),
    .A1(\core_pipeline.pipeline_registers.registers[21][13] ),
    .A2(\core_pipeline.pipeline_registers.registers[22][13] ),
    .A3(\core_pipeline.pipeline_registers.registers[23][13] ),
    .S0(net552),
    .S1(net532),
    .X(_05215_));
 sky130_fd_sc_hd__mux2_1 _09174_ (.A0(\core_pipeline.pipeline_registers.registers[18][13] ),
    .A1(\core_pipeline.pipeline_registers.registers[19][13] ),
    .S(net552),
    .X(_05216_));
 sky130_fd_sc_hd__a31o_1 _09175_ (.A1(net532),
    .A2(net429),
    .A3(_05216_),
    .B1(net461),
    .X(_05217_));
 sky130_fd_sc_hd__a221o_1 _09176_ (.A1(\core_pipeline.pipeline_registers.registers[16][13] ),
    .A2(net279),
    .B1(net277),
    .B2(\core_pipeline.pipeline_registers.registers[17][13] ),
    .C1(_05217_),
    .X(_05218_));
 sky130_fd_sc_hd__a21o_1 _09177_ (.A1(net368),
    .A2(_05215_),
    .B1(_05218_),
    .X(_05219_));
 sky130_fd_sc_hd__o22a_2 _09178_ (.A1(_05204_),
    .A2(_05207_),
    .B1(_05214_),
    .B2(_05219_),
    .X(_05220_));
 sky130_fd_sc_hd__mux2_1 _09179_ (.A0(\core_pipeline.decode_to_execute_rs2_data[13] ),
    .A1(_05220_),
    .S(net139),
    .X(_00545_));
 sky130_fd_sc_hd__mux4_1 _09180_ (.A0(\core_pipeline.pipeline_registers.registers[8][14] ),
    .A1(\core_pipeline.pipeline_registers.registers[9][14] ),
    .A2(\core_pipeline.pipeline_registers.registers[10][14] ),
    .A3(\core_pipeline.pipeline_registers.registers[11][14] ),
    .S0(net552),
    .S1(net532),
    .X(_05221_));
 sky130_fd_sc_hd__or2_1 _09181_ (.A(net521),
    .B(_05221_),
    .X(_05222_));
 sky130_fd_sc_hd__mux4_1 _09182_ (.A0(\core_pipeline.pipeline_registers.registers[12][14] ),
    .A1(\core_pipeline.pipeline_registers.registers[13][14] ),
    .A2(\core_pipeline.pipeline_registers.registers[14][14] ),
    .A3(\core_pipeline.pipeline_registers.registers[15][14] ),
    .S0(net552),
    .S1(net533),
    .X(_05223_));
 sky130_fd_sc_hd__o211a_1 _09183_ (.A1(net463),
    .A2(_05223_),
    .B1(_05222_),
    .C1(net515),
    .X(_05224_));
 sky130_fd_sc_hd__mux4_2 _09184_ (.A0(\core_pipeline.pipeline_registers.registers[0][14] ),
    .A1(\core_pipeline.pipeline_registers.registers[1][14] ),
    .A2(\core_pipeline.pipeline_registers.registers[2][14] ),
    .A3(\core_pipeline.pipeline_registers.registers[3][14] ),
    .S0(net554),
    .S1(net533),
    .X(_05225_));
 sky130_fd_sc_hd__mux4_2 _09185_ (.A0(\core_pipeline.pipeline_registers.registers[4][14] ),
    .A1(\core_pipeline.pipeline_registers.registers[5][14] ),
    .A2(\core_pipeline.pipeline_registers.registers[6][14] ),
    .A3(\core_pipeline.pipeline_registers.registers[7][14] ),
    .S0(net554),
    .S1(net533),
    .X(_05226_));
 sky130_fd_sc_hd__a221o_4 _09186_ (.A1(net429),
    .A2(_05225_),
    .B1(_05226_),
    .B2(net368),
    .C1(_05224_),
    .X(_05227_));
 sky130_fd_sc_hd__mux2_1 _09187_ (.A0(\core_pipeline.pipeline_registers.registers[26][14] ),
    .A1(\core_pipeline.pipeline_registers.registers[27][14] ),
    .S(net547),
    .X(_05228_));
 sky130_fd_sc_hd__a221o_1 _09188_ (.A1(\core_pipeline.pipeline_registers.registers[24][14] ),
    .A2(net424),
    .B1(net363),
    .B2(\core_pipeline.pipeline_registers.registers[25][14] ),
    .C1(net519),
    .X(_05229_));
 sky130_fd_sc_hd__a21o_1 _09189_ (.A1(net527),
    .A2(_05228_),
    .B1(_05229_),
    .X(_05230_));
 sky130_fd_sc_hd__mux2_1 _09190_ (.A0(\core_pipeline.pipeline_registers.registers[30][14] ),
    .A1(\core_pipeline.pipeline_registers.registers[31][14] ),
    .S(net546),
    .X(_05231_));
 sky130_fd_sc_hd__a221o_1 _09191_ (.A1(\core_pipeline.pipeline_registers.registers[28][14] ),
    .A2(net424),
    .B1(net363),
    .B2(\core_pipeline.pipeline_registers.registers[29][14] ),
    .C1(net463),
    .X(_05232_));
 sky130_fd_sc_hd__a21o_1 _09192_ (.A1(net527),
    .A2(_05231_),
    .B1(_05232_),
    .X(_05233_));
 sky130_fd_sc_hd__mux4_1 _09193_ (.A0(\core_pipeline.pipeline_registers.registers[16][14] ),
    .A1(\core_pipeline.pipeline_registers.registers[17][14] ),
    .A2(\core_pipeline.pipeline_registers.registers[18][14] ),
    .A3(\core_pipeline.pipeline_registers.registers[19][14] ),
    .S0(net546),
    .S1(net526),
    .X(_05234_));
 sky130_fd_sc_hd__mux4_1 _09194_ (.A0(\core_pipeline.pipeline_registers.registers[20][14] ),
    .A1(\core_pipeline.pipeline_registers.registers[21][14] ),
    .A2(\core_pipeline.pipeline_registers.registers[22][14] ),
    .A3(\core_pipeline.pipeline_registers.registers[23][14] ),
    .S0(net546),
    .S1(net526),
    .X(_05235_));
 sky130_fd_sc_hd__a22o_1 _09195_ (.A1(net428),
    .A2(_05234_),
    .B1(_05235_),
    .B2(net367),
    .X(_05236_));
 sky130_fd_sc_hd__a31o_1 _09196_ (.A1(net514),
    .A2(_05230_),
    .A3(_05233_),
    .B1(net461),
    .X(_05237_));
 sky130_fd_sc_hd__o22a_2 _09197_ (.A1(net511),
    .A2(_05227_),
    .B1(_05236_),
    .B2(_05237_),
    .X(_05238_));
 sky130_fd_sc_hd__mux2_1 _09198_ (.A0(\core_pipeline.decode_to_execute_rs2_data[14] ),
    .A1(_05238_),
    .S(net139),
    .X(_00546_));
 sky130_fd_sc_hd__mux4_1 _09199_ (.A0(\core_pipeline.pipeline_registers.registers[12][15] ),
    .A1(\core_pipeline.pipeline_registers.registers[13][15] ),
    .A2(\core_pipeline.pipeline_registers.registers[14][15] ),
    .A3(\core_pipeline.pipeline_registers.registers[15][15] ),
    .S0(net553),
    .S1(net533),
    .X(_05239_));
 sky130_fd_sc_hd__mux4_1 _09200_ (.A0(\core_pipeline.pipeline_registers.registers[8][15] ),
    .A1(\core_pipeline.pipeline_registers.registers[9][15] ),
    .A2(\core_pipeline.pipeline_registers.registers[10][15] ),
    .A3(\core_pipeline.pipeline_registers.registers[11][15] ),
    .S0(net554),
    .S1(net533),
    .X(_05240_));
 sky130_fd_sc_hd__or2_1 _09201_ (.A(net521),
    .B(_05240_),
    .X(_05241_));
 sky130_fd_sc_hd__o211a_1 _09202_ (.A1(net463),
    .A2(_05239_),
    .B1(_05241_),
    .C1(net515),
    .X(_05242_));
 sky130_fd_sc_hd__mux4_1 _09203_ (.A0(\core_pipeline.pipeline_registers.registers[4][15] ),
    .A1(\core_pipeline.pipeline_registers.registers[5][15] ),
    .A2(\core_pipeline.pipeline_registers.registers[6][15] ),
    .A3(\core_pipeline.pipeline_registers.registers[7][15] ),
    .S0(net554),
    .S1(net533),
    .X(_05243_));
 sky130_fd_sc_hd__mux4_1 _09204_ (.A0(\core_pipeline.pipeline_registers.registers[0][15] ),
    .A1(\core_pipeline.pipeline_registers.registers[1][15] ),
    .A2(\core_pipeline.pipeline_registers.registers[2][15] ),
    .A3(\core_pipeline.pipeline_registers.registers[3][15] ),
    .S0(net553),
    .S1(net533),
    .X(_05244_));
 sky130_fd_sc_hd__a221o_1 _09205_ (.A1(net368),
    .A2(_05243_),
    .B1(_05244_),
    .B2(net429),
    .C1(\core_pipeline.decode_to_csr_read_address[4] ),
    .X(_05245_));
 sky130_fd_sc_hd__mux2_1 _09206_ (.A0(\core_pipeline.pipeline_registers.registers[30][15] ),
    .A1(\core_pipeline.pipeline_registers.registers[31][15] ),
    .S(net550),
    .X(_05246_));
 sky130_fd_sc_hd__a221o_1 _09207_ (.A1(\core_pipeline.pipeline_registers.registers[28][15] ),
    .A2(net425),
    .B1(net364),
    .B2(\core_pipeline.pipeline_registers.registers[29][15] ),
    .C1(net463),
    .X(_05247_));
 sky130_fd_sc_hd__a21o_1 _09208_ (.A1(net543),
    .A2(_05246_),
    .B1(_05247_),
    .X(_05248_));
 sky130_fd_sc_hd__mux2_1 _09209_ (.A0(\core_pipeline.pipeline_registers.registers[26][15] ),
    .A1(\core_pipeline.pipeline_registers.registers[27][15] ),
    .S(net550),
    .X(_05249_));
 sky130_fd_sc_hd__a221o_1 _09210_ (.A1(\core_pipeline.pipeline_registers.registers[24][15] ),
    .A2(net425),
    .B1(net364),
    .B2(\core_pipeline.pipeline_registers.registers[25][15] ),
    .C1(net519),
    .X(_05250_));
 sky130_fd_sc_hd__a21o_1 _09211_ (.A1(net530),
    .A2(_05249_),
    .B1(_05250_),
    .X(_05251_));
 sky130_fd_sc_hd__and3_1 _09212_ (.A(net515),
    .B(_05248_),
    .C(_05251_),
    .X(_05252_));
 sky130_fd_sc_hd__mux4_1 _09213_ (.A0(\core_pipeline.pipeline_registers.registers[20][15] ),
    .A1(\core_pipeline.pipeline_registers.registers[21][15] ),
    .A2(\core_pipeline.pipeline_registers.registers[22][15] ),
    .A3(\core_pipeline.pipeline_registers.registers[23][15] ),
    .S0(net553),
    .S1(net532),
    .X(_05253_));
 sky130_fd_sc_hd__a31o_1 _09214_ (.A1(\core_pipeline.pipeline_registers.registers[16][15] ),
    .A2(net428),
    .A3(net425),
    .B1(net461),
    .X(_05254_));
 sky130_fd_sc_hd__mux2_1 _09215_ (.A0(\core_pipeline.pipeline_registers.registers[18][15] ),
    .A1(\core_pipeline.pipeline_registers.registers[19][15] ),
    .S(net553),
    .X(_05255_));
 sky130_fd_sc_hd__a22o_1 _09216_ (.A1(\core_pipeline.pipeline_registers.registers[17][15] ),
    .A2(net277),
    .B1(net361),
    .B2(_05255_),
    .X(_05256_));
 sky130_fd_sc_hd__a211o_1 _09217_ (.A1(net367),
    .A2(_05253_),
    .B1(_05254_),
    .C1(_05256_),
    .X(_05257_));
 sky130_fd_sc_hd__o22a_1 _09218_ (.A1(_05242_),
    .A2(_05245_),
    .B1(_05252_),
    .B2(_05257_),
    .X(_05258_));
 sky130_fd_sc_hd__mux2_1 _09219_ (.A0(\core_pipeline.decode_to_execute_rs2_data[15] ),
    .A1(_05258_),
    .S(net140),
    .X(_00547_));
 sky130_fd_sc_hd__mux4_1 _09220_ (.A0(\core_pipeline.pipeline_registers.registers[8][16] ),
    .A1(\core_pipeline.pipeline_registers.registers[9][16] ),
    .A2(\core_pipeline.pipeline_registers.registers[10][16] ),
    .A3(\core_pipeline.pipeline_registers.registers[11][16] ),
    .S0(net545),
    .S1(net525),
    .X(_05259_));
 sky130_fd_sc_hd__or2_1 _09221_ (.A(net519),
    .B(_05259_),
    .X(_05260_));
 sky130_fd_sc_hd__mux4_1 _09222_ (.A0(\core_pipeline.pipeline_registers.registers[12][16] ),
    .A1(\core_pipeline.pipeline_registers.registers[13][16] ),
    .A2(\core_pipeline.pipeline_registers.registers[14][16] ),
    .A3(\core_pipeline.pipeline_registers.registers[15][16] ),
    .S0(net544),
    .S1(net525),
    .X(_05261_));
 sky130_fd_sc_hd__o211a_1 _09223_ (.A1(net462),
    .A2(_05261_),
    .B1(_05260_),
    .C1(net514),
    .X(_05262_));
 sky130_fd_sc_hd__mux4_1 _09224_ (.A0(\core_pipeline.pipeline_registers.registers[0][16] ),
    .A1(\core_pipeline.pipeline_registers.registers[1][16] ),
    .A2(\core_pipeline.pipeline_registers.registers[2][16] ),
    .A3(\core_pipeline.pipeline_registers.registers[3][16] ),
    .S0(net544),
    .S1(net525),
    .X(_05263_));
 sky130_fd_sc_hd__mux4_1 _09225_ (.A0(\core_pipeline.pipeline_registers.registers[4][16] ),
    .A1(\core_pipeline.pipeline_registers.registers[5][16] ),
    .A2(\core_pipeline.pipeline_registers.registers[6][16] ),
    .A3(\core_pipeline.pipeline_registers.registers[7][16] ),
    .S0(net544),
    .S1(net525),
    .X(_05264_));
 sky130_fd_sc_hd__a221o_1 _09226_ (.A1(net428),
    .A2(_05263_),
    .B1(_05264_),
    .B2(net367),
    .C1(_05262_),
    .X(_05265_));
 sky130_fd_sc_hd__mux2_1 _09227_ (.A0(\core_pipeline.pipeline_registers.registers[26][16] ),
    .A1(\core_pipeline.pipeline_registers.registers[27][16] ),
    .S(net548),
    .X(_05266_));
 sky130_fd_sc_hd__a221o_1 _09228_ (.A1(\core_pipeline.pipeline_registers.registers[24][16] ),
    .A2(net424),
    .B1(net363),
    .B2(\core_pipeline.pipeline_registers.registers[25][16] ),
    .C1(net520),
    .X(_05267_));
 sky130_fd_sc_hd__a21o_1 _09229_ (.A1(net529),
    .A2(_05266_),
    .B1(_05267_),
    .X(_05268_));
 sky130_fd_sc_hd__mux2_1 _09230_ (.A0(\core_pipeline.pipeline_registers.registers[30][16] ),
    .A1(\core_pipeline.pipeline_registers.registers[31][16] ),
    .S(net548),
    .X(_05269_));
 sky130_fd_sc_hd__a221o_1 _09231_ (.A1(\core_pipeline.pipeline_registers.registers[28][16] ),
    .A2(net424),
    .B1(net363),
    .B2(\core_pipeline.pipeline_registers.registers[29][16] ),
    .C1(net462),
    .X(_05270_));
 sky130_fd_sc_hd__a21o_1 _09232_ (.A1(net529),
    .A2(_05269_),
    .B1(_05270_),
    .X(_05271_));
 sky130_fd_sc_hd__mux4_1 _09233_ (.A0(\core_pipeline.pipeline_registers.registers[16][16] ),
    .A1(\core_pipeline.pipeline_registers.registers[17][16] ),
    .A2(\core_pipeline.pipeline_registers.registers[18][16] ),
    .A3(\core_pipeline.pipeline_registers.registers[19][16] ),
    .S0(net548),
    .S1(net529),
    .X(_05272_));
 sky130_fd_sc_hd__mux4_1 _09234_ (.A0(\core_pipeline.pipeline_registers.registers[20][16] ),
    .A1(\core_pipeline.pipeline_registers.registers[21][16] ),
    .A2(\core_pipeline.pipeline_registers.registers[22][16] ),
    .A3(\core_pipeline.pipeline_registers.registers[23][16] ),
    .S0(net548),
    .S1(net529),
    .X(_05273_));
 sky130_fd_sc_hd__a22o_1 _09235_ (.A1(net429),
    .A2(_05272_),
    .B1(_05273_),
    .B2(net368),
    .X(_05274_));
 sky130_fd_sc_hd__a31o_1 _09236_ (.A1(net515),
    .A2(_05268_),
    .A3(_05271_),
    .B1(net461),
    .X(_05275_));
 sky130_fd_sc_hd__o22a_1 _09237_ (.A1(net511),
    .A2(_05265_),
    .B1(_05274_),
    .B2(_05275_),
    .X(_05276_));
 sky130_fd_sc_hd__mux2_1 _09238_ (.A0(\core_pipeline.decode_to_execute_rs2_data[16] ),
    .A1(_05276_),
    .S(net144),
    .X(_00548_));
 sky130_fd_sc_hd__mux4_1 _09239_ (.A0(\core_pipeline.pipeline_registers.registers[12][17] ),
    .A1(\core_pipeline.pipeline_registers.registers[13][17] ),
    .A2(\core_pipeline.pipeline_registers.registers[14][17] ),
    .A3(\core_pipeline.pipeline_registers.registers[15][17] ),
    .S0(net557),
    .S1(net535),
    .X(_05277_));
 sky130_fd_sc_hd__mux4_1 _09240_ (.A0(\core_pipeline.pipeline_registers.registers[8][17] ),
    .A1(\core_pipeline.pipeline_registers.registers[9][17] ),
    .A2(\core_pipeline.pipeline_registers.registers[10][17] ),
    .A3(\core_pipeline.pipeline_registers.registers[11][17] ),
    .S0(net557),
    .S1(net535),
    .X(_05278_));
 sky130_fd_sc_hd__or2_1 _09241_ (.A(net523),
    .B(_05278_),
    .X(_05279_));
 sky130_fd_sc_hd__o211a_1 _09242_ (.A1(net464),
    .A2(_05277_),
    .B1(_05279_),
    .C1(net516),
    .X(_05280_));
 sky130_fd_sc_hd__mux4_1 _09243_ (.A0(\core_pipeline.pipeline_registers.registers[4][17] ),
    .A1(\core_pipeline.pipeline_registers.registers[5][17] ),
    .A2(\core_pipeline.pipeline_registers.registers[6][17] ),
    .A3(\core_pipeline.pipeline_registers.registers[7][17] ),
    .S0(net561),
    .S1(net538),
    .X(_05281_));
 sky130_fd_sc_hd__mux4_1 _09244_ (.A0(\core_pipeline.pipeline_registers.registers[0][17] ),
    .A1(\core_pipeline.pipeline_registers.registers[1][17] ),
    .A2(\core_pipeline.pipeline_registers.registers[2][17] ),
    .A3(\core_pipeline.pipeline_registers.registers[3][17] ),
    .S0(net561),
    .S1(net538),
    .X(_05282_));
 sky130_fd_sc_hd__a221o_1 _09245_ (.A1(net369),
    .A2(_05281_),
    .B1(_05282_),
    .B2(net430),
    .C1(net512),
    .X(_05283_));
 sky130_fd_sc_hd__mux2_1 _09246_ (.A0(\core_pipeline.pipeline_registers.registers[30][17] ),
    .A1(\core_pipeline.pipeline_registers.registers[31][17] ),
    .S(net561),
    .X(_05284_));
 sky130_fd_sc_hd__a221o_1 _09247_ (.A1(\core_pipeline.pipeline_registers.registers[28][17] ),
    .A2(net426),
    .B1(net366),
    .B2(\core_pipeline.pipeline_registers.registers[29][17] ),
    .C1(net464),
    .X(_05285_));
 sky130_fd_sc_hd__a21o_1 _09248_ (.A1(net538),
    .A2(_05284_),
    .B1(_05285_),
    .X(_05286_));
 sky130_fd_sc_hd__mux2_1 _09249_ (.A0(\core_pipeline.pipeline_registers.registers[26][17] ),
    .A1(\core_pipeline.pipeline_registers.registers[27][17] ),
    .S(net559),
    .X(_05287_));
 sky130_fd_sc_hd__a221o_1 _09250_ (.A1(\core_pipeline.pipeline_registers.registers[24][17] ),
    .A2(net426),
    .B1(net365),
    .B2(\core_pipeline.pipeline_registers.registers[25][17] ),
    .C1(net522),
    .X(_05288_));
 sky130_fd_sc_hd__a21o_1 _09251_ (.A1(net538),
    .A2(_05287_),
    .B1(_05288_),
    .X(_05289_));
 sky130_fd_sc_hd__and3_1 _09252_ (.A(net516),
    .B(_05286_),
    .C(_05289_),
    .X(_05290_));
 sky130_fd_sc_hd__mux4_1 _09253_ (.A0(\core_pipeline.pipeline_registers.registers[20][17] ),
    .A1(\core_pipeline.pipeline_registers.registers[21][17] ),
    .A2(\core_pipeline.pipeline_registers.registers[22][17] ),
    .A3(\core_pipeline.pipeline_registers.registers[23][17] ),
    .S0(net561),
    .S1(net538),
    .X(_05291_));
 sky130_fd_sc_hd__mux2_1 _09254_ (.A0(\core_pipeline.pipeline_registers.registers[18][17] ),
    .A1(\core_pipeline.pipeline_registers.registers[19][17] ),
    .S(net558),
    .X(_05292_));
 sky130_fd_sc_hd__a31o_1 _09255_ (.A1(net536),
    .A2(net430),
    .A3(_05292_),
    .B1(net460),
    .X(_05293_));
 sky130_fd_sc_hd__a221o_1 _09256_ (.A1(\core_pipeline.pipeline_registers.registers[16][17] ),
    .A2(net278),
    .B1(net276),
    .B2(\core_pipeline.pipeline_registers.registers[17][17] ),
    .C1(_05293_),
    .X(_05294_));
 sky130_fd_sc_hd__a21o_1 _09257_ (.A1(net369),
    .A2(_05291_),
    .B1(_05294_),
    .X(_05295_));
 sky130_fd_sc_hd__o22a_1 _09258_ (.A1(_05280_),
    .A2(_05283_),
    .B1(_05290_),
    .B2(_05295_),
    .X(_05296_));
 sky130_fd_sc_hd__mux2_1 _09259_ (.A0(\core_pipeline.decode_to_execute_rs2_data[17] ),
    .A1(_05296_),
    .S(net145),
    .X(_00549_));
 sky130_fd_sc_hd__mux4_1 _09260_ (.A0(\core_pipeline.pipeline_registers.registers[8][18] ),
    .A1(\core_pipeline.pipeline_registers.registers[9][18] ),
    .A2(\core_pipeline.pipeline_registers.registers[10][18] ),
    .A3(\core_pipeline.pipeline_registers.registers[11][18] ),
    .S0(net560),
    .S1(net537),
    .X(_05297_));
 sky130_fd_sc_hd__or2_1 _09261_ (.A(net523),
    .B(_05297_),
    .X(_05298_));
 sky130_fd_sc_hd__mux4_1 _09262_ (.A0(\core_pipeline.pipeline_registers.registers[12][18] ),
    .A1(\core_pipeline.pipeline_registers.registers[13][18] ),
    .A2(\core_pipeline.pipeline_registers.registers[14][18] ),
    .A3(\core_pipeline.pipeline_registers.registers[15][18] ),
    .S0(net559),
    .S1(net538),
    .X(_05299_));
 sky130_fd_sc_hd__o211a_1 _09263_ (.A1(net464),
    .A2(_05299_),
    .B1(_05298_),
    .C1(net516),
    .X(_05300_));
 sky130_fd_sc_hd__mux4_1 _09264_ (.A0(\core_pipeline.pipeline_registers.registers[4][18] ),
    .A1(\core_pipeline.pipeline_registers.registers[5][18] ),
    .A2(\core_pipeline.pipeline_registers.registers[6][18] ),
    .A3(\core_pipeline.pipeline_registers.registers[7][18] ),
    .S0(net561),
    .S1(net538),
    .X(_05301_));
 sky130_fd_sc_hd__mux2_1 _09265_ (.A0(\core_pipeline.pipeline_registers.registers[2][18] ),
    .A1(\core_pipeline.pipeline_registers.registers[3][18] ),
    .S(net561),
    .X(_05302_));
 sky130_fd_sc_hd__a22o_1 _09266_ (.A1(\core_pipeline.pipeline_registers.registers[1][18] ),
    .A2(net276),
    .B1(net361),
    .B2(_05302_),
    .X(_05303_));
 sky130_fd_sc_hd__a211o_1 _09267_ (.A1(\core_pipeline.pipeline_registers.registers[0][18] ),
    .A2(net278),
    .B1(_05303_),
    .C1(net512),
    .X(_05304_));
 sky130_fd_sc_hd__a211o_1 _09268_ (.A1(net369),
    .A2(_05301_),
    .B1(_05304_),
    .C1(_05300_),
    .X(_05305_));
 sky130_fd_sc_hd__mux2_1 _09269_ (.A0(\core_pipeline.pipeline_registers.registers[30][18] ),
    .A1(\core_pipeline.pipeline_registers.registers[31][18] ),
    .S(net561),
    .X(_05306_));
 sky130_fd_sc_hd__a221o_1 _09270_ (.A1(\core_pipeline.pipeline_registers.registers[28][18] ),
    .A2(net426),
    .B1(net366),
    .B2(\core_pipeline.pipeline_registers.registers[29][18] ),
    .C1(net464),
    .X(_05307_));
 sky130_fd_sc_hd__a21o_1 _09271_ (.A1(net538),
    .A2(_05306_),
    .B1(_05307_),
    .X(_05308_));
 sky130_fd_sc_hd__mux2_1 _09272_ (.A0(\core_pipeline.pipeline_registers.registers[26][18] ),
    .A1(\core_pipeline.pipeline_registers.registers[27][18] ),
    .S(net561),
    .X(_05309_));
 sky130_fd_sc_hd__a221o_1 _09273_ (.A1(\core_pipeline.pipeline_registers.registers[24][18] ),
    .A2(net426),
    .B1(net366),
    .B2(\core_pipeline.pipeline_registers.registers[25][18] ),
    .C1(net523),
    .X(_05310_));
 sky130_fd_sc_hd__a21o_1 _09274_ (.A1(net538),
    .A2(_05309_),
    .B1(_05310_),
    .X(_05311_));
 sky130_fd_sc_hd__and3_1 _09275_ (.A(net518),
    .B(_05308_),
    .C(_05311_),
    .X(_05312_));
 sky130_fd_sc_hd__mux4_1 _09276_ (.A0(\core_pipeline.pipeline_registers.registers[20][18] ),
    .A1(\core_pipeline.pipeline_registers.registers[21][18] ),
    .A2(\core_pipeline.pipeline_registers.registers[22][18] ),
    .A3(\core_pipeline.pipeline_registers.registers[23][18] ),
    .S0(net561),
    .S1(net538),
    .X(_05313_));
 sky130_fd_sc_hd__mux2_1 _09277_ (.A0(\core_pipeline.pipeline_registers.registers[18][18] ),
    .A1(\core_pipeline.pipeline_registers.registers[19][18] ),
    .S(net561),
    .X(_05314_));
 sky130_fd_sc_hd__a22o_1 _09278_ (.A1(\core_pipeline.pipeline_registers.registers[16][18] ),
    .A2(net278),
    .B1(net362),
    .B2(_05314_),
    .X(_05315_));
 sky130_fd_sc_hd__a211o_1 _09279_ (.A1(\core_pipeline.pipeline_registers.registers[17][18] ),
    .A2(net276),
    .B1(_05315_),
    .C1(net460),
    .X(_05316_));
 sky130_fd_sc_hd__a211o_1 _09280_ (.A1(net369),
    .A2(_05313_),
    .B1(_05316_),
    .C1(_05312_),
    .X(_05317_));
 sky130_fd_sc_hd__and3_1 _09281_ (.A(net145),
    .B(_05305_),
    .C(_05317_),
    .X(_05318_));
 sky130_fd_sc_hd__a21o_1 _09282_ (.A1(\core_pipeline.decode_to_execute_rs2_data[18] ),
    .A2(net135),
    .B1(_05318_),
    .X(_00550_));
 sky130_fd_sc_hd__mux4_1 _09283_ (.A0(\core_pipeline.pipeline_registers.registers[8][19] ),
    .A1(\core_pipeline.pipeline_registers.registers[9][19] ),
    .A2(\core_pipeline.pipeline_registers.registers[10][19] ),
    .A3(\core_pipeline.pipeline_registers.registers[11][19] ),
    .S0(net559),
    .S1(net537),
    .X(_05319_));
 sky130_fd_sc_hd__or2_1 _09284_ (.A(net523),
    .B(_05319_),
    .X(_05320_));
 sky130_fd_sc_hd__mux4_1 _09285_ (.A0(\core_pipeline.pipeline_registers.registers[12][19] ),
    .A1(\core_pipeline.pipeline_registers.registers[13][19] ),
    .A2(\core_pipeline.pipeline_registers.registers[14][19] ),
    .A3(\core_pipeline.pipeline_registers.registers[15][19] ),
    .S0(net559),
    .S1(net537),
    .X(_05321_));
 sky130_fd_sc_hd__o211a_1 _09286_ (.A1(net465),
    .A2(_05321_),
    .B1(_05320_),
    .C1(net518),
    .X(_05322_));
 sky130_fd_sc_hd__mux4_1 _09287_ (.A0(\core_pipeline.pipeline_registers.registers[4][19] ),
    .A1(\core_pipeline.pipeline_registers.registers[5][19] ),
    .A2(\core_pipeline.pipeline_registers.registers[6][19] ),
    .A3(\core_pipeline.pipeline_registers.registers[7][19] ),
    .S0(net559),
    .S1(net537),
    .X(_05323_));
 sky130_fd_sc_hd__mux2_1 _09288_ (.A0(\core_pipeline.pipeline_registers.registers[2][19] ),
    .A1(\core_pipeline.pipeline_registers.registers[3][19] ),
    .S(net559),
    .X(_05324_));
 sky130_fd_sc_hd__a22o_1 _09289_ (.A1(\core_pipeline.pipeline_registers.registers[1][19] ),
    .A2(net276),
    .B1(net361),
    .B2(_05324_),
    .X(_05325_));
 sky130_fd_sc_hd__a211o_1 _09290_ (.A1(\core_pipeline.pipeline_registers.registers[0][19] ),
    .A2(net278),
    .B1(_05325_),
    .C1(net512),
    .X(_05326_));
 sky130_fd_sc_hd__a211o_1 _09291_ (.A1(net369),
    .A2(_05323_),
    .B1(_05326_),
    .C1(_05322_),
    .X(_05327_));
 sky130_fd_sc_hd__mux2_1 _09292_ (.A0(\core_pipeline.pipeline_registers.registers[26][19] ),
    .A1(\core_pipeline.pipeline_registers.registers[27][19] ),
    .S(net559),
    .X(_05328_));
 sky130_fd_sc_hd__a221o_1 _09293_ (.A1(\core_pipeline.pipeline_registers.registers[24][19] ),
    .A2(net426),
    .B1(net366),
    .B2(\core_pipeline.pipeline_registers.registers[25][19] ),
    .C1(net522),
    .X(_05329_));
 sky130_fd_sc_hd__a21o_1 _09294_ (.A1(net537),
    .A2(_05328_),
    .B1(_05329_),
    .X(_05330_));
 sky130_fd_sc_hd__mux2_1 _09295_ (.A0(\core_pipeline.pipeline_registers.registers[30][19] ),
    .A1(\core_pipeline.pipeline_registers.registers[31][19] ),
    .S(net559),
    .X(_05331_));
 sky130_fd_sc_hd__a221o_1 _09296_ (.A1(\core_pipeline.pipeline_registers.registers[28][19] ),
    .A2(net426),
    .B1(net366),
    .B2(\core_pipeline.pipeline_registers.registers[29][19] ),
    .C1(net465),
    .X(_05332_));
 sky130_fd_sc_hd__a21o_1 _09297_ (.A1(net537),
    .A2(_05331_),
    .B1(_05332_),
    .X(_05333_));
 sky130_fd_sc_hd__mux4_1 _09298_ (.A0(\core_pipeline.pipeline_registers.registers[16][19] ),
    .A1(\core_pipeline.pipeline_registers.registers[17][19] ),
    .A2(\core_pipeline.pipeline_registers.registers[18][19] ),
    .A3(\core_pipeline.pipeline_registers.registers[19][19] ),
    .S0(net559),
    .S1(net537),
    .X(_05334_));
 sky130_fd_sc_hd__mux4_1 _09299_ (.A0(\core_pipeline.pipeline_registers.registers[20][19] ),
    .A1(\core_pipeline.pipeline_registers.registers[21][19] ),
    .A2(\core_pipeline.pipeline_registers.registers[22][19] ),
    .A3(\core_pipeline.pipeline_registers.registers[23][19] ),
    .S0(net559),
    .S1(net537),
    .X(_05335_));
 sky130_fd_sc_hd__a22o_1 _09300_ (.A1(net430),
    .A2(_05334_),
    .B1(_05335_),
    .B2(net369),
    .X(_05336_));
 sky130_fd_sc_hd__a31o_1 _09301_ (.A1(net516),
    .A2(_05330_),
    .A3(_05333_),
    .B1(net460),
    .X(_05337_));
 sky130_fd_sc_hd__o211a_2 _09302_ (.A1(_05336_),
    .A2(_05337_),
    .B1(net145),
    .C1(_05327_),
    .X(_05338_));
 sky130_fd_sc_hd__a21o_1 _09303_ (.A1(\core_pipeline.decode_to_execute_rs2_data[19] ),
    .A2(net135),
    .B1(_05338_),
    .X(_00551_));
 sky130_fd_sc_hd__mux4_1 _09304_ (.A0(\core_pipeline.pipeline_registers.registers[12][20] ),
    .A1(\core_pipeline.pipeline_registers.registers[13][20] ),
    .A2(\core_pipeline.pipeline_registers.registers[14][20] ),
    .A3(\core_pipeline.pipeline_registers.registers[15][20] ),
    .S0(net560),
    .S1(net539),
    .X(_05339_));
 sky130_fd_sc_hd__mux4_1 _09305_ (.A0(\core_pipeline.pipeline_registers.registers[8][20] ),
    .A1(\core_pipeline.pipeline_registers.registers[9][20] ),
    .A2(\core_pipeline.pipeline_registers.registers[10][20] ),
    .A3(\core_pipeline.pipeline_registers.registers[11][20] ),
    .S0(net560),
    .S1(net537),
    .X(_05340_));
 sky130_fd_sc_hd__or2_1 _09306_ (.A(net523),
    .B(_05340_),
    .X(_05341_));
 sky130_fd_sc_hd__o211a_1 _09307_ (.A1(net464),
    .A2(_05339_),
    .B1(_05341_),
    .C1(net518),
    .X(_05342_));
 sky130_fd_sc_hd__mux4_1 _09308_ (.A0(\core_pipeline.pipeline_registers.registers[4][20] ),
    .A1(\core_pipeline.pipeline_registers.registers[5][20] ),
    .A2(\core_pipeline.pipeline_registers.registers[6][20] ),
    .A3(\core_pipeline.pipeline_registers.registers[7][20] ),
    .S0(net560),
    .S1(net539),
    .X(_05343_));
 sky130_fd_sc_hd__mux4_1 _09309_ (.A0(\core_pipeline.pipeline_registers.registers[0][20] ),
    .A1(\core_pipeline.pipeline_registers.registers[1][20] ),
    .A2(\core_pipeline.pipeline_registers.registers[2][20] ),
    .A3(\core_pipeline.pipeline_registers.registers[3][20] ),
    .S0(net560),
    .S1(net539),
    .X(_05344_));
 sky130_fd_sc_hd__a221o_1 _09310_ (.A1(net369),
    .A2(_05343_),
    .B1(_05344_),
    .B2(net430),
    .C1(net512),
    .X(_05345_));
 sky130_fd_sc_hd__mux2_1 _09311_ (.A0(\core_pipeline.pipeline_registers.registers[30][20] ),
    .A1(\core_pipeline.pipeline_registers.registers[31][20] ),
    .S(net560),
    .X(_05346_));
 sky130_fd_sc_hd__a221o_1 _09312_ (.A1(\core_pipeline.pipeline_registers.registers[28][20] ),
    .A2(net426),
    .B1(net365),
    .B2(\core_pipeline.pipeline_registers.registers[29][20] ),
    .C1(net464),
    .X(_05347_));
 sky130_fd_sc_hd__a21o_1 _09313_ (.A1(net537),
    .A2(_05346_),
    .B1(_05347_),
    .X(_05348_));
 sky130_fd_sc_hd__mux2_1 _09314_ (.A0(\core_pipeline.pipeline_registers.registers[26][20] ),
    .A1(\core_pipeline.pipeline_registers.registers[27][20] ),
    .S(net560),
    .X(_05349_));
 sky130_fd_sc_hd__a221o_1 _09315_ (.A1(\core_pipeline.pipeline_registers.registers[24][20] ),
    .A2(net427),
    .B1(net365),
    .B2(\core_pipeline.pipeline_registers.registers[25][20] ),
    .C1(net523),
    .X(_05350_));
 sky130_fd_sc_hd__a21o_1 _09316_ (.A1(net537),
    .A2(_05349_),
    .B1(_05350_),
    .X(_05351_));
 sky130_fd_sc_hd__and3_1 _09317_ (.A(net518),
    .B(_05348_),
    .C(_05351_),
    .X(_05352_));
 sky130_fd_sc_hd__mux4_1 _09318_ (.A0(\core_pipeline.pipeline_registers.registers[20][20] ),
    .A1(\core_pipeline.pipeline_registers.registers[21][20] ),
    .A2(\core_pipeline.pipeline_registers.registers[22][20] ),
    .A3(\core_pipeline.pipeline_registers.registers[23][20] ),
    .S0(net560),
    .S1(net537),
    .X(_05353_));
 sky130_fd_sc_hd__a31o_1 _09319_ (.A1(\core_pipeline.pipeline_registers.registers[17][20] ),
    .A2(net430),
    .A3(net365),
    .B1(net460),
    .X(_05354_));
 sky130_fd_sc_hd__mux2_1 _09320_ (.A0(\core_pipeline.pipeline_registers.registers[18][20] ),
    .A1(\core_pipeline.pipeline_registers.registers[19][20] ),
    .S(net560),
    .X(_05355_));
 sky130_fd_sc_hd__a22o_1 _09321_ (.A1(\core_pipeline.pipeline_registers.registers[16][20] ),
    .A2(net278),
    .B1(net362),
    .B2(_05355_),
    .X(_05356_));
 sky130_fd_sc_hd__a211o_1 _09322_ (.A1(net369),
    .A2(_05353_),
    .B1(_05354_),
    .C1(_05356_),
    .X(_05357_));
 sky130_fd_sc_hd__o22a_1 _09323_ (.A1(_05342_),
    .A2(_05345_),
    .B1(_05352_),
    .B2(_05357_),
    .X(_05358_));
 sky130_fd_sc_hd__mux2_1 _09324_ (.A0(\core_pipeline.decode_to_execute_rs2_data[20] ),
    .A1(_05358_),
    .S(net145),
    .X(_00552_));
 sky130_fd_sc_hd__mux4_1 _09325_ (.A0(\core_pipeline.pipeline_registers.registers[8][21] ),
    .A1(\core_pipeline.pipeline_registers.registers[9][21] ),
    .A2(\core_pipeline.pipeline_registers.registers[10][21] ),
    .A3(\core_pipeline.pipeline_registers.registers[11][21] ),
    .S0(net564),
    .S1(net541),
    .X(_05359_));
 sky130_fd_sc_hd__or2_1 _09326_ (.A(net524),
    .B(_05359_),
    .X(_05360_));
 sky130_fd_sc_hd__mux4_1 _09327_ (.A0(\core_pipeline.pipeline_registers.registers[12][21] ),
    .A1(\core_pipeline.pipeline_registers.registers[13][21] ),
    .A2(\core_pipeline.pipeline_registers.registers[14][21] ),
    .A3(\core_pipeline.pipeline_registers.registers[15][21] ),
    .S0(net563),
    .S1(net540),
    .X(_05361_));
 sky130_fd_sc_hd__o211a_1 _09328_ (.A1(net465),
    .A2(_05361_),
    .B1(_05360_),
    .C1(net517),
    .X(_05362_));
 sky130_fd_sc_hd__mux4_1 _09329_ (.A0(\core_pipeline.pipeline_registers.registers[4][21] ),
    .A1(\core_pipeline.pipeline_registers.registers[5][21] ),
    .A2(\core_pipeline.pipeline_registers.registers[6][21] ),
    .A3(\core_pipeline.pipeline_registers.registers[7][21] ),
    .S0(net563),
    .S1(net540),
    .X(_05363_));
 sky130_fd_sc_hd__mux2_1 _09330_ (.A0(\core_pipeline.pipeline_registers.registers[2][21] ),
    .A1(\core_pipeline.pipeline_registers.registers[3][21] ),
    .S(net563),
    .X(_05364_));
 sky130_fd_sc_hd__a22o_1 _09331_ (.A1(\core_pipeline.pipeline_registers.registers[1][21] ),
    .A2(net276),
    .B1(net362),
    .B2(_05364_),
    .X(_05365_));
 sky130_fd_sc_hd__a211o_1 _09332_ (.A1(\core_pipeline.pipeline_registers.registers[0][21] ),
    .A2(net279),
    .B1(_05365_),
    .C1(net513),
    .X(_05366_));
 sky130_fd_sc_hd__a211o_1 _09333_ (.A1(net369),
    .A2(_05363_),
    .B1(_05366_),
    .C1(_05362_),
    .X(_05367_));
 sky130_fd_sc_hd__mux2_1 _09334_ (.A0(\core_pipeline.pipeline_registers.registers[30][21] ),
    .A1(\core_pipeline.pipeline_registers.registers[31][21] ),
    .S(net564),
    .X(_05368_));
 sky130_fd_sc_hd__a221o_1 _09335_ (.A1(\core_pipeline.pipeline_registers.registers[28][21] ),
    .A2(net427),
    .B1(net366),
    .B2(\core_pipeline.pipeline_registers.registers[29][21] ),
    .C1(net465),
    .X(_05369_));
 sky130_fd_sc_hd__a21o_1 _09336_ (.A1(net541),
    .A2(_05368_),
    .B1(_05369_),
    .X(_05370_));
 sky130_fd_sc_hd__mux2_1 _09337_ (.A0(\core_pipeline.pipeline_registers.registers[26][21] ),
    .A1(\core_pipeline.pipeline_registers.registers[27][21] ),
    .S(net564),
    .X(_05371_));
 sky130_fd_sc_hd__a221o_1 _09338_ (.A1(\core_pipeline.pipeline_registers.registers[24][21] ),
    .A2(net427),
    .B1(net366),
    .B2(\core_pipeline.pipeline_registers.registers[25][21] ),
    .C1(net524),
    .X(_05372_));
 sky130_fd_sc_hd__a21o_1 _09339_ (.A1(net540),
    .A2(_05371_),
    .B1(_05372_),
    .X(_05373_));
 sky130_fd_sc_hd__and3_1 _09340_ (.A(net517),
    .B(_05370_),
    .C(_05373_),
    .X(_05374_));
 sky130_fd_sc_hd__mux4_1 _09341_ (.A0(\core_pipeline.pipeline_registers.registers[20][21] ),
    .A1(\core_pipeline.pipeline_registers.registers[21][21] ),
    .A2(\core_pipeline.pipeline_registers.registers[22][21] ),
    .A3(\core_pipeline.pipeline_registers.registers[23][21] ),
    .S0(net564),
    .S1(net540),
    .X(_05375_));
 sky130_fd_sc_hd__mux2_1 _09342_ (.A0(\core_pipeline.pipeline_registers.registers[18][21] ),
    .A1(\core_pipeline.pipeline_registers.registers[19][21] ),
    .S(net564),
    .X(_05376_));
 sky130_fd_sc_hd__a22o_1 _09343_ (.A1(\core_pipeline.pipeline_registers.registers[16][21] ),
    .A2(net279),
    .B1(net362),
    .B2(_05376_),
    .X(_05377_));
 sky130_fd_sc_hd__a211o_1 _09344_ (.A1(\core_pipeline.pipeline_registers.registers[17][21] ),
    .A2(net276),
    .B1(_05377_),
    .C1(net460),
    .X(_05378_));
 sky130_fd_sc_hd__a211o_1 _09345_ (.A1(net369),
    .A2(_05375_),
    .B1(_05378_),
    .C1(_05374_),
    .X(_05379_));
 sky130_fd_sc_hd__and3_1 _09346_ (.A(net146),
    .B(_05367_),
    .C(_05379_),
    .X(_05380_));
 sky130_fd_sc_hd__a21o_1 _09347_ (.A1(\core_pipeline.decode_to_execute_rs2_data[21] ),
    .A2(net134),
    .B1(_05380_),
    .X(_00553_));
 sky130_fd_sc_hd__mux4_1 _09348_ (.A0(\core_pipeline.pipeline_registers.registers[8][22] ),
    .A1(\core_pipeline.pipeline_registers.registers[9][22] ),
    .A2(\core_pipeline.pipeline_registers.registers[10][22] ),
    .A3(\core_pipeline.pipeline_registers.registers[11][22] ),
    .S0(net555),
    .S1(net534),
    .X(_05381_));
 sky130_fd_sc_hd__or2_1 _09349_ (.A(net522),
    .B(_05381_),
    .X(_05382_));
 sky130_fd_sc_hd__mux4_1 _09350_ (.A0(\core_pipeline.pipeline_registers.registers[12][22] ),
    .A1(\core_pipeline.pipeline_registers.registers[13][22] ),
    .A2(\core_pipeline.pipeline_registers.registers[14][22] ),
    .A3(\core_pipeline.pipeline_registers.registers[15][22] ),
    .S0(net555),
    .S1(net534),
    .X(_05383_));
 sky130_fd_sc_hd__o211a_1 _09351_ (.A1(net464),
    .A2(_05383_),
    .B1(_05382_),
    .C1(net516),
    .X(_05384_));
 sky130_fd_sc_hd__mux4_1 _09352_ (.A0(\core_pipeline.pipeline_registers.registers[4][22] ),
    .A1(\core_pipeline.pipeline_registers.registers[5][22] ),
    .A2(\core_pipeline.pipeline_registers.registers[6][22] ),
    .A3(\core_pipeline.pipeline_registers.registers[7][22] ),
    .S0(net555),
    .S1(net534),
    .X(_05385_));
 sky130_fd_sc_hd__mux2_1 _09353_ (.A0(\core_pipeline.pipeline_registers.registers[2][22] ),
    .A1(\core_pipeline.pipeline_registers.registers[3][22] ),
    .S(net555),
    .X(_05386_));
 sky130_fd_sc_hd__a22o_1 _09354_ (.A1(\core_pipeline.pipeline_registers.registers[1][22] ),
    .A2(net276),
    .B1(net361),
    .B2(_05386_),
    .X(_05387_));
 sky130_fd_sc_hd__a211o_1 _09355_ (.A1(\core_pipeline.pipeline_registers.registers[0][22] ),
    .A2(net278),
    .B1(_05387_),
    .C1(net512),
    .X(_05388_));
 sky130_fd_sc_hd__a211o_1 _09356_ (.A1(net370),
    .A2(_05385_),
    .B1(_05388_),
    .C1(_05384_),
    .X(_05389_));
 sky130_fd_sc_hd__mux2_1 _09357_ (.A0(\core_pipeline.pipeline_registers.registers[26][22] ),
    .A1(\core_pipeline.pipeline_registers.registers[27][22] ),
    .S(net555),
    .X(_05390_));
 sky130_fd_sc_hd__a221o_1 _09358_ (.A1(\core_pipeline.pipeline_registers.registers[24][22] ),
    .A2(net426),
    .B1(net365),
    .B2(\core_pipeline.pipeline_registers.registers[25][22] ),
    .C1(net522),
    .X(_05391_));
 sky130_fd_sc_hd__a21o_1 _09359_ (.A1(net536),
    .A2(_05390_),
    .B1(_05391_),
    .X(_05392_));
 sky130_fd_sc_hd__mux2_1 _09360_ (.A0(\core_pipeline.pipeline_registers.registers[30][22] ),
    .A1(\core_pipeline.pipeline_registers.registers[31][22] ),
    .S(net555),
    .X(_05393_));
 sky130_fd_sc_hd__a221o_1 _09361_ (.A1(\core_pipeline.pipeline_registers.registers[28][22] ),
    .A2(net426),
    .B1(net365),
    .B2(\core_pipeline.pipeline_registers.registers[29][22] ),
    .C1(net464),
    .X(_05394_));
 sky130_fd_sc_hd__a21o_1 _09362_ (.A1(net534),
    .A2(_05393_),
    .B1(_05394_),
    .X(_05395_));
 sky130_fd_sc_hd__mux4_1 _09363_ (.A0(\core_pipeline.pipeline_registers.registers[16][22] ),
    .A1(\core_pipeline.pipeline_registers.registers[17][22] ),
    .A2(\core_pipeline.pipeline_registers.registers[18][22] ),
    .A3(\core_pipeline.pipeline_registers.registers[19][22] ),
    .S0(net555),
    .S1(net534),
    .X(_05396_));
 sky130_fd_sc_hd__mux4_1 _09364_ (.A0(\core_pipeline.pipeline_registers.registers[20][22] ),
    .A1(\core_pipeline.pipeline_registers.registers[21][22] ),
    .A2(\core_pipeline.pipeline_registers.registers[22][22] ),
    .A3(\core_pipeline.pipeline_registers.registers[23][22] ),
    .S0(net555),
    .S1(net534),
    .X(_05397_));
 sky130_fd_sc_hd__a22o_1 _09365_ (.A1(net430),
    .A2(_05396_),
    .B1(_05397_),
    .B2(net370),
    .X(_05398_));
 sky130_fd_sc_hd__a31o_1 _09366_ (.A1(net516),
    .A2(_05392_),
    .A3(_05395_),
    .B1(net460),
    .X(_05399_));
 sky130_fd_sc_hd__o211a_1 _09367_ (.A1(_05398_),
    .A2(_05399_),
    .B1(net145),
    .C1(_05389_),
    .X(_05400_));
 sky130_fd_sc_hd__a21o_1 _09368_ (.A1(\core_pipeline.decode_to_execute_rs2_data[22] ),
    .A2(net131),
    .B1(_05400_),
    .X(_00554_));
 sky130_fd_sc_hd__mux4_1 _09369_ (.A0(\core_pipeline.pipeline_registers.registers[12][23] ),
    .A1(\core_pipeline.pipeline_registers.registers[13][23] ),
    .A2(\core_pipeline.pipeline_registers.registers[14][23] ),
    .A3(\core_pipeline.pipeline_registers.registers[15][23] ),
    .S0(net557),
    .S1(net535),
    .X(_05401_));
 sky130_fd_sc_hd__mux4_1 _09370_ (.A0(\core_pipeline.pipeline_registers.registers[8][23] ),
    .A1(\core_pipeline.pipeline_registers.registers[9][23] ),
    .A2(\core_pipeline.pipeline_registers.registers[10][23] ),
    .A3(\core_pipeline.pipeline_registers.registers[11][23] ),
    .S0(net557),
    .S1(net535),
    .X(_05402_));
 sky130_fd_sc_hd__or2_1 _09371_ (.A(net522),
    .B(_05402_),
    .X(_05403_));
 sky130_fd_sc_hd__o211a_1 _09372_ (.A1(_03329_),
    .A2(_05401_),
    .B1(_05403_),
    .C1(net517),
    .X(_05404_));
 sky130_fd_sc_hd__mux4_1 _09373_ (.A0(\core_pipeline.pipeline_registers.registers[4][23] ),
    .A1(\core_pipeline.pipeline_registers.registers[5][23] ),
    .A2(\core_pipeline.pipeline_registers.registers[6][23] ),
    .A3(\core_pipeline.pipeline_registers.registers[7][23] ),
    .S0(net557),
    .S1(net535),
    .X(_05405_));
 sky130_fd_sc_hd__mux4_1 _09374_ (.A0(\core_pipeline.pipeline_registers.registers[0][23] ),
    .A1(\core_pipeline.pipeline_registers.registers[1][23] ),
    .A2(\core_pipeline.pipeline_registers.registers[2][23] ),
    .A3(\core_pipeline.pipeline_registers.registers[3][23] ),
    .S0(net557),
    .S1(net542),
    .X(_05406_));
 sky130_fd_sc_hd__a221o_1 _09375_ (.A1(net370),
    .A2(_05405_),
    .B1(_05406_),
    .B2(net430),
    .C1(net512),
    .X(_05407_));
 sky130_fd_sc_hd__mux2_1 _09376_ (.A0(\core_pipeline.pipeline_registers.registers[30][23] ),
    .A1(\core_pipeline.pipeline_registers.registers[31][23] ),
    .S(net558),
    .X(_05408_));
 sky130_fd_sc_hd__a221o_1 _09377_ (.A1(\core_pipeline.pipeline_registers.registers[28][23] ),
    .A2(net427),
    .B1(net366),
    .B2(\core_pipeline.pipeline_registers.registers[29][23] ),
    .C1(net465),
    .X(_05409_));
 sky130_fd_sc_hd__a21o_1 _09378_ (.A1(net535),
    .A2(_05408_),
    .B1(_05409_),
    .X(_05410_));
 sky130_fd_sc_hd__mux2_1 _09379_ (.A0(\core_pipeline.pipeline_registers.registers[26][23] ),
    .A1(\core_pipeline.pipeline_registers.registers[27][23] ),
    .S(net558),
    .X(_05411_));
 sky130_fd_sc_hd__a221o_1 _09380_ (.A1(\core_pipeline.pipeline_registers.registers[24][23] ),
    .A2(net427),
    .B1(_04695_),
    .B2(\core_pipeline.pipeline_registers.registers[25][23] ),
    .C1(net522),
    .X(_05412_));
 sky130_fd_sc_hd__a21o_1 _09381_ (.A1(net535),
    .A2(_05411_),
    .B1(_05412_),
    .X(_05413_));
 sky130_fd_sc_hd__and3_1 _09382_ (.A(net517),
    .B(_05410_),
    .C(_05413_),
    .X(_05414_));
 sky130_fd_sc_hd__mux4_1 _09383_ (.A0(\core_pipeline.pipeline_registers.registers[20][23] ),
    .A1(\core_pipeline.pipeline_registers.registers[21][23] ),
    .A2(\core_pipeline.pipeline_registers.registers[22][23] ),
    .A3(\core_pipeline.pipeline_registers.registers[23][23] ),
    .S0(net557),
    .S1(net535),
    .X(_05415_));
 sky130_fd_sc_hd__a31o_1 _09384_ (.A1(\core_pipeline.pipeline_registers.registers[17][23] ),
    .A2(net430),
    .A3(net365),
    .B1(net460),
    .X(_05416_));
 sky130_fd_sc_hd__mux2_1 _09385_ (.A0(\core_pipeline.pipeline_registers.registers[18][23] ),
    .A1(\core_pipeline.pipeline_registers.registers[19][23] ),
    .S(net557),
    .X(_05417_));
 sky130_fd_sc_hd__a22o_1 _09386_ (.A1(\core_pipeline.pipeline_registers.registers[16][23] ),
    .A2(net278),
    .B1(net361),
    .B2(_05417_),
    .X(_05418_));
 sky130_fd_sc_hd__a211o_1 _09387_ (.A1(net370),
    .A2(_05415_),
    .B1(_05416_),
    .C1(_05418_),
    .X(_05419_));
 sky130_fd_sc_hd__o22a_1 _09388_ (.A1(_05404_),
    .A2(_05407_),
    .B1(_05414_),
    .B2(_05419_),
    .X(_05420_));
 sky130_fd_sc_hd__mux2_1 _09389_ (.A0(\core_pipeline.decode_to_execute_rs2_data[23] ),
    .A1(_05420_),
    .S(net141),
    .X(_00555_));
 sky130_fd_sc_hd__mux4_1 _09390_ (.A0(\core_pipeline.pipeline_registers.registers[8][24] ),
    .A1(\core_pipeline.pipeline_registers.registers[9][24] ),
    .A2(\core_pipeline.pipeline_registers.registers[10][24] ),
    .A3(\core_pipeline.pipeline_registers.registers[11][24] ),
    .S0(net550),
    .S1(net530),
    .X(_05421_));
 sky130_fd_sc_hd__or2_1 _09391_ (.A(net520),
    .B(_05421_),
    .X(_05422_));
 sky130_fd_sc_hd__mux4_1 _09392_ (.A0(\core_pipeline.pipeline_registers.registers[12][24] ),
    .A1(\core_pipeline.pipeline_registers.registers[13][24] ),
    .A2(\core_pipeline.pipeline_registers.registers[14][24] ),
    .A3(\core_pipeline.pipeline_registers.registers[15][24] ),
    .S0(net551),
    .S1(net530),
    .X(_05423_));
 sky130_fd_sc_hd__o211a_1 _09393_ (.A1(net463),
    .A2(_05423_),
    .B1(_05422_),
    .C1(net514),
    .X(_05424_));
 sky130_fd_sc_hd__mux4_1 _09394_ (.A0(\core_pipeline.pipeline_registers.registers[4][24] ),
    .A1(\core_pipeline.pipeline_registers.registers[5][24] ),
    .A2(\core_pipeline.pipeline_registers.registers[6][24] ),
    .A3(\core_pipeline.pipeline_registers.registers[7][24] ),
    .S0(net550),
    .S1(net530),
    .X(_05425_));
 sky130_fd_sc_hd__mux2_1 _09395_ (.A0(\core_pipeline.pipeline_registers.registers[2][24] ),
    .A1(\core_pipeline.pipeline_registers.registers[3][24] ),
    .S(net550),
    .X(_05426_));
 sky130_fd_sc_hd__a31o_1 _09396_ (.A1(net530),
    .A2(net429),
    .A3(_05426_),
    .B1(net511),
    .X(_05427_));
 sky130_fd_sc_hd__a221o_1 _09397_ (.A1(\core_pipeline.pipeline_registers.registers[0][24] ),
    .A2(net279),
    .B1(net277),
    .B2(\core_pipeline.pipeline_registers.registers[1][24] ),
    .C1(_05427_),
    .X(_05428_));
 sky130_fd_sc_hd__a211o_1 _09398_ (.A1(net368),
    .A2(_05425_),
    .B1(_05428_),
    .C1(_05424_),
    .X(_05429_));
 sky130_fd_sc_hd__mux2_1 _09399_ (.A0(\core_pipeline.pipeline_registers.registers[30][24] ),
    .A1(\core_pipeline.pipeline_registers.registers[31][24] ),
    .S(net557),
    .X(_05430_));
 sky130_fd_sc_hd__a221o_1 _09400_ (.A1(\core_pipeline.pipeline_registers.registers[28][24] ),
    .A2(net425),
    .B1(net364),
    .B2(\core_pipeline.pipeline_registers.registers[29][24] ),
    .C1(net462),
    .X(_05431_));
 sky130_fd_sc_hd__a21o_1 _09401_ (.A1(net530),
    .A2(_05430_),
    .B1(_05431_),
    .X(_05432_));
 sky130_fd_sc_hd__mux2_1 _09402_ (.A0(\core_pipeline.pipeline_registers.registers[26][24] ),
    .A1(\core_pipeline.pipeline_registers.registers[27][24] ),
    .S(net550),
    .X(_05433_));
 sky130_fd_sc_hd__a221o_1 _09403_ (.A1(\core_pipeline.pipeline_registers.registers[24][24] ),
    .A2(_04681_),
    .B1(net363),
    .B2(\core_pipeline.pipeline_registers.registers[25][24] ),
    .C1(net520),
    .X(_05434_));
 sky130_fd_sc_hd__a21o_1 _09404_ (.A1(net530),
    .A2(_05433_),
    .B1(_05434_),
    .X(_05435_));
 sky130_fd_sc_hd__and3_1 _09405_ (.A(net515),
    .B(_05432_),
    .C(_05435_),
    .X(_05436_));
 sky130_fd_sc_hd__mux4_1 _09406_ (.A0(\core_pipeline.pipeline_registers.registers[20][24] ),
    .A1(\core_pipeline.pipeline_registers.registers[21][24] ),
    .A2(\core_pipeline.pipeline_registers.registers[22][24] ),
    .A3(\core_pipeline.pipeline_registers.registers[23][24] ),
    .S0(net550),
    .S1(net530),
    .X(_05437_));
 sky130_fd_sc_hd__mux2_1 _09407_ (.A0(\core_pipeline.pipeline_registers.registers[18][24] ),
    .A1(\core_pipeline.pipeline_registers.registers[19][24] ),
    .S(net550),
    .X(_05438_));
 sky130_fd_sc_hd__a22o_1 _09408_ (.A1(\core_pipeline.pipeline_registers.registers[16][24] ),
    .A2(net279),
    .B1(net361),
    .B2(_05438_),
    .X(_05439_));
 sky130_fd_sc_hd__a211o_1 _09409_ (.A1(\core_pipeline.pipeline_registers.registers[17][24] ),
    .A2(net277),
    .B1(_05439_),
    .C1(net461),
    .X(_05440_));
 sky130_fd_sc_hd__a211o_1 _09410_ (.A1(net368),
    .A2(_05437_),
    .B1(_05440_),
    .C1(_05436_),
    .X(_05441_));
 sky130_fd_sc_hd__and3_1 _09411_ (.A(net141),
    .B(_05429_),
    .C(_05441_),
    .X(_05442_));
 sky130_fd_sc_hd__a21o_1 _09412_ (.A1(\core_pipeline.decode_to_execute_rs2_data[24] ),
    .A2(net124),
    .B1(_05442_),
    .X(_00556_));
 sky130_fd_sc_hd__mux4_1 _09413_ (.A0(\core_pipeline.pipeline_registers.registers[8][25] ),
    .A1(\core_pipeline.pipeline_registers.registers[9][25] ),
    .A2(\core_pipeline.pipeline_registers.registers[10][25] ),
    .A3(\core_pipeline.pipeline_registers.registers[11][25] ),
    .S0(net546),
    .S1(net532),
    .X(_05443_));
 sky130_fd_sc_hd__or2_1 _09414_ (.A(net521),
    .B(_05443_),
    .X(_05444_));
 sky130_fd_sc_hd__mux4_1 _09415_ (.A0(\core_pipeline.pipeline_registers.registers[12][25] ),
    .A1(\core_pipeline.pipeline_registers.registers[13][25] ),
    .A2(\core_pipeline.pipeline_registers.registers[14][25] ),
    .A3(\core_pipeline.pipeline_registers.registers[15][25] ),
    .S0(net552),
    .S1(net532),
    .X(_05445_));
 sky130_fd_sc_hd__o211a_1 _09416_ (.A1(net463),
    .A2(_05445_),
    .B1(_05444_),
    .C1(net515),
    .X(_05446_));
 sky130_fd_sc_hd__mux4_1 _09417_ (.A0(\core_pipeline.pipeline_registers.registers[4][25] ),
    .A1(\core_pipeline.pipeline_registers.registers[5][25] ),
    .A2(\core_pipeline.pipeline_registers.registers[6][25] ),
    .A3(\core_pipeline.pipeline_registers.registers[7][25] ),
    .S0(net552),
    .S1(net532),
    .X(_05447_));
 sky130_fd_sc_hd__mux2_1 _09418_ (.A0(\core_pipeline.pipeline_registers.registers[2][25] ),
    .A1(\core_pipeline.pipeline_registers.registers[3][25] ),
    .S(net552),
    .X(_05448_));
 sky130_fd_sc_hd__a31o_1 _09419_ (.A1(net532),
    .A2(net429),
    .A3(_05448_),
    .B1(net511),
    .X(_05449_));
 sky130_fd_sc_hd__a221o_1 _09420_ (.A1(\core_pipeline.pipeline_registers.registers[0][25] ),
    .A2(net279),
    .B1(net277),
    .B2(\core_pipeline.pipeline_registers.registers[1][25] ),
    .C1(_05449_),
    .X(_05450_));
 sky130_fd_sc_hd__a211o_1 _09421_ (.A1(net368),
    .A2(_05447_),
    .B1(_05450_),
    .C1(_05446_),
    .X(_05451_));
 sky130_fd_sc_hd__mux2_1 _09422_ (.A0(\core_pipeline.pipeline_registers.registers[26][25] ),
    .A1(\core_pipeline.pipeline_registers.registers[27][25] ),
    .S(net547),
    .X(_05452_));
 sky130_fd_sc_hd__a221o_1 _09423_ (.A1(\core_pipeline.pipeline_registers.registers[24][25] ),
    .A2(net425),
    .B1(_04695_),
    .B2(\core_pipeline.pipeline_registers.registers[25][25] ),
    .C1(net519),
    .X(_05453_));
 sky130_fd_sc_hd__a21o_1 _09424_ (.A1(net527),
    .A2(_05452_),
    .B1(_05453_),
    .X(_05454_));
 sky130_fd_sc_hd__mux2_1 _09425_ (.A0(\core_pipeline.pipeline_registers.registers[30][25] ),
    .A1(\core_pipeline.pipeline_registers.registers[31][25] ),
    .S(net547),
    .X(_05455_));
 sky130_fd_sc_hd__a221o_1 _09426_ (.A1(\core_pipeline.pipeline_registers.registers[28][25] ),
    .A2(net425),
    .B1(net364),
    .B2(\core_pipeline.pipeline_registers.registers[29][25] ),
    .C1(net463),
    .X(_05456_));
 sky130_fd_sc_hd__a21o_1 _09427_ (.A1(net527),
    .A2(_05455_),
    .B1(_05456_),
    .X(_05457_));
 sky130_fd_sc_hd__mux4_1 _09428_ (.A0(\core_pipeline.pipeline_registers.registers[16][25] ),
    .A1(\core_pipeline.pipeline_registers.registers[17][25] ),
    .A2(\core_pipeline.pipeline_registers.registers[18][25] ),
    .A3(\core_pipeline.pipeline_registers.registers[19][25] ),
    .S0(net546),
    .S1(net526),
    .X(_05458_));
 sky130_fd_sc_hd__mux4_1 _09429_ (.A0(\core_pipeline.pipeline_registers.registers[20][25] ),
    .A1(\core_pipeline.pipeline_registers.registers[21][25] ),
    .A2(\core_pipeline.pipeline_registers.registers[22][25] ),
    .A3(\core_pipeline.pipeline_registers.registers[23][25] ),
    .S0(net546),
    .S1(net526),
    .X(_05459_));
 sky130_fd_sc_hd__a22o_1 _09430_ (.A1(net428),
    .A2(_05458_),
    .B1(_05459_),
    .B2(net367),
    .X(_05460_));
 sky130_fd_sc_hd__a31o_1 _09431_ (.A1(net515),
    .A2(_05454_),
    .A3(_05457_),
    .B1(net461),
    .X(_05461_));
 sky130_fd_sc_hd__o211a_1 _09432_ (.A1(_05460_),
    .A2(_05461_),
    .B1(net139),
    .C1(_05451_),
    .X(_05462_));
 sky130_fd_sc_hd__a21o_1 _09433_ (.A1(\core_pipeline.decode_to_execute_rs2_data[25] ),
    .A2(net121),
    .B1(_05462_),
    .X(_00557_));
 sky130_fd_sc_hd__mux4_1 _09434_ (.A0(\core_pipeline.pipeline_registers.registers[8][26] ),
    .A1(\core_pipeline.pipeline_registers.registers[9][26] ),
    .A2(\core_pipeline.pipeline_registers.registers[10][26] ),
    .A3(\core_pipeline.pipeline_registers.registers[11][26] ),
    .S0(net552),
    .S1(net532),
    .X(_05463_));
 sky130_fd_sc_hd__or2_1 _09435_ (.A(net521),
    .B(_05463_),
    .X(_05464_));
 sky130_fd_sc_hd__mux4_1 _09436_ (.A0(\core_pipeline.pipeline_registers.registers[12][26] ),
    .A1(\core_pipeline.pipeline_registers.registers[13][26] ),
    .A2(\core_pipeline.pipeline_registers.registers[14][26] ),
    .A3(\core_pipeline.pipeline_registers.registers[15][26] ),
    .S0(net552),
    .S1(net532),
    .X(_05465_));
 sky130_fd_sc_hd__o211a_1 _09437_ (.A1(net463),
    .A2(_05465_),
    .B1(_05464_),
    .C1(\core_pipeline.decode_to_csr_read_address[3] ),
    .X(_05466_));
 sky130_fd_sc_hd__mux4_1 _09438_ (.A0(\core_pipeline.pipeline_registers.registers[0][26] ),
    .A1(\core_pipeline.pipeline_registers.registers[1][26] ),
    .A2(\core_pipeline.pipeline_registers.registers[2][26] ),
    .A3(\core_pipeline.pipeline_registers.registers[3][26] ),
    .S0(net554),
    .S1(net533),
    .X(_05467_));
 sky130_fd_sc_hd__mux4_1 _09439_ (.A0(\core_pipeline.pipeline_registers.registers[4][26] ),
    .A1(\core_pipeline.pipeline_registers.registers[5][26] ),
    .A2(\core_pipeline.pipeline_registers.registers[6][26] ),
    .A3(\core_pipeline.pipeline_registers.registers[7][26] ),
    .S0(net552),
    .S1(net533),
    .X(_05468_));
 sky130_fd_sc_hd__a221o_1 _09440_ (.A1(net428),
    .A2(_05467_),
    .B1(_05468_),
    .B2(net367),
    .C1(_05466_),
    .X(_05469_));
 sky130_fd_sc_hd__mux2_1 _09441_ (.A0(\core_pipeline.pipeline_registers.registers[26][26] ),
    .A1(\core_pipeline.pipeline_registers.registers[27][26] ),
    .S(net553),
    .X(_05470_));
 sky130_fd_sc_hd__a221o_1 _09442_ (.A1(\core_pipeline.pipeline_registers.registers[24][26] ),
    .A2(net425),
    .B1(net364),
    .B2(\core_pipeline.pipeline_registers.registers[25][26] ),
    .C1(net521),
    .X(_05471_));
 sky130_fd_sc_hd__a21o_1 _09443_ (.A1(net532),
    .A2(_05470_),
    .B1(_05471_),
    .X(_05472_));
 sky130_fd_sc_hd__mux2_1 _09444_ (.A0(\core_pipeline.pipeline_registers.registers[30][26] ),
    .A1(\core_pipeline.pipeline_registers.registers[31][26] ),
    .S(net552),
    .X(_05473_));
 sky130_fd_sc_hd__a221o_1 _09445_ (.A1(\core_pipeline.pipeline_registers.registers[28][26] ),
    .A2(net425),
    .B1(net364),
    .B2(\core_pipeline.pipeline_registers.registers[29][26] ),
    .C1(net462),
    .X(_05474_));
 sky130_fd_sc_hd__a21o_1 _09446_ (.A1(net532),
    .A2(_05473_),
    .B1(_05474_),
    .X(_05475_));
 sky130_fd_sc_hd__mux4_1 _09447_ (.A0(\core_pipeline.pipeline_registers.registers[16][26] ),
    .A1(\core_pipeline.pipeline_registers.registers[17][26] ),
    .A2(\core_pipeline.pipeline_registers.registers[18][26] ),
    .A3(\core_pipeline.pipeline_registers.registers[19][26] ),
    .S0(net553),
    .S1(net533),
    .X(_05476_));
 sky130_fd_sc_hd__mux4_1 _09448_ (.A0(\core_pipeline.pipeline_registers.registers[20][26] ),
    .A1(\core_pipeline.pipeline_registers.registers[21][26] ),
    .A2(\core_pipeline.pipeline_registers.registers[22][26] ),
    .A3(\core_pipeline.pipeline_registers.registers[23][26] ),
    .S0(net553),
    .S1(net533),
    .X(_05477_));
 sky130_fd_sc_hd__a22o_1 _09449_ (.A1(net428),
    .A2(_05476_),
    .B1(_05477_),
    .B2(net367),
    .X(_05478_));
 sky130_fd_sc_hd__a31o_1 _09450_ (.A1(net515),
    .A2(_05472_),
    .A3(_05475_),
    .B1(net461),
    .X(_05479_));
 sky130_fd_sc_hd__o22a_1 _09451_ (.A1(\core_pipeline.decode_to_csr_read_address[4] ),
    .A2(_05469_),
    .B1(_05478_),
    .B2(_05479_),
    .X(_05480_));
 sky130_fd_sc_hd__mux2_1 _09452_ (.A0(\core_pipeline.decode_to_execute_rs2_data[26] ),
    .A1(_05480_),
    .S(net139),
    .X(_00558_));
 sky130_fd_sc_hd__and2_1 _09453_ (.A(\core_pipeline.decode_to_execute_rs2_data[27] ),
    .B(net134),
    .X(_05481_));
 sky130_fd_sc_hd__mux2_1 _09454_ (.A0(\core_pipeline.pipeline_registers.registers[30][27] ),
    .A1(\core_pipeline.pipeline_registers.registers[31][27] ),
    .S(net563),
    .X(_05482_));
 sky130_fd_sc_hd__a221o_1 _09455_ (.A1(\core_pipeline.pipeline_registers.registers[28][27] ),
    .A2(net427),
    .B1(net366),
    .B2(\core_pipeline.pipeline_registers.registers[29][27] ),
    .C1(net465),
    .X(_05483_));
 sky130_fd_sc_hd__a21o_1 _09456_ (.A1(net540),
    .A2(_05482_),
    .B1(_05483_),
    .X(_05484_));
 sky130_fd_sc_hd__mux2_1 _09457_ (.A0(\core_pipeline.pipeline_registers.registers[26][27] ),
    .A1(\core_pipeline.pipeline_registers.registers[27][27] ),
    .S(net563),
    .X(_05485_));
 sky130_fd_sc_hd__a221o_1 _09458_ (.A1(\core_pipeline.pipeline_registers.registers[24][27] ),
    .A2(net427),
    .B1(net366),
    .B2(\core_pipeline.pipeline_registers.registers[25][27] ),
    .C1(net524),
    .X(_05486_));
 sky130_fd_sc_hd__a21o_1 _09459_ (.A1(net540),
    .A2(_05485_),
    .B1(_05486_),
    .X(_05487_));
 sky130_fd_sc_hd__mux4_1 _09460_ (.A0(\core_pipeline.pipeline_registers.registers[20][27] ),
    .A1(\core_pipeline.pipeline_registers.registers[21][27] ),
    .A2(\core_pipeline.pipeline_registers.registers[22][27] ),
    .A3(\core_pipeline.pipeline_registers.registers[23][27] ),
    .S0(net563),
    .S1(net540),
    .X(_05488_));
 sky130_fd_sc_hd__mux4_1 _09461_ (.A0(\core_pipeline.pipeline_registers.registers[16][27] ),
    .A1(\core_pipeline.pipeline_registers.registers[17][27] ),
    .A2(\core_pipeline.pipeline_registers.registers[18][27] ),
    .A3(\core_pipeline.pipeline_registers.registers[19][27] ),
    .S0(net563),
    .S1(net540),
    .X(_05489_));
 sky130_fd_sc_hd__a221o_1 _09462_ (.A1(net369),
    .A2(_05488_),
    .B1(_05489_),
    .B2(net430),
    .C1(_03330_),
    .X(_05490_));
 sky130_fd_sc_hd__a31o_1 _09463_ (.A1(net517),
    .A2(_05484_),
    .A3(_05487_),
    .B1(_05490_),
    .X(_05491_));
 sky130_fd_sc_hd__mux4_1 _09464_ (.A0(\core_pipeline.pipeline_registers.registers[12][27] ),
    .A1(\core_pipeline.pipeline_registers.registers[13][27] ),
    .A2(\core_pipeline.pipeline_registers.registers[14][27] ),
    .A3(\core_pipeline.pipeline_registers.registers[15][27] ),
    .S0(net563),
    .S1(net540),
    .X(_05492_));
 sky130_fd_sc_hd__mux4_1 _09465_ (.A0(\core_pipeline.pipeline_registers.registers[8][27] ),
    .A1(\core_pipeline.pipeline_registers.registers[9][27] ),
    .A2(\core_pipeline.pipeline_registers.registers[10][27] ),
    .A3(\core_pipeline.pipeline_registers.registers[11][27] ),
    .S0(net563),
    .S1(net541),
    .X(_05493_));
 sky130_fd_sc_hd__or2_1 _09466_ (.A(net524),
    .B(_05493_),
    .X(_05494_));
 sky130_fd_sc_hd__o211a_1 _09467_ (.A1(net465),
    .A2(_05492_),
    .B1(_05494_),
    .C1(net517),
    .X(_05495_));
 sky130_fd_sc_hd__mux4_1 _09468_ (.A0(\core_pipeline.pipeline_registers.registers[4][27] ),
    .A1(\core_pipeline.pipeline_registers.registers[5][27] ),
    .A2(\core_pipeline.pipeline_registers.registers[6][27] ),
    .A3(\core_pipeline.pipeline_registers.registers[7][27] ),
    .S0(net564),
    .S1(net541),
    .X(_05496_));
 sky130_fd_sc_hd__mux2_1 _09469_ (.A0(\core_pipeline.pipeline_registers.registers[2][27] ),
    .A1(\core_pipeline.pipeline_registers.registers[3][27] ),
    .S(net563),
    .X(_05497_));
 sky130_fd_sc_hd__a22o_1 _09470_ (.A1(\core_pipeline.pipeline_registers.registers[1][27] ),
    .A2(net276),
    .B1(net362),
    .B2(_05497_),
    .X(_05498_));
 sky130_fd_sc_hd__a211o_1 _09471_ (.A1(\core_pipeline.pipeline_registers.registers[0][27] ),
    .A2(net279),
    .B1(_05498_),
    .C1(net512),
    .X(_05499_));
 sky130_fd_sc_hd__a211o_1 _09472_ (.A1(net369),
    .A2(_05496_),
    .B1(_05499_),
    .C1(_05495_),
    .X(_05500_));
 sky130_fd_sc_hd__a31o_1 _09473_ (.A1(net148),
    .A2(_05491_),
    .A3(_05500_),
    .B1(_05481_),
    .X(_00559_));
 sky130_fd_sc_hd__mux4_1 _09474_ (.A0(\core_pipeline.pipeline_registers.registers[12][28] ),
    .A1(\core_pipeline.pipeline_registers.registers[13][28] ),
    .A2(\core_pipeline.pipeline_registers.registers[14][28] ),
    .A3(\core_pipeline.pipeline_registers.registers[15][28] ),
    .S0(net562),
    .S1(net538),
    .X(_05501_));
 sky130_fd_sc_hd__mux4_1 _09475_ (.A0(\core_pipeline.pipeline_registers.registers[8][28] ),
    .A1(\core_pipeline.pipeline_registers.registers[9][28] ),
    .A2(\core_pipeline.pipeline_registers.registers[10][28] ),
    .A3(\core_pipeline.pipeline_registers.registers[11][28] ),
    .S0(net562),
    .S1(net538),
    .X(_05502_));
 sky130_fd_sc_hd__or2_1 _09476_ (.A(net523),
    .B(_05502_),
    .X(_05503_));
 sky130_fd_sc_hd__o211a_1 _09477_ (.A1(net465),
    .A2(_05501_),
    .B1(_05503_),
    .C1(net518),
    .X(_05504_));
 sky130_fd_sc_hd__mux4_1 _09478_ (.A0(\core_pipeline.pipeline_registers.registers[4][28] ),
    .A1(\core_pipeline.pipeline_registers.registers[5][28] ),
    .A2(\core_pipeline.pipeline_registers.registers[6][28] ),
    .A3(\core_pipeline.pipeline_registers.registers[7][28] ),
    .S0(net562),
    .S1(net539),
    .X(_05505_));
 sky130_fd_sc_hd__mux4_1 _09479_ (.A0(\core_pipeline.pipeline_registers.registers[0][28] ),
    .A1(\core_pipeline.pipeline_registers.registers[1][28] ),
    .A2(\core_pipeline.pipeline_registers.registers[2][28] ),
    .A3(\core_pipeline.pipeline_registers.registers[3][28] ),
    .S0(net561),
    .S1(net538),
    .X(_05506_));
 sky130_fd_sc_hd__a221o_1 _09480_ (.A1(net369),
    .A2(_05505_),
    .B1(_05506_),
    .B2(net430),
    .C1(net512),
    .X(_05507_));
 sky130_fd_sc_hd__mux2_1 _09481_ (.A0(\core_pipeline.pipeline_registers.registers[30][28] ),
    .A1(\core_pipeline.pipeline_registers.registers[31][28] ),
    .S(net560),
    .X(_05508_));
 sky130_fd_sc_hd__a221o_1 _09482_ (.A1(\core_pipeline.pipeline_registers.registers[28][28] ),
    .A2(net427),
    .B1(net365),
    .B2(\core_pipeline.pipeline_registers.registers[29][28] ),
    .C1(net465),
    .X(_05509_));
 sky130_fd_sc_hd__a21o_1 _09483_ (.A1(net539),
    .A2(_05508_),
    .B1(_05509_),
    .X(_05510_));
 sky130_fd_sc_hd__mux2_1 _09484_ (.A0(\core_pipeline.pipeline_registers.registers[26][28] ),
    .A1(\core_pipeline.pipeline_registers.registers[27][28] ),
    .S(net559),
    .X(_05511_));
 sky130_fd_sc_hd__a221o_1 _09485_ (.A1(\core_pipeline.pipeline_registers.registers[24][28] ),
    .A2(net426),
    .B1(net365),
    .B2(\core_pipeline.pipeline_registers.registers[25][28] ),
    .C1(net523),
    .X(_05512_));
 sky130_fd_sc_hd__a21o_1 _09486_ (.A1(net538),
    .A2(_05511_),
    .B1(_05512_),
    .X(_05513_));
 sky130_fd_sc_hd__and3_1 _09487_ (.A(net518),
    .B(_05510_),
    .C(_05513_),
    .X(_05514_));
 sky130_fd_sc_hd__mux4_1 _09488_ (.A0(\core_pipeline.pipeline_registers.registers[20][28] ),
    .A1(\core_pipeline.pipeline_registers.registers[21][28] ),
    .A2(\core_pipeline.pipeline_registers.registers[22][28] ),
    .A3(\core_pipeline.pipeline_registers.registers[23][28] ),
    .S0(net562),
    .S1(net538),
    .X(_05515_));
 sky130_fd_sc_hd__a31o_1 _09489_ (.A1(\core_pipeline.pipeline_registers.registers[17][28] ),
    .A2(_04680_),
    .A3(net365),
    .B1(net460),
    .X(_05516_));
 sky130_fd_sc_hd__mux2_1 _09490_ (.A0(\core_pipeline.pipeline_registers.registers[18][28] ),
    .A1(\core_pipeline.pipeline_registers.registers[19][28] ),
    .S(net562),
    .X(_05517_));
 sky130_fd_sc_hd__a22o_1 _09491_ (.A1(\core_pipeline.pipeline_registers.registers[16][28] ),
    .A2(net278),
    .B1(net362),
    .B2(_05517_),
    .X(_05518_));
 sky130_fd_sc_hd__a211o_1 _09492_ (.A1(net369),
    .A2(_05515_),
    .B1(_05516_),
    .C1(_05518_),
    .X(_05519_));
 sky130_fd_sc_hd__o22a_1 _09493_ (.A1(_05504_),
    .A2(_05507_),
    .B1(_05514_),
    .B2(_05519_),
    .X(_05520_));
 sky130_fd_sc_hd__mux2_1 _09494_ (.A0(\core_pipeline.decode_to_execute_rs2_data[28] ),
    .A1(_05520_),
    .S(net145),
    .X(_00560_));
 sky130_fd_sc_hd__mux4_1 _09495_ (.A0(\core_pipeline.pipeline_registers.registers[8][29] ),
    .A1(\core_pipeline.pipeline_registers.registers[9][29] ),
    .A2(\core_pipeline.pipeline_registers.registers[10][29] ),
    .A3(\core_pipeline.pipeline_registers.registers[11][29] ),
    .S0(net558),
    .S1(net535),
    .X(_05521_));
 sky130_fd_sc_hd__or2_1 _09496_ (.A(net522),
    .B(_05521_),
    .X(_05522_));
 sky130_fd_sc_hd__mux4_1 _09497_ (.A0(\core_pipeline.pipeline_registers.registers[12][29] ),
    .A1(\core_pipeline.pipeline_registers.registers[13][29] ),
    .A2(\core_pipeline.pipeline_registers.registers[14][29] ),
    .A3(\core_pipeline.pipeline_registers.registers[15][29] ),
    .S0(net558),
    .S1(net536),
    .X(_05523_));
 sky130_fd_sc_hd__o211a_1 _09498_ (.A1(_03329_),
    .A2(_05523_),
    .B1(_05522_),
    .C1(net516),
    .X(_05524_));
 sky130_fd_sc_hd__mux4_1 _09499_ (.A0(\core_pipeline.pipeline_registers.registers[4][29] ),
    .A1(\core_pipeline.pipeline_registers.registers[5][29] ),
    .A2(\core_pipeline.pipeline_registers.registers[6][29] ),
    .A3(\core_pipeline.pipeline_registers.registers[7][29] ),
    .S0(net557),
    .S1(net535),
    .X(_05525_));
 sky130_fd_sc_hd__mux2_1 _09500_ (.A0(\core_pipeline.pipeline_registers.registers[2][29] ),
    .A1(\core_pipeline.pipeline_registers.registers[3][29] ),
    .S(net557),
    .X(_05526_));
 sky130_fd_sc_hd__a31o_1 _09501_ (.A1(net535),
    .A2(net430),
    .A3(_05526_),
    .B1(net512),
    .X(_05527_));
 sky130_fd_sc_hd__a221o_1 _09502_ (.A1(\core_pipeline.pipeline_registers.registers[0][29] ),
    .A2(net278),
    .B1(net277),
    .B2(\core_pipeline.pipeline_registers.registers[1][29] ),
    .C1(_05527_),
    .X(_05528_));
 sky130_fd_sc_hd__a211o_1 _09503_ (.A1(net370),
    .A2(_05525_),
    .B1(_05528_),
    .C1(_05524_),
    .X(_05529_));
 sky130_fd_sc_hd__mux2_1 _09504_ (.A0(\core_pipeline.pipeline_registers.registers[30][29] ),
    .A1(\core_pipeline.pipeline_registers.registers[31][29] ),
    .S(net557),
    .X(_05530_));
 sky130_fd_sc_hd__a221o_1 _09505_ (.A1(\core_pipeline.pipeline_registers.registers[28][29] ),
    .A2(net426),
    .B1(net365),
    .B2(\core_pipeline.pipeline_registers.registers[29][29] ),
    .C1(net464),
    .X(_05531_));
 sky130_fd_sc_hd__a21o_1 _09506_ (.A1(net535),
    .A2(_05530_),
    .B1(_05531_),
    .X(_05532_));
 sky130_fd_sc_hd__mux2_1 _09507_ (.A0(\core_pipeline.pipeline_registers.registers[26][29] ),
    .A1(\core_pipeline.pipeline_registers.registers[27][29] ),
    .S(net557),
    .X(_05533_));
 sky130_fd_sc_hd__a221o_1 _09508_ (.A1(\core_pipeline.pipeline_registers.registers[24][29] ),
    .A2(net426),
    .B1(net365),
    .B2(\core_pipeline.pipeline_registers.registers[25][29] ),
    .C1(net522),
    .X(_05534_));
 sky130_fd_sc_hd__a21o_1 _09509_ (.A1(net535),
    .A2(_05533_),
    .B1(_05534_),
    .X(_05535_));
 sky130_fd_sc_hd__and3_1 _09510_ (.A(net516),
    .B(_05532_),
    .C(_05535_),
    .X(_05536_));
 sky130_fd_sc_hd__mux4_1 _09511_ (.A0(\core_pipeline.pipeline_registers.registers[20][29] ),
    .A1(\core_pipeline.pipeline_registers.registers[21][29] ),
    .A2(\core_pipeline.pipeline_registers.registers[22][29] ),
    .A3(\core_pipeline.pipeline_registers.registers[23][29] ),
    .S0(net558),
    .S1(net536),
    .X(_05537_));
 sky130_fd_sc_hd__mux2_1 _09512_ (.A0(\core_pipeline.pipeline_registers.registers[18][29] ),
    .A1(\core_pipeline.pipeline_registers.registers[19][29] ),
    .S(net558),
    .X(_05538_));
 sky130_fd_sc_hd__a22o_1 _09513_ (.A1(\core_pipeline.pipeline_registers.registers[17][29] ),
    .A2(net276),
    .B1(net362),
    .B2(_05538_),
    .X(_05539_));
 sky130_fd_sc_hd__a211o_1 _09514_ (.A1(\core_pipeline.pipeline_registers.registers[16][29] ),
    .A2(net278),
    .B1(_05539_),
    .C1(net460),
    .X(_05540_));
 sky130_fd_sc_hd__a211o_1 _09515_ (.A1(net370),
    .A2(_05537_),
    .B1(_05540_),
    .C1(_05536_),
    .X(_05541_));
 sky130_fd_sc_hd__and3_1 _09516_ (.A(net145),
    .B(_05529_),
    .C(_05541_),
    .X(_05542_));
 sky130_fd_sc_hd__a21o_1 _09517_ (.A1(\core_pipeline.decode_to_execute_rs2_data[29] ),
    .A2(net131),
    .B1(_05542_),
    .X(_00561_));
 sky130_fd_sc_hd__mux2_1 _09518_ (.A0(\core_pipeline.pipeline_registers.registers[30][30] ),
    .A1(\core_pipeline.pipeline_registers.registers[31][30] ),
    .S(net555),
    .X(_05543_));
 sky130_fd_sc_hd__a221o_1 _09519_ (.A1(\core_pipeline.pipeline_registers.registers[28][30] ),
    .A2(net426),
    .B1(net365),
    .B2(\core_pipeline.pipeline_registers.registers[29][30] ),
    .C1(net464),
    .X(_05544_));
 sky130_fd_sc_hd__a21o_1 _09520_ (.A1(net534),
    .A2(_05543_),
    .B1(_05544_),
    .X(_05545_));
 sky130_fd_sc_hd__mux2_1 _09521_ (.A0(\core_pipeline.pipeline_registers.registers[26][30] ),
    .A1(\core_pipeline.pipeline_registers.registers[27][30] ),
    .S(net555),
    .X(_05546_));
 sky130_fd_sc_hd__a221o_1 _09522_ (.A1(\core_pipeline.pipeline_registers.registers[24][30] ),
    .A2(net426),
    .B1(net364),
    .B2(\core_pipeline.pipeline_registers.registers[25][30] ),
    .C1(net522),
    .X(_05547_));
 sky130_fd_sc_hd__a21o_1 _09523_ (.A1(net534),
    .A2(_05546_),
    .B1(_05547_),
    .X(_05548_));
 sky130_fd_sc_hd__and3_1 _09524_ (.A(net516),
    .B(_05545_),
    .C(_05548_),
    .X(_05549_));
 sky130_fd_sc_hd__mux4_1 _09525_ (.A0(\core_pipeline.pipeline_registers.registers[20][30] ),
    .A1(\core_pipeline.pipeline_registers.registers[21][30] ),
    .A2(\core_pipeline.pipeline_registers.registers[22][30] ),
    .A3(\core_pipeline.pipeline_registers.registers[23][30] ),
    .S0(net557),
    .S1(net535),
    .X(_05550_));
 sky130_fd_sc_hd__mux2_1 _09526_ (.A0(\core_pipeline.pipeline_registers.registers[18][30] ),
    .A1(\core_pipeline.pipeline_registers.registers[19][30] ),
    .S(net557),
    .X(_05551_));
 sky130_fd_sc_hd__a22o_1 _09527_ (.A1(\core_pipeline.pipeline_registers.registers[16][30] ),
    .A2(net278),
    .B1(net361),
    .B2(_05551_),
    .X(_05552_));
 sky130_fd_sc_hd__a211o_1 _09528_ (.A1(\core_pipeline.pipeline_registers.registers[17][30] ),
    .A2(net276),
    .B1(_05552_),
    .C1(net460),
    .X(_05553_));
 sky130_fd_sc_hd__a211o_1 _09529_ (.A1(net370),
    .A2(_05550_),
    .B1(_05553_),
    .C1(_05549_),
    .X(_05554_));
 sky130_fd_sc_hd__mux4_1 _09530_ (.A0(\core_pipeline.pipeline_registers.registers[12][30] ),
    .A1(\core_pipeline.pipeline_registers.registers[13][30] ),
    .A2(\core_pipeline.pipeline_registers.registers[14][30] ),
    .A3(\core_pipeline.pipeline_registers.registers[15][30] ),
    .S0(net551),
    .S1(net531),
    .X(_05555_));
 sky130_fd_sc_hd__mux4_1 _09531_ (.A0(\core_pipeline.pipeline_registers.registers[8][30] ),
    .A1(\core_pipeline.pipeline_registers.registers[9][30] ),
    .A2(\core_pipeline.pipeline_registers.registers[10][30] ),
    .A3(\core_pipeline.pipeline_registers.registers[11][30] ),
    .S0(net555),
    .S1(net535),
    .X(_05556_));
 sky130_fd_sc_hd__or2_1 _09532_ (.A(net522),
    .B(_05556_),
    .X(_05557_));
 sky130_fd_sc_hd__o211a_1 _09533_ (.A1(net464),
    .A2(_05555_),
    .B1(_05557_),
    .C1(net516),
    .X(_05558_));
 sky130_fd_sc_hd__mux4_1 _09534_ (.A0(\core_pipeline.pipeline_registers.registers[4][30] ),
    .A1(\core_pipeline.pipeline_registers.registers[5][30] ),
    .A2(\core_pipeline.pipeline_registers.registers[6][30] ),
    .A3(\core_pipeline.pipeline_registers.registers[7][30] ),
    .S0(net557),
    .S1(net535),
    .X(_05559_));
 sky130_fd_sc_hd__mux2_1 _09535_ (.A0(\core_pipeline.pipeline_registers.registers[2][30] ),
    .A1(\core_pipeline.pipeline_registers.registers[3][30] ),
    .S(net557),
    .X(_05560_));
 sky130_fd_sc_hd__a221o_1 _09536_ (.A1(\core_pipeline.pipeline_registers.registers[0][30] ),
    .A2(net279),
    .B1(net277),
    .B2(\core_pipeline.pipeline_registers.registers[1][30] ),
    .C1(net511),
    .X(_05561_));
 sky130_fd_sc_hd__a21o_1 _09537_ (.A1(net370),
    .A2(_05559_),
    .B1(_05561_),
    .X(_05562_));
 sky130_fd_sc_hd__a211o_1 _09538_ (.A1(net361),
    .A2(_05560_),
    .B1(_05562_),
    .C1(_05558_),
    .X(_05563_));
 sky130_fd_sc_hd__and3_1 _09539_ (.A(net144),
    .B(_05554_),
    .C(_05563_),
    .X(_05564_));
 sky130_fd_sc_hd__a21o_1 _09540_ (.A1(\core_pipeline.decode_to_execute_rs2_data[30] ),
    .A2(net125),
    .B1(_05564_),
    .X(_00562_));
 sky130_fd_sc_hd__mux4_1 _09541_ (.A0(\core_pipeline.pipeline_registers.registers[12][31] ),
    .A1(\core_pipeline.pipeline_registers.registers[13][31] ),
    .A2(\core_pipeline.pipeline_registers.registers[14][31] ),
    .A3(\core_pipeline.pipeline_registers.registers[15][31] ),
    .S0(net563),
    .S1(net540),
    .X(_05565_));
 sky130_fd_sc_hd__mux4_1 _09542_ (.A0(\core_pipeline.pipeline_registers.registers[8][31] ),
    .A1(\core_pipeline.pipeline_registers.registers[9][31] ),
    .A2(\core_pipeline.pipeline_registers.registers[10][31] ),
    .A3(\core_pipeline.pipeline_registers.registers[11][31] ),
    .S0(net561),
    .S1(net541),
    .X(_05566_));
 sky130_fd_sc_hd__or2_1 _09543_ (.A(net523),
    .B(_05566_),
    .X(_05567_));
 sky130_fd_sc_hd__o211a_1 _09544_ (.A1(net465),
    .A2(_05565_),
    .B1(_05567_),
    .C1(net518),
    .X(_05568_));
 sky130_fd_sc_hd__mux4_1 _09545_ (.A0(\core_pipeline.pipeline_registers.registers[0][31] ),
    .A1(\core_pipeline.pipeline_registers.registers[1][31] ),
    .A2(\core_pipeline.pipeline_registers.registers[2][31] ),
    .A3(\core_pipeline.pipeline_registers.registers[3][31] ),
    .S0(net563),
    .S1(net540),
    .X(_05569_));
 sky130_fd_sc_hd__mux4_1 _09546_ (.A0(\core_pipeline.pipeline_registers.registers[4][31] ),
    .A1(\core_pipeline.pipeline_registers.registers[5][31] ),
    .A2(\core_pipeline.pipeline_registers.registers[6][31] ),
    .A3(\core_pipeline.pipeline_registers.registers[7][31] ),
    .S0(net563),
    .S1(net540),
    .X(_05570_));
 sky130_fd_sc_hd__a221o_1 _09547_ (.A1(_04680_),
    .A2(_05569_),
    .B1(_05570_),
    .B2(_04694_),
    .C1(net512),
    .X(_05571_));
 sky130_fd_sc_hd__mux2_1 _09548_ (.A0(\core_pipeline.pipeline_registers.registers[30][31] ),
    .A1(\core_pipeline.pipeline_registers.registers[31][31] ),
    .S(net561),
    .X(_05572_));
 sky130_fd_sc_hd__a221o_1 _09549_ (.A1(\core_pipeline.pipeline_registers.registers[28][31] ),
    .A2(_04681_),
    .B1(net366),
    .B2(\core_pipeline.pipeline_registers.registers[29][31] ),
    .C1(net465),
    .X(_05573_));
 sky130_fd_sc_hd__a21o_1 _09550_ (.A1(net538),
    .A2(_05572_),
    .B1(_05573_),
    .X(_05574_));
 sky130_fd_sc_hd__mux2_1 _09551_ (.A0(\core_pipeline.pipeline_registers.registers[26][31] ),
    .A1(\core_pipeline.pipeline_registers.registers[27][31] ),
    .S(net562),
    .X(_05575_));
 sky130_fd_sc_hd__a221o_1 _09552_ (.A1(\core_pipeline.pipeline_registers.registers[24][31] ),
    .A2(_04681_),
    .B1(net366),
    .B2(\core_pipeline.pipeline_registers.registers[25][31] ),
    .C1(net523),
    .X(_05576_));
 sky130_fd_sc_hd__a21o_1 _09553_ (.A1(net539),
    .A2(_05575_),
    .B1(_05576_),
    .X(_05577_));
 sky130_fd_sc_hd__and3_1 _09554_ (.A(net518),
    .B(_05574_),
    .C(_05577_),
    .X(_05578_));
 sky130_fd_sc_hd__mux4_1 _09555_ (.A0(\core_pipeline.pipeline_registers.registers[20][31] ),
    .A1(\core_pipeline.pipeline_registers.registers[21][31] ),
    .A2(\core_pipeline.pipeline_registers.registers[22][31] ),
    .A3(\core_pipeline.pipeline_registers.registers[23][31] ),
    .S0(net561),
    .S1(net541),
    .X(_05579_));
 sky130_fd_sc_hd__a31o_1 _09556_ (.A1(\core_pipeline.pipeline_registers.registers[17][31] ),
    .A2(_04680_),
    .A3(_04695_),
    .B1(_03330_),
    .X(_05580_));
 sky130_fd_sc_hd__mux2_1 _09557_ (.A0(\core_pipeline.pipeline_registers.registers[18][31] ),
    .A1(\core_pipeline.pipeline_registers.registers[19][31] ),
    .S(net561),
    .X(_05581_));
 sky130_fd_sc_hd__a22o_1 _09558_ (.A1(\core_pipeline.pipeline_registers.registers[16][31] ),
    .A2(net278),
    .B1(net362),
    .B2(_05581_),
    .X(_05582_));
 sky130_fd_sc_hd__a211o_1 _09559_ (.A1(_04694_),
    .A2(_05579_),
    .B1(_05580_),
    .C1(_05582_),
    .X(_05583_));
 sky130_fd_sc_hd__o22a_2 _09560_ (.A1(_05568_),
    .A2(_05571_),
    .B1(_05578_),
    .B2(_05583_),
    .X(_05584_));
 sky130_fd_sc_hd__mux2_1 _09561_ (.A0(\core_pipeline.decode_to_execute_rs2_data[31] ),
    .A1(_05584_),
    .S(net147),
    .X(_00563_));
 sky130_fd_sc_hd__nor2_8 _09562_ (.A(_04469_),
    .B(_04934_),
    .Y(_05585_));
 sky130_fd_sc_hd__mux2_1 _09563_ (.A0(\core_pipeline.pipeline_registers.registers[30][0] ),
    .A1(net349),
    .S(net213),
    .X(_00564_));
 sky130_fd_sc_hd__mux2_1 _09564_ (.A0(\core_pipeline.pipeline_registers.registers[30][1] ),
    .A1(net346),
    .S(net214),
    .X(_00565_));
 sky130_fd_sc_hd__mux2_1 _09565_ (.A0(\core_pipeline.pipeline_registers.registers[30][2] ),
    .A1(net344),
    .S(net214),
    .X(_00566_));
 sky130_fd_sc_hd__mux2_1 _09566_ (.A0(\core_pipeline.pipeline_registers.registers[30][3] ),
    .A1(net342),
    .S(net213),
    .X(_00567_));
 sky130_fd_sc_hd__mux2_1 _09567_ (.A0(\core_pipeline.pipeline_registers.registers[30][4] ),
    .A1(net341),
    .S(net213),
    .X(_00568_));
 sky130_fd_sc_hd__mux2_1 _09568_ (.A0(\core_pipeline.pipeline_registers.registers[30][5] ),
    .A1(net338),
    .S(net214),
    .X(_00569_));
 sky130_fd_sc_hd__mux2_1 _09569_ (.A0(\core_pipeline.pipeline_registers.registers[30][6] ),
    .A1(net336),
    .S(net214),
    .X(_00570_));
 sky130_fd_sc_hd__mux2_1 _09570_ (.A0(\core_pipeline.pipeline_registers.registers[30][7] ),
    .A1(net333),
    .S(net213),
    .X(_00571_));
 sky130_fd_sc_hd__mux2_1 _09571_ (.A0(\core_pipeline.pipeline_registers.registers[30][8] ),
    .A1(net331),
    .S(net213),
    .X(_00572_));
 sky130_fd_sc_hd__mux2_1 _09572_ (.A0(\core_pipeline.pipeline_registers.registers[30][9] ),
    .A1(net330),
    .S(net213),
    .X(_00573_));
 sky130_fd_sc_hd__mux2_1 _09573_ (.A0(\core_pipeline.pipeline_registers.registers[30][10] ),
    .A1(net328),
    .S(net213),
    .X(_00574_));
 sky130_fd_sc_hd__mux2_1 _09574_ (.A0(\core_pipeline.pipeline_registers.registers[30][11] ),
    .A1(net326),
    .S(net213),
    .X(_00575_));
 sky130_fd_sc_hd__mux2_1 _09575_ (.A0(\core_pipeline.pipeline_registers.registers[30][12] ),
    .A1(net324),
    .S(net213),
    .X(_00576_));
 sky130_fd_sc_hd__mux2_1 _09576_ (.A0(\core_pipeline.pipeline_registers.registers[30][13] ),
    .A1(net322),
    .S(net213),
    .X(_00577_));
 sky130_fd_sc_hd__mux2_1 _09577_ (.A0(\core_pipeline.pipeline_registers.registers[30][14] ),
    .A1(net319),
    .S(net213),
    .X(_00578_));
 sky130_fd_sc_hd__mux2_1 _09578_ (.A0(\core_pipeline.pipeline_registers.registers[30][15] ),
    .A1(net318),
    .S(net213),
    .X(_00579_));
 sky130_fd_sc_hd__mux2_1 _09579_ (.A0(\core_pipeline.pipeline_registers.registers[30][16] ),
    .A1(net316),
    .S(net213),
    .X(_00580_));
 sky130_fd_sc_hd__mux2_1 _09580_ (.A0(\core_pipeline.pipeline_registers.registers[30][17] ),
    .A1(net312),
    .S(net214),
    .X(_00581_));
 sky130_fd_sc_hd__mux2_1 _09581_ (.A0(\core_pipeline.pipeline_registers.registers[30][18] ),
    .A1(net310),
    .S(net214),
    .X(_00582_));
 sky130_fd_sc_hd__mux2_1 _09582_ (.A0(\core_pipeline.pipeline_registers.registers[30][19] ),
    .A1(net309),
    .S(net214),
    .X(_00583_));
 sky130_fd_sc_hd__mux2_1 _09583_ (.A0(\core_pipeline.pipeline_registers.registers[30][20] ),
    .A1(net305),
    .S(net214),
    .X(_00584_));
 sky130_fd_sc_hd__mux2_1 _09584_ (.A0(\core_pipeline.pipeline_registers.registers[30][21] ),
    .A1(net303),
    .S(net214),
    .X(_00585_));
 sky130_fd_sc_hd__mux2_1 _09585_ (.A0(\core_pipeline.pipeline_registers.registers[30][22] ),
    .A1(net302),
    .S(net213),
    .X(_00586_));
 sky130_fd_sc_hd__mux2_1 _09586_ (.A0(\core_pipeline.pipeline_registers.registers[30][23] ),
    .A1(net299),
    .S(net214),
    .X(_00587_));
 sky130_fd_sc_hd__mux2_1 _09587_ (.A0(\core_pipeline.pipeline_registers.registers[30][24] ),
    .A1(net298),
    .S(net213),
    .X(_00588_));
 sky130_fd_sc_hd__mux2_1 _09588_ (.A0(\core_pipeline.pipeline_registers.registers[30][25] ),
    .A1(net296),
    .S(net213),
    .X(_00589_));
 sky130_fd_sc_hd__mux2_1 _09589_ (.A0(\core_pipeline.pipeline_registers.registers[30][26] ),
    .A1(net294),
    .S(net213),
    .X(_00590_));
 sky130_fd_sc_hd__mux2_1 _09590_ (.A0(\core_pipeline.pipeline_registers.registers[30][27] ),
    .A1(net291),
    .S(net214),
    .X(_00591_));
 sky130_fd_sc_hd__mux2_1 _09591_ (.A0(\core_pipeline.pipeline_registers.registers[30][28] ),
    .A1(net289),
    .S(net214),
    .X(_00592_));
 sky130_fd_sc_hd__mux2_1 _09592_ (.A0(\core_pipeline.pipeline_registers.registers[30][29] ),
    .A1(net286),
    .S(net214),
    .X(_00593_));
 sky130_fd_sc_hd__mux2_1 _09593_ (.A0(\core_pipeline.pipeline_registers.registers[30][30] ),
    .A1(net284),
    .S(net214),
    .X(_00594_));
 sky130_fd_sc_hd__mux2_1 _09594_ (.A0(\core_pipeline.pipeline_registers.registers[30][31] ),
    .A1(net282),
    .S(net214),
    .X(_00595_));
 sky130_fd_sc_hd__or3b_4 _09595_ (.A(_04468_),
    .B(\core_pipeline.memory_to_writeback_rd_address[2] ),
    .C_N(\core_pipeline.memory_to_writeback_rd_address[4] ),
    .X(_05586_));
 sky130_fd_sc_hd__nor2_8 _09596_ (.A(_03915_),
    .B(_05586_),
    .Y(_05587_));
 sky130_fd_sc_hd__mux2_1 _09597_ (.A0(\core_pipeline.pipeline_registers.registers[27][0] ),
    .A1(net349),
    .S(net211),
    .X(_00596_));
 sky130_fd_sc_hd__mux2_1 _09598_ (.A0(\core_pipeline.pipeline_registers.registers[27][1] ),
    .A1(net346),
    .S(net212),
    .X(_00597_));
 sky130_fd_sc_hd__mux2_1 _09599_ (.A0(\core_pipeline.pipeline_registers.registers[27][2] ),
    .A1(net344),
    .S(net212),
    .X(_00598_));
 sky130_fd_sc_hd__mux2_1 _09600_ (.A0(\core_pipeline.pipeline_registers.registers[27][3] ),
    .A1(net342),
    .S(net211),
    .X(_00599_));
 sky130_fd_sc_hd__mux2_1 _09601_ (.A0(\core_pipeline.pipeline_registers.registers[27][4] ),
    .A1(net341),
    .S(net211),
    .X(_00600_));
 sky130_fd_sc_hd__mux2_1 _09602_ (.A0(\core_pipeline.pipeline_registers.registers[27][5] ),
    .A1(net337),
    .S(net212),
    .X(_00601_));
 sky130_fd_sc_hd__mux2_1 _09603_ (.A0(\core_pipeline.pipeline_registers.registers[27][6] ),
    .A1(net336),
    .S(net212),
    .X(_00602_));
 sky130_fd_sc_hd__mux2_1 _09604_ (.A0(\core_pipeline.pipeline_registers.registers[27][7] ),
    .A1(net333),
    .S(net211),
    .X(_00603_));
 sky130_fd_sc_hd__mux2_1 _09605_ (.A0(\core_pipeline.pipeline_registers.registers[27][8] ),
    .A1(net331),
    .S(net211),
    .X(_00604_));
 sky130_fd_sc_hd__mux2_1 _09606_ (.A0(\core_pipeline.pipeline_registers.registers[27][9] ),
    .A1(net330),
    .S(net211),
    .X(_00605_));
 sky130_fd_sc_hd__mux2_1 _09607_ (.A0(\core_pipeline.pipeline_registers.registers[27][10] ),
    .A1(net328),
    .S(net211),
    .X(_00606_));
 sky130_fd_sc_hd__mux2_1 _09608_ (.A0(\core_pipeline.pipeline_registers.registers[27][11] ),
    .A1(net326),
    .S(net211),
    .X(_00607_));
 sky130_fd_sc_hd__mux2_1 _09609_ (.A0(\core_pipeline.pipeline_registers.registers[27][12] ),
    .A1(net324),
    .S(net211),
    .X(_00608_));
 sky130_fd_sc_hd__mux2_1 _09610_ (.A0(\core_pipeline.pipeline_registers.registers[27][13] ),
    .A1(net322),
    .S(net211),
    .X(_00609_));
 sky130_fd_sc_hd__mux2_1 _09611_ (.A0(\core_pipeline.pipeline_registers.registers[27][14] ),
    .A1(net319),
    .S(net211),
    .X(_00610_));
 sky130_fd_sc_hd__mux2_1 _09612_ (.A0(\core_pipeline.pipeline_registers.registers[27][15] ),
    .A1(net318),
    .S(net211),
    .X(_00611_));
 sky130_fd_sc_hd__mux2_1 _09613_ (.A0(\core_pipeline.pipeline_registers.registers[27][16] ),
    .A1(net316),
    .S(net211),
    .X(_00612_));
 sky130_fd_sc_hd__mux2_1 _09614_ (.A0(\core_pipeline.pipeline_registers.registers[27][17] ),
    .A1(net312),
    .S(net212),
    .X(_00613_));
 sky130_fd_sc_hd__mux2_1 _09615_ (.A0(\core_pipeline.pipeline_registers.registers[27][18] ),
    .A1(net310),
    .S(net212),
    .X(_00614_));
 sky130_fd_sc_hd__mux2_1 _09616_ (.A0(\core_pipeline.pipeline_registers.registers[27][19] ),
    .A1(net308),
    .S(net212),
    .X(_00615_));
 sky130_fd_sc_hd__mux2_1 _09617_ (.A0(\core_pipeline.pipeline_registers.registers[27][20] ),
    .A1(net307),
    .S(net212),
    .X(_00616_));
 sky130_fd_sc_hd__mux2_1 _09618_ (.A0(\core_pipeline.pipeline_registers.registers[27][21] ),
    .A1(net304),
    .S(net212),
    .X(_00617_));
 sky130_fd_sc_hd__mux2_1 _09619_ (.A0(\core_pipeline.pipeline_registers.registers[27][22] ),
    .A1(net301),
    .S(net212),
    .X(_00618_));
 sky130_fd_sc_hd__mux2_1 _09620_ (.A0(\core_pipeline.pipeline_registers.registers[27][23] ),
    .A1(net300),
    .S(net212),
    .X(_00619_));
 sky130_fd_sc_hd__mux2_1 _09621_ (.A0(\core_pipeline.pipeline_registers.registers[27][24] ),
    .A1(net297),
    .S(net211),
    .X(_00620_));
 sky130_fd_sc_hd__mux2_1 _09622_ (.A0(\core_pipeline.pipeline_registers.registers[27][25] ),
    .A1(net296),
    .S(net211),
    .X(_00621_));
 sky130_fd_sc_hd__mux2_1 _09623_ (.A0(\core_pipeline.pipeline_registers.registers[27][26] ),
    .A1(net294),
    .S(net211),
    .X(_00622_));
 sky130_fd_sc_hd__mux2_1 _09624_ (.A0(\core_pipeline.pipeline_registers.registers[27][27] ),
    .A1(net291),
    .S(net212),
    .X(_00623_));
 sky130_fd_sc_hd__mux2_1 _09625_ (.A0(\core_pipeline.pipeline_registers.registers[27][28] ),
    .A1(net290),
    .S(net212),
    .X(_00624_));
 sky130_fd_sc_hd__mux2_1 _09626_ (.A0(\core_pipeline.pipeline_registers.registers[27][29] ),
    .A1(net286),
    .S(net212),
    .X(_00625_));
 sky130_fd_sc_hd__mux2_1 _09627_ (.A0(\core_pipeline.pipeline_registers.registers[27][30] ),
    .A1(net284),
    .S(net211),
    .X(_00626_));
 sky130_fd_sc_hd__mux2_1 _09628_ (.A0(\core_pipeline.pipeline_registers.registers[27][31] ),
    .A1(net283),
    .S(net212),
    .X(_00627_));
 sky130_fd_sc_hd__nor2_8 _09629_ (.A(_04934_),
    .B(_05586_),
    .Y(_05588_));
 sky130_fd_sc_hd__mux2_1 _09630_ (.A0(\core_pipeline.pipeline_registers.registers[26][0] ),
    .A1(net349),
    .S(net209),
    .X(_00628_));
 sky130_fd_sc_hd__mux2_1 _09631_ (.A0(\core_pipeline.pipeline_registers.registers[26][1] ),
    .A1(net346),
    .S(net210),
    .X(_00629_));
 sky130_fd_sc_hd__mux2_1 _09632_ (.A0(\core_pipeline.pipeline_registers.registers[26][2] ),
    .A1(net344),
    .S(net210),
    .X(_00630_));
 sky130_fd_sc_hd__mux2_1 _09633_ (.A0(\core_pipeline.pipeline_registers.registers[26][3] ),
    .A1(net342),
    .S(net209),
    .X(_00631_));
 sky130_fd_sc_hd__mux2_1 _09634_ (.A0(\core_pipeline.pipeline_registers.registers[26][4] ),
    .A1(net341),
    .S(net209),
    .X(_00632_));
 sky130_fd_sc_hd__mux2_1 _09635_ (.A0(\core_pipeline.pipeline_registers.registers[26][5] ),
    .A1(net337),
    .S(net210),
    .X(_00633_));
 sky130_fd_sc_hd__mux2_1 _09636_ (.A0(\core_pipeline.pipeline_registers.registers[26][6] ),
    .A1(net336),
    .S(net210),
    .X(_00634_));
 sky130_fd_sc_hd__mux2_1 _09637_ (.A0(\core_pipeline.pipeline_registers.registers[26][7] ),
    .A1(net333),
    .S(net209),
    .X(_00635_));
 sky130_fd_sc_hd__mux2_1 _09638_ (.A0(\core_pipeline.pipeline_registers.registers[26][8] ),
    .A1(net331),
    .S(net209),
    .X(_00636_));
 sky130_fd_sc_hd__mux2_1 _09639_ (.A0(\core_pipeline.pipeline_registers.registers[26][9] ),
    .A1(net330),
    .S(net209),
    .X(_00637_));
 sky130_fd_sc_hd__mux2_1 _09640_ (.A0(\core_pipeline.pipeline_registers.registers[26][10] ),
    .A1(net328),
    .S(net209),
    .X(_00638_));
 sky130_fd_sc_hd__mux2_1 _09641_ (.A0(\core_pipeline.pipeline_registers.registers[26][11] ),
    .A1(net326),
    .S(net209),
    .X(_00639_));
 sky130_fd_sc_hd__mux2_1 _09642_ (.A0(\core_pipeline.pipeline_registers.registers[26][12] ),
    .A1(net324),
    .S(net209),
    .X(_00640_));
 sky130_fd_sc_hd__mux2_1 _09643_ (.A0(\core_pipeline.pipeline_registers.registers[26][13] ),
    .A1(net322),
    .S(net209),
    .X(_00641_));
 sky130_fd_sc_hd__mux2_1 _09644_ (.A0(\core_pipeline.pipeline_registers.registers[26][14] ),
    .A1(net319),
    .S(net209),
    .X(_00642_));
 sky130_fd_sc_hd__mux2_1 _09645_ (.A0(\core_pipeline.pipeline_registers.registers[26][15] ),
    .A1(net318),
    .S(net209),
    .X(_00643_));
 sky130_fd_sc_hd__mux2_1 _09646_ (.A0(\core_pipeline.pipeline_registers.registers[26][16] ),
    .A1(net316),
    .S(net209),
    .X(_00644_));
 sky130_fd_sc_hd__mux2_1 _09647_ (.A0(\core_pipeline.pipeline_registers.registers[26][17] ),
    .A1(net312),
    .S(net210),
    .X(_00645_));
 sky130_fd_sc_hd__mux2_1 _09648_ (.A0(\core_pipeline.pipeline_registers.registers[26][18] ),
    .A1(net310),
    .S(net210),
    .X(_00646_));
 sky130_fd_sc_hd__mux2_1 _09649_ (.A0(\core_pipeline.pipeline_registers.registers[26][19] ),
    .A1(net308),
    .S(net210),
    .X(_00647_));
 sky130_fd_sc_hd__mux2_1 _09650_ (.A0(\core_pipeline.pipeline_registers.registers[26][20] ),
    .A1(net307),
    .S(net210),
    .X(_00648_));
 sky130_fd_sc_hd__mux2_1 _09651_ (.A0(\core_pipeline.pipeline_registers.registers[26][21] ),
    .A1(net304),
    .S(net210),
    .X(_00649_));
 sky130_fd_sc_hd__mux2_1 _09652_ (.A0(\core_pipeline.pipeline_registers.registers[26][22] ),
    .A1(net302),
    .S(net210),
    .X(_00650_));
 sky130_fd_sc_hd__mux2_1 _09653_ (.A0(\core_pipeline.pipeline_registers.registers[26][23] ),
    .A1(net299),
    .S(net210),
    .X(_00651_));
 sky130_fd_sc_hd__mux2_1 _09654_ (.A0(\core_pipeline.pipeline_registers.registers[26][24] ),
    .A1(net297),
    .S(net209),
    .X(_00652_));
 sky130_fd_sc_hd__mux2_1 _09655_ (.A0(\core_pipeline.pipeline_registers.registers[26][25] ),
    .A1(net296),
    .S(net209),
    .X(_00653_));
 sky130_fd_sc_hd__mux2_1 _09656_ (.A0(\core_pipeline.pipeline_registers.registers[26][26] ),
    .A1(net294),
    .S(net209),
    .X(_00654_));
 sky130_fd_sc_hd__mux2_1 _09657_ (.A0(\core_pipeline.pipeline_registers.registers[26][27] ),
    .A1(net291),
    .S(net210),
    .X(_00655_));
 sky130_fd_sc_hd__mux2_1 _09658_ (.A0(\core_pipeline.pipeline_registers.registers[26][28] ),
    .A1(net290),
    .S(net210),
    .X(_00656_));
 sky130_fd_sc_hd__mux2_1 _09659_ (.A0(\core_pipeline.pipeline_registers.registers[26][29] ),
    .A1(net286),
    .S(net210),
    .X(_00657_));
 sky130_fd_sc_hd__mux2_1 _09660_ (.A0(\core_pipeline.pipeline_registers.registers[26][30] ),
    .A1(net284),
    .S(net209),
    .X(_00658_));
 sky130_fd_sc_hd__mux2_1 _09661_ (.A0(\core_pipeline.pipeline_registers.registers[26][31] ),
    .A1(net283),
    .S(net210),
    .X(_00659_));
 sky130_fd_sc_hd__or2_4 _09662_ (.A(\core_pipeline.memory_to_writeback_rd_address[1] ),
    .B(_03913_),
    .X(_05589_));
 sky130_fd_sc_hd__nor2_8 _09663_ (.A(_05586_),
    .B(_05589_),
    .Y(_05590_));
 sky130_fd_sc_hd__mux2_1 _09664_ (.A0(\core_pipeline.pipeline_registers.registers[25][0] ),
    .A1(net349),
    .S(net207),
    .X(_00660_));
 sky130_fd_sc_hd__mux2_1 _09665_ (.A0(\core_pipeline.pipeline_registers.registers[25][1] ),
    .A1(net346),
    .S(net208),
    .X(_00661_));
 sky130_fd_sc_hd__mux2_1 _09666_ (.A0(\core_pipeline.pipeline_registers.registers[25][2] ),
    .A1(net344),
    .S(net208),
    .X(_00662_));
 sky130_fd_sc_hd__mux2_1 _09667_ (.A0(\core_pipeline.pipeline_registers.registers[25][3] ),
    .A1(net342),
    .S(net207),
    .X(_00663_));
 sky130_fd_sc_hd__mux2_1 _09668_ (.A0(\core_pipeline.pipeline_registers.registers[25][4] ),
    .A1(net341),
    .S(net207),
    .X(_00664_));
 sky130_fd_sc_hd__mux2_1 _09669_ (.A0(\core_pipeline.pipeline_registers.registers[25][5] ),
    .A1(net337),
    .S(net208),
    .X(_00665_));
 sky130_fd_sc_hd__mux2_1 _09670_ (.A0(\core_pipeline.pipeline_registers.registers[25][6] ),
    .A1(net336),
    .S(net207),
    .X(_00666_));
 sky130_fd_sc_hd__mux2_1 _09671_ (.A0(\core_pipeline.pipeline_registers.registers[25][7] ),
    .A1(net333),
    .S(net207),
    .X(_00667_));
 sky130_fd_sc_hd__mux2_1 _09672_ (.A0(\core_pipeline.pipeline_registers.registers[25][8] ),
    .A1(net331),
    .S(net207),
    .X(_00668_));
 sky130_fd_sc_hd__mux2_1 _09673_ (.A0(\core_pipeline.pipeline_registers.registers[25][9] ),
    .A1(net330),
    .S(net207),
    .X(_00669_));
 sky130_fd_sc_hd__mux2_1 _09674_ (.A0(\core_pipeline.pipeline_registers.registers[25][10] ),
    .A1(net328),
    .S(net207),
    .X(_00670_));
 sky130_fd_sc_hd__mux2_1 _09675_ (.A0(\core_pipeline.pipeline_registers.registers[25][11] ),
    .A1(net326),
    .S(net207),
    .X(_00671_));
 sky130_fd_sc_hd__mux2_1 _09676_ (.A0(\core_pipeline.pipeline_registers.registers[25][12] ),
    .A1(net324),
    .S(net207),
    .X(_00672_));
 sky130_fd_sc_hd__mux2_1 _09677_ (.A0(\core_pipeline.pipeline_registers.registers[25][13] ),
    .A1(net322),
    .S(net207),
    .X(_00673_));
 sky130_fd_sc_hd__mux2_1 _09678_ (.A0(\core_pipeline.pipeline_registers.registers[25][14] ),
    .A1(net319),
    .S(net207),
    .X(_00674_));
 sky130_fd_sc_hd__mux2_1 _09679_ (.A0(\core_pipeline.pipeline_registers.registers[25][15] ),
    .A1(net318),
    .S(net207),
    .X(_00675_));
 sky130_fd_sc_hd__mux2_1 _09680_ (.A0(\core_pipeline.pipeline_registers.registers[25][16] ),
    .A1(net316),
    .S(net207),
    .X(_00676_));
 sky130_fd_sc_hd__mux2_1 _09681_ (.A0(\core_pipeline.pipeline_registers.registers[25][17] ),
    .A1(net312),
    .S(net208),
    .X(_00677_));
 sky130_fd_sc_hd__mux2_1 _09682_ (.A0(\core_pipeline.pipeline_registers.registers[25][18] ),
    .A1(net310),
    .S(net208),
    .X(_00678_));
 sky130_fd_sc_hd__mux2_1 _09683_ (.A0(\core_pipeline.pipeline_registers.registers[25][19] ),
    .A1(net308),
    .S(net208),
    .X(_00679_));
 sky130_fd_sc_hd__mux2_1 _09684_ (.A0(\core_pipeline.pipeline_registers.registers[25][20] ),
    .A1(net307),
    .S(net208),
    .X(_00680_));
 sky130_fd_sc_hd__mux2_1 _09685_ (.A0(\core_pipeline.pipeline_registers.registers[25][21] ),
    .A1(net304),
    .S(net208),
    .X(_00681_));
 sky130_fd_sc_hd__mux2_1 _09686_ (.A0(\core_pipeline.pipeline_registers.registers[25][22] ),
    .A1(net302),
    .S(net208),
    .X(_00682_));
 sky130_fd_sc_hd__mux2_1 _09687_ (.A0(\core_pipeline.pipeline_registers.registers[25][23] ),
    .A1(net299),
    .S(net208),
    .X(_00683_));
 sky130_fd_sc_hd__mux2_1 _09688_ (.A0(\core_pipeline.pipeline_registers.registers[25][24] ),
    .A1(net298),
    .S(net207),
    .X(_00684_));
 sky130_fd_sc_hd__mux2_1 _09689_ (.A0(\core_pipeline.pipeline_registers.registers[25][25] ),
    .A1(net296),
    .S(net207),
    .X(_00685_));
 sky130_fd_sc_hd__mux2_1 _09690_ (.A0(\core_pipeline.pipeline_registers.registers[25][26] ),
    .A1(net294),
    .S(net207),
    .X(_00686_));
 sky130_fd_sc_hd__mux2_1 _09691_ (.A0(\core_pipeline.pipeline_registers.registers[25][27] ),
    .A1(net291),
    .S(net208),
    .X(_00687_));
 sky130_fd_sc_hd__mux2_1 _09692_ (.A0(\core_pipeline.pipeline_registers.registers[25][28] ),
    .A1(net290),
    .S(net208),
    .X(_00688_));
 sky130_fd_sc_hd__mux2_1 _09693_ (.A0(\core_pipeline.pipeline_registers.registers[25][29] ),
    .A1(net286),
    .S(net208),
    .X(_00689_));
 sky130_fd_sc_hd__mux2_1 _09694_ (.A0(\core_pipeline.pipeline_registers.registers[25][30] ),
    .A1(net284),
    .S(net208),
    .X(_00690_));
 sky130_fd_sc_hd__mux2_1 _09695_ (.A0(\core_pipeline.pipeline_registers.registers[25][31] ),
    .A1(net283),
    .S(net208),
    .X(_00691_));
 sky130_fd_sc_hd__or2_4 _09696_ (.A(_04939_),
    .B(_05586_),
    .X(_05591_));
 sky130_fd_sc_hd__mux2_1 _09697_ (.A0(net349),
    .A1(\core_pipeline.pipeline_registers.registers[24][0] ),
    .S(net205),
    .X(_00692_));
 sky130_fd_sc_hd__mux2_1 _09698_ (.A0(net346),
    .A1(\core_pipeline.pipeline_registers.registers[24][1] ),
    .S(net206),
    .X(_00693_));
 sky130_fd_sc_hd__mux2_1 _09699_ (.A0(net344),
    .A1(\core_pipeline.pipeline_registers.registers[24][2] ),
    .S(net206),
    .X(_00694_));
 sky130_fd_sc_hd__mux2_1 _09700_ (.A0(net342),
    .A1(\core_pipeline.pipeline_registers.registers[24][3] ),
    .S(net205),
    .X(_00695_));
 sky130_fd_sc_hd__mux2_1 _09701_ (.A0(net341),
    .A1(\core_pipeline.pipeline_registers.registers[24][4] ),
    .S(net205),
    .X(_00696_));
 sky130_fd_sc_hd__mux2_1 _09702_ (.A0(net337),
    .A1(\core_pipeline.pipeline_registers.registers[24][5] ),
    .S(net206),
    .X(_00697_));
 sky130_fd_sc_hd__mux2_1 _09703_ (.A0(net336),
    .A1(\core_pipeline.pipeline_registers.registers[24][6] ),
    .S(net205),
    .X(_00698_));
 sky130_fd_sc_hd__mux2_1 _09704_ (.A0(net333),
    .A1(\core_pipeline.pipeline_registers.registers[24][7] ),
    .S(net205),
    .X(_00699_));
 sky130_fd_sc_hd__mux2_1 _09705_ (.A0(net331),
    .A1(\core_pipeline.pipeline_registers.registers[24][8] ),
    .S(net205),
    .X(_00700_));
 sky130_fd_sc_hd__mux2_1 _09706_ (.A0(net330),
    .A1(\core_pipeline.pipeline_registers.registers[24][9] ),
    .S(net205),
    .X(_00701_));
 sky130_fd_sc_hd__mux2_1 _09707_ (.A0(net328),
    .A1(\core_pipeline.pipeline_registers.registers[24][10] ),
    .S(net205),
    .X(_00702_));
 sky130_fd_sc_hd__mux2_1 _09708_ (.A0(net326),
    .A1(\core_pipeline.pipeline_registers.registers[24][11] ),
    .S(net205),
    .X(_00703_));
 sky130_fd_sc_hd__mux2_1 _09709_ (.A0(net324),
    .A1(\core_pipeline.pipeline_registers.registers[24][12] ),
    .S(net205),
    .X(_00704_));
 sky130_fd_sc_hd__mux2_1 _09710_ (.A0(net322),
    .A1(\core_pipeline.pipeline_registers.registers[24][13] ),
    .S(net205),
    .X(_00705_));
 sky130_fd_sc_hd__mux2_1 _09711_ (.A0(net319),
    .A1(\core_pipeline.pipeline_registers.registers[24][14] ),
    .S(net205),
    .X(_00706_));
 sky130_fd_sc_hd__mux2_1 _09712_ (.A0(net318),
    .A1(\core_pipeline.pipeline_registers.registers[24][15] ),
    .S(net205),
    .X(_00707_));
 sky130_fd_sc_hd__mux2_1 _09713_ (.A0(net316),
    .A1(\core_pipeline.pipeline_registers.registers[24][16] ),
    .S(net205),
    .X(_00708_));
 sky130_fd_sc_hd__mux2_1 _09714_ (.A0(net312),
    .A1(\core_pipeline.pipeline_registers.registers[24][17] ),
    .S(net206),
    .X(_00709_));
 sky130_fd_sc_hd__mux2_1 _09715_ (.A0(net310),
    .A1(\core_pipeline.pipeline_registers.registers[24][18] ),
    .S(net206),
    .X(_00710_));
 sky130_fd_sc_hd__mux2_1 _09716_ (.A0(net308),
    .A1(\core_pipeline.pipeline_registers.registers[24][19] ),
    .S(net206),
    .X(_00711_));
 sky130_fd_sc_hd__mux2_1 _09717_ (.A0(net307),
    .A1(\core_pipeline.pipeline_registers.registers[24][20] ),
    .S(net206),
    .X(_00712_));
 sky130_fd_sc_hd__mux2_1 _09718_ (.A0(net304),
    .A1(\core_pipeline.pipeline_registers.registers[24][21] ),
    .S(net206),
    .X(_00713_));
 sky130_fd_sc_hd__mux2_1 _09719_ (.A0(net302),
    .A1(\core_pipeline.pipeline_registers.registers[24][22] ),
    .S(net206),
    .X(_00714_));
 sky130_fd_sc_hd__mux2_1 _09720_ (.A0(net299),
    .A1(\core_pipeline.pipeline_registers.registers[24][23] ),
    .S(net206),
    .X(_00715_));
 sky130_fd_sc_hd__mux2_1 _09721_ (.A0(net298),
    .A1(\core_pipeline.pipeline_registers.registers[24][24] ),
    .S(net205),
    .X(_00716_));
 sky130_fd_sc_hd__mux2_1 _09722_ (.A0(net296),
    .A1(\core_pipeline.pipeline_registers.registers[24][25] ),
    .S(net205),
    .X(_00717_));
 sky130_fd_sc_hd__mux2_1 _09723_ (.A0(net294),
    .A1(\core_pipeline.pipeline_registers.registers[24][26] ),
    .S(net205),
    .X(_00718_));
 sky130_fd_sc_hd__mux2_1 _09724_ (.A0(net291),
    .A1(\core_pipeline.pipeline_registers.registers[24][27] ),
    .S(net206),
    .X(_00719_));
 sky130_fd_sc_hd__mux2_1 _09725_ (.A0(net290),
    .A1(\core_pipeline.pipeline_registers.registers[24][28] ),
    .S(net206),
    .X(_00720_));
 sky130_fd_sc_hd__mux2_1 _09726_ (.A0(net286),
    .A1(\core_pipeline.pipeline_registers.registers[24][29] ),
    .S(net206),
    .X(_00721_));
 sky130_fd_sc_hd__mux2_1 _09727_ (.A0(net284),
    .A1(\core_pipeline.pipeline_registers.registers[24][30] ),
    .S(net206),
    .X(_00722_));
 sky130_fd_sc_hd__mux2_1 _09728_ (.A0(net283),
    .A1(\core_pipeline.pipeline_registers.registers[24][31] ),
    .S(net206),
    .X(_00723_));
 sky130_fd_sc_hd__or3b_4 _09729_ (.A(\core_pipeline.memory_to_writeback_rd_address[3] ),
    .B(_03912_),
    .C_N(\core_pipeline.memory_to_writeback_rd_address[2] ),
    .X(_05592_));
 sky130_fd_sc_hd__nor2_8 _09730_ (.A(_03915_),
    .B(_05592_),
    .Y(_05593_));
 sky130_fd_sc_hd__mux2_1 _09731_ (.A0(\core_pipeline.pipeline_registers.registers[23][0] ),
    .A1(net349),
    .S(net203),
    .X(_00724_));
 sky130_fd_sc_hd__mux2_1 _09732_ (.A0(\core_pipeline.pipeline_registers.registers[23][1] ),
    .A1(net347),
    .S(net204),
    .X(_00725_));
 sky130_fd_sc_hd__mux2_1 _09733_ (.A0(\core_pipeline.pipeline_registers.registers[23][2] ),
    .A1(net345),
    .S(net204),
    .X(_00726_));
 sky130_fd_sc_hd__mux2_1 _09734_ (.A0(\core_pipeline.pipeline_registers.registers[23][3] ),
    .A1(net342),
    .S(net203),
    .X(_00727_));
 sky130_fd_sc_hd__mux2_1 _09735_ (.A0(\core_pipeline.pipeline_registers.registers[23][4] ),
    .A1(net340),
    .S(net203),
    .X(_00728_));
 sky130_fd_sc_hd__mux2_1 _09736_ (.A0(\core_pipeline.pipeline_registers.registers[23][5] ),
    .A1(net339),
    .S(net204),
    .X(_00729_));
 sky130_fd_sc_hd__mux2_1 _09737_ (.A0(\core_pipeline.pipeline_registers.registers[23][6] ),
    .A1(net336),
    .S(net203),
    .X(_00730_));
 sky130_fd_sc_hd__mux2_1 _09738_ (.A0(\core_pipeline.pipeline_registers.registers[23][7] ),
    .A1(net333),
    .S(net203),
    .X(_00731_));
 sky130_fd_sc_hd__mux2_1 _09739_ (.A0(\core_pipeline.pipeline_registers.registers[23][8] ),
    .A1(net331),
    .S(net203),
    .X(_00732_));
 sky130_fd_sc_hd__mux2_1 _09740_ (.A0(\core_pipeline.pipeline_registers.registers[23][9] ),
    .A1(net329),
    .S(net203),
    .X(_00733_));
 sky130_fd_sc_hd__mux2_1 _09741_ (.A0(\core_pipeline.pipeline_registers.registers[23][10] ),
    .A1(net327),
    .S(net203),
    .X(_00734_));
 sky130_fd_sc_hd__mux2_1 _09742_ (.A0(\core_pipeline.pipeline_registers.registers[23][11] ),
    .A1(net326),
    .S(net203),
    .X(_00735_));
 sky130_fd_sc_hd__mux2_1 _09743_ (.A0(\core_pipeline.pipeline_registers.registers[23][12] ),
    .A1(net323),
    .S(net203),
    .X(_00736_));
 sky130_fd_sc_hd__mux2_1 _09744_ (.A0(\core_pipeline.pipeline_registers.registers[23][13] ),
    .A1(net321),
    .S(net203),
    .X(_00737_));
 sky130_fd_sc_hd__mux2_1 _09745_ (.A0(\core_pipeline.pipeline_registers.registers[23][14] ),
    .A1(net319),
    .S(net203),
    .X(_00738_));
 sky130_fd_sc_hd__mux2_1 _09746_ (.A0(\core_pipeline.pipeline_registers.registers[23][15] ),
    .A1(net317),
    .S(net203),
    .X(_00739_));
 sky130_fd_sc_hd__mux2_1 _09747_ (.A0(\core_pipeline.pipeline_registers.registers[23][16] ),
    .A1(net316),
    .S(net203),
    .X(_00740_));
 sky130_fd_sc_hd__mux2_1 _09748_ (.A0(\core_pipeline.pipeline_registers.registers[23][17] ),
    .A1(net314),
    .S(net204),
    .X(_00741_));
 sky130_fd_sc_hd__mux2_1 _09749_ (.A0(\core_pipeline.pipeline_registers.registers[23][18] ),
    .A1(net310),
    .S(net204),
    .X(_00742_));
 sky130_fd_sc_hd__mux2_1 _09750_ (.A0(\core_pipeline.pipeline_registers.registers[23][19] ),
    .A1(net309),
    .S(net204),
    .X(_00743_));
 sky130_fd_sc_hd__mux2_1 _09751_ (.A0(\core_pipeline.pipeline_registers.registers[23][20] ),
    .A1(net307),
    .S(net204),
    .X(_00744_));
 sky130_fd_sc_hd__mux2_1 _09752_ (.A0(\core_pipeline.pipeline_registers.registers[23][21] ),
    .A1(net304),
    .S(net204),
    .X(_00745_));
 sky130_fd_sc_hd__mux2_1 _09753_ (.A0(\core_pipeline.pipeline_registers.registers[23][22] ),
    .A1(net302),
    .S(net204),
    .X(_00746_));
 sky130_fd_sc_hd__mux2_1 _09754_ (.A0(\core_pipeline.pipeline_registers.registers[23][23] ),
    .A1(net299),
    .S(net204),
    .X(_00747_));
 sky130_fd_sc_hd__mux2_1 _09755_ (.A0(\core_pipeline.pipeline_registers.registers[23][24] ),
    .A1(net297),
    .S(net203),
    .X(_00748_));
 sky130_fd_sc_hd__mux2_1 _09756_ (.A0(\core_pipeline.pipeline_registers.registers[23][25] ),
    .A1(net295),
    .S(net203),
    .X(_00749_));
 sky130_fd_sc_hd__mux2_1 _09757_ (.A0(\core_pipeline.pipeline_registers.registers[23][26] ),
    .A1(net293),
    .S(net203),
    .X(_00750_));
 sky130_fd_sc_hd__mux2_1 _09758_ (.A0(\core_pipeline.pipeline_registers.registers[23][27] ),
    .A1(net291),
    .S(net204),
    .X(_00751_));
 sky130_fd_sc_hd__mux2_1 _09759_ (.A0(\core_pipeline.pipeline_registers.registers[23][28] ),
    .A1(net290),
    .S(net204),
    .X(_00752_));
 sky130_fd_sc_hd__mux2_1 _09760_ (.A0(\core_pipeline.pipeline_registers.registers[23][29] ),
    .A1(net287),
    .S(net204),
    .X(_00753_));
 sky130_fd_sc_hd__mux2_1 _09761_ (.A0(\core_pipeline.pipeline_registers.registers[23][30] ),
    .A1(net285),
    .S(net204),
    .X(_00754_));
 sky130_fd_sc_hd__mux2_1 _09762_ (.A0(\core_pipeline.pipeline_registers.registers[23][31] ),
    .A1(net283),
    .S(net204),
    .X(_00755_));
 sky130_fd_sc_hd__nor2_8 _09763_ (.A(_05589_),
    .B(_05592_),
    .Y(_05594_));
 sky130_fd_sc_hd__mux2_1 _09764_ (.A0(\core_pipeline.pipeline_registers.registers[21][0] ),
    .A1(net349),
    .S(net201),
    .X(_00756_));
 sky130_fd_sc_hd__mux2_1 _09765_ (.A0(\core_pipeline.pipeline_registers.registers[21][1] ),
    .A1(net347),
    .S(net202),
    .X(_00757_));
 sky130_fd_sc_hd__mux2_1 _09766_ (.A0(\core_pipeline.pipeline_registers.registers[21][2] ),
    .A1(net345),
    .S(net202),
    .X(_00758_));
 sky130_fd_sc_hd__mux2_1 _09767_ (.A0(\core_pipeline.pipeline_registers.registers[21][3] ),
    .A1(net342),
    .S(net201),
    .X(_00759_));
 sky130_fd_sc_hd__mux2_1 _09768_ (.A0(\core_pipeline.pipeline_registers.registers[21][4] ),
    .A1(net341),
    .S(net201),
    .X(_00760_));
 sky130_fd_sc_hd__mux2_1 _09769_ (.A0(\core_pipeline.pipeline_registers.registers[21][5] ),
    .A1(net338),
    .S(net202),
    .X(_00761_));
 sky130_fd_sc_hd__mux2_1 _09770_ (.A0(\core_pipeline.pipeline_registers.registers[21][6] ),
    .A1(net336),
    .S(net201),
    .X(_00762_));
 sky130_fd_sc_hd__mux2_1 _09771_ (.A0(\core_pipeline.pipeline_registers.registers[21][7] ),
    .A1(net333),
    .S(net201),
    .X(_00763_));
 sky130_fd_sc_hd__mux2_1 _09772_ (.A0(\core_pipeline.pipeline_registers.registers[21][8] ),
    .A1(net331),
    .S(net201),
    .X(_00764_));
 sky130_fd_sc_hd__mux2_1 _09773_ (.A0(\core_pipeline.pipeline_registers.registers[21][9] ),
    .A1(net330),
    .S(net201),
    .X(_00765_));
 sky130_fd_sc_hd__mux2_1 _09774_ (.A0(\core_pipeline.pipeline_registers.registers[21][10] ),
    .A1(net327),
    .S(net201),
    .X(_00766_));
 sky130_fd_sc_hd__mux2_1 _09775_ (.A0(\core_pipeline.pipeline_registers.registers[21][11] ),
    .A1(net326),
    .S(net201),
    .X(_00767_));
 sky130_fd_sc_hd__mux2_1 _09776_ (.A0(\core_pipeline.pipeline_registers.registers[21][12] ),
    .A1(net324),
    .S(net201),
    .X(_00768_));
 sky130_fd_sc_hd__mux2_1 _09777_ (.A0(\core_pipeline.pipeline_registers.registers[21][13] ),
    .A1(net321),
    .S(net201),
    .X(_00769_));
 sky130_fd_sc_hd__mux2_1 _09778_ (.A0(\core_pipeline.pipeline_registers.registers[21][14] ),
    .A1(net319),
    .S(net201),
    .X(_00770_));
 sky130_fd_sc_hd__mux2_1 _09779_ (.A0(\core_pipeline.pipeline_registers.registers[21][15] ),
    .A1(net318),
    .S(net201),
    .X(_00771_));
 sky130_fd_sc_hd__mux2_1 _09780_ (.A0(\core_pipeline.pipeline_registers.registers[21][16] ),
    .A1(net316),
    .S(net201),
    .X(_00772_));
 sky130_fd_sc_hd__mux2_1 _09781_ (.A0(\core_pipeline.pipeline_registers.registers[21][17] ),
    .A1(net314),
    .S(net202),
    .X(_00773_));
 sky130_fd_sc_hd__mux2_1 _09782_ (.A0(\core_pipeline.pipeline_registers.registers[21][18] ),
    .A1(_03976_),
    .S(net202),
    .X(_00774_));
 sky130_fd_sc_hd__mux2_1 _09783_ (.A0(\core_pipeline.pipeline_registers.registers[21][19] ),
    .A1(net309),
    .S(net202),
    .X(_00775_));
 sky130_fd_sc_hd__mux2_1 _09784_ (.A0(\core_pipeline.pipeline_registers.registers[21][20] ),
    .A1(net305),
    .S(net202),
    .X(_00776_));
 sky130_fd_sc_hd__mux2_1 _09785_ (.A0(\core_pipeline.pipeline_registers.registers[21][21] ),
    .A1(net304),
    .S(net202),
    .X(_00777_));
 sky130_fd_sc_hd__mux2_1 _09786_ (.A0(\core_pipeline.pipeline_registers.registers[21][22] ),
    .A1(net302),
    .S(net202),
    .X(_00778_));
 sky130_fd_sc_hd__mux2_1 _09787_ (.A0(\core_pipeline.pipeline_registers.registers[21][23] ),
    .A1(net299),
    .S(net202),
    .X(_00779_));
 sky130_fd_sc_hd__mux2_1 _09788_ (.A0(\core_pipeline.pipeline_registers.registers[21][24] ),
    .A1(net298),
    .S(net201),
    .X(_00780_));
 sky130_fd_sc_hd__mux2_1 _09789_ (.A0(\core_pipeline.pipeline_registers.registers[21][25] ),
    .A1(net295),
    .S(net201),
    .X(_00781_));
 sky130_fd_sc_hd__mux2_1 _09790_ (.A0(\core_pipeline.pipeline_registers.registers[21][26] ),
    .A1(net293),
    .S(net201),
    .X(_00782_));
 sky130_fd_sc_hd__mux2_1 _09791_ (.A0(\core_pipeline.pipeline_registers.registers[21][27] ),
    .A1(net291),
    .S(net202),
    .X(_00783_));
 sky130_fd_sc_hd__mux2_1 _09792_ (.A0(\core_pipeline.pipeline_registers.registers[21][28] ),
    .A1(net290),
    .S(net202),
    .X(_00784_));
 sky130_fd_sc_hd__mux2_1 _09793_ (.A0(\core_pipeline.pipeline_registers.registers[21][29] ),
    .A1(net287),
    .S(net202),
    .X(_00785_));
 sky130_fd_sc_hd__mux2_1 _09794_ (.A0(\core_pipeline.pipeline_registers.registers[21][30] ),
    .A1(net285),
    .S(net202),
    .X(_00786_));
 sky130_fd_sc_hd__mux2_1 _09795_ (.A0(\core_pipeline.pipeline_registers.registers[21][31] ),
    .A1(net283),
    .S(net202),
    .X(_00787_));
 sky130_fd_sc_hd__nor2_8 _09796_ (.A(_04934_),
    .B(_05592_),
    .Y(_05595_));
 sky130_fd_sc_hd__mux2_1 _09797_ (.A0(\core_pipeline.pipeline_registers.registers[22][0] ),
    .A1(net349),
    .S(net199),
    .X(_00788_));
 sky130_fd_sc_hd__mux2_1 _09798_ (.A0(\core_pipeline.pipeline_registers.registers[22][1] ),
    .A1(net347),
    .S(net200),
    .X(_00789_));
 sky130_fd_sc_hd__mux2_1 _09799_ (.A0(\core_pipeline.pipeline_registers.registers[22][2] ),
    .A1(net345),
    .S(net200),
    .X(_00790_));
 sky130_fd_sc_hd__mux2_1 _09800_ (.A0(\core_pipeline.pipeline_registers.registers[22][3] ),
    .A1(net342),
    .S(net199),
    .X(_00791_));
 sky130_fd_sc_hd__mux2_1 _09801_ (.A0(\core_pipeline.pipeline_registers.registers[22][4] ),
    .A1(net340),
    .S(net199),
    .X(_00792_));
 sky130_fd_sc_hd__mux2_1 _09802_ (.A0(\core_pipeline.pipeline_registers.registers[22][5] ),
    .A1(net339),
    .S(net200),
    .X(_00793_));
 sky130_fd_sc_hd__mux2_1 _09803_ (.A0(\core_pipeline.pipeline_registers.registers[22][6] ),
    .A1(net336),
    .S(net199),
    .X(_00794_));
 sky130_fd_sc_hd__mux2_1 _09804_ (.A0(\core_pipeline.pipeline_registers.registers[22][7] ),
    .A1(net333),
    .S(net199),
    .X(_00795_));
 sky130_fd_sc_hd__mux2_1 _09805_ (.A0(\core_pipeline.pipeline_registers.registers[22][8] ),
    .A1(net331),
    .S(net199),
    .X(_00796_));
 sky130_fd_sc_hd__mux2_1 _09806_ (.A0(\core_pipeline.pipeline_registers.registers[22][9] ),
    .A1(net329),
    .S(net199),
    .X(_00797_));
 sky130_fd_sc_hd__mux2_1 _09807_ (.A0(\core_pipeline.pipeline_registers.registers[22][10] ),
    .A1(net327),
    .S(net199),
    .X(_00798_));
 sky130_fd_sc_hd__mux2_1 _09808_ (.A0(\core_pipeline.pipeline_registers.registers[22][11] ),
    .A1(net326),
    .S(net199),
    .X(_00799_));
 sky130_fd_sc_hd__mux2_1 _09809_ (.A0(\core_pipeline.pipeline_registers.registers[22][12] ),
    .A1(net323),
    .S(net199),
    .X(_00800_));
 sky130_fd_sc_hd__mux2_1 _09810_ (.A0(\core_pipeline.pipeline_registers.registers[22][13] ),
    .A1(net321),
    .S(net199),
    .X(_00801_));
 sky130_fd_sc_hd__mux2_1 _09811_ (.A0(\core_pipeline.pipeline_registers.registers[22][14] ),
    .A1(net319),
    .S(net199),
    .X(_00802_));
 sky130_fd_sc_hd__mux2_1 _09812_ (.A0(\core_pipeline.pipeline_registers.registers[22][15] ),
    .A1(net317),
    .S(net199),
    .X(_00803_));
 sky130_fd_sc_hd__mux2_1 _09813_ (.A0(\core_pipeline.pipeline_registers.registers[22][16] ),
    .A1(net316),
    .S(net199),
    .X(_00804_));
 sky130_fd_sc_hd__mux2_1 _09814_ (.A0(\core_pipeline.pipeline_registers.registers[22][17] ),
    .A1(net314),
    .S(net200),
    .X(_00805_));
 sky130_fd_sc_hd__mux2_1 _09815_ (.A0(\core_pipeline.pipeline_registers.registers[22][18] ),
    .A1(net310),
    .S(net200),
    .X(_00806_));
 sky130_fd_sc_hd__mux2_1 _09816_ (.A0(\core_pipeline.pipeline_registers.registers[22][19] ),
    .A1(net309),
    .S(net200),
    .X(_00807_));
 sky130_fd_sc_hd__mux2_1 _09817_ (.A0(\core_pipeline.pipeline_registers.registers[22][20] ),
    .A1(net307),
    .S(net200),
    .X(_00808_));
 sky130_fd_sc_hd__mux2_1 _09818_ (.A0(\core_pipeline.pipeline_registers.registers[22][21] ),
    .A1(net304),
    .S(net200),
    .X(_00809_));
 sky130_fd_sc_hd__mux2_1 _09819_ (.A0(\core_pipeline.pipeline_registers.registers[22][22] ),
    .A1(net302),
    .S(net200),
    .X(_00810_));
 sky130_fd_sc_hd__mux2_1 _09820_ (.A0(\core_pipeline.pipeline_registers.registers[22][23] ),
    .A1(net299),
    .S(net200),
    .X(_00811_));
 sky130_fd_sc_hd__mux2_1 _09821_ (.A0(\core_pipeline.pipeline_registers.registers[22][24] ),
    .A1(net297),
    .S(net199),
    .X(_00812_));
 sky130_fd_sc_hd__mux2_1 _09822_ (.A0(\core_pipeline.pipeline_registers.registers[22][25] ),
    .A1(net295),
    .S(net199),
    .X(_00813_));
 sky130_fd_sc_hd__mux2_1 _09823_ (.A0(\core_pipeline.pipeline_registers.registers[22][26] ),
    .A1(net293),
    .S(net199),
    .X(_00814_));
 sky130_fd_sc_hd__mux2_1 _09824_ (.A0(\core_pipeline.pipeline_registers.registers[22][27] ),
    .A1(net291),
    .S(net200),
    .X(_00815_));
 sky130_fd_sc_hd__mux2_1 _09825_ (.A0(\core_pipeline.pipeline_registers.registers[22][28] ),
    .A1(net290),
    .S(net200),
    .X(_00816_));
 sky130_fd_sc_hd__mux2_1 _09826_ (.A0(\core_pipeline.pipeline_registers.registers[22][29] ),
    .A1(net287),
    .S(net200),
    .X(_00817_));
 sky130_fd_sc_hd__mux2_1 _09827_ (.A0(\core_pipeline.pipeline_registers.registers[22][30] ),
    .A1(net284),
    .S(net200),
    .X(_00818_));
 sky130_fd_sc_hd__mux2_1 _09828_ (.A0(\core_pipeline.pipeline_registers.registers[22][31] ),
    .A1(net283),
    .S(net200),
    .X(_00819_));
 sky130_fd_sc_hd__or3_1 _09829_ (.A(net126),
    .B(_03445_),
    .C(_03638_),
    .X(_05596_));
 sky130_fd_sc_hd__o21a_1 _09830_ (.A1(net630),
    .A2(net142),
    .B1(_05596_),
    .X(_00820_));
 sky130_fd_sc_hd__nor2_8 _09831_ (.A(_03915_),
    .B(_04937_),
    .Y(_05597_));
 sky130_fd_sc_hd__mux2_1 _09832_ (.A0(\core_pipeline.pipeline_registers.registers[3][0] ),
    .A1(net348),
    .S(net243),
    .X(_00821_));
 sky130_fd_sc_hd__mux2_1 _09833_ (.A0(\core_pipeline.pipeline_registers.registers[3][1] ),
    .A1(net347),
    .S(net244),
    .X(_00822_));
 sky130_fd_sc_hd__mux2_1 _09834_ (.A0(\core_pipeline.pipeline_registers.registers[3][2] ),
    .A1(net345),
    .S(net244),
    .X(_00823_));
 sky130_fd_sc_hd__mux2_1 _09835_ (.A0(\core_pipeline.pipeline_registers.registers[3][3] ),
    .A1(net342),
    .S(net243),
    .X(_00824_));
 sky130_fd_sc_hd__mux2_1 _09836_ (.A0(\core_pipeline.pipeline_registers.registers[3][4] ),
    .A1(net340),
    .S(net243),
    .X(_00825_));
 sky130_fd_sc_hd__mux2_1 _09837_ (.A0(\core_pipeline.pipeline_registers.registers[3][5] ),
    .A1(net338),
    .S(net244),
    .X(_00826_));
 sky130_fd_sc_hd__mux2_1 _09838_ (.A0(\core_pipeline.pipeline_registers.registers[3][6] ),
    .A1(net335),
    .S(net243),
    .X(_00827_));
 sky130_fd_sc_hd__mux2_1 _09839_ (.A0(\core_pipeline.pipeline_registers.registers[3][7] ),
    .A1(net334),
    .S(net243),
    .X(_00828_));
 sky130_fd_sc_hd__mux2_1 _09840_ (.A0(\core_pipeline.pipeline_registers.registers[3][8] ),
    .A1(net332),
    .S(net243),
    .X(_00829_));
 sky130_fd_sc_hd__mux2_1 _09841_ (.A0(\core_pipeline.pipeline_registers.registers[3][9] ),
    .A1(net329),
    .S(net243),
    .X(_00830_));
 sky130_fd_sc_hd__mux2_1 _09842_ (.A0(\core_pipeline.pipeline_registers.registers[3][10] ),
    .A1(net327),
    .S(net243),
    .X(_00831_));
 sky130_fd_sc_hd__mux2_1 _09843_ (.A0(\core_pipeline.pipeline_registers.registers[3][11] ),
    .A1(net325),
    .S(net243),
    .X(_00832_));
 sky130_fd_sc_hd__mux2_1 _09844_ (.A0(\core_pipeline.pipeline_registers.registers[3][12] ),
    .A1(net324),
    .S(net243),
    .X(_00833_));
 sky130_fd_sc_hd__mux2_1 _09845_ (.A0(\core_pipeline.pipeline_registers.registers[3][13] ),
    .A1(net322),
    .S(net243),
    .X(_00834_));
 sky130_fd_sc_hd__mux2_1 _09846_ (.A0(\core_pipeline.pipeline_registers.registers[3][14] ),
    .A1(net320),
    .S(net243),
    .X(_00835_));
 sky130_fd_sc_hd__mux2_1 _09847_ (.A0(\core_pipeline.pipeline_registers.registers[3][15] ),
    .A1(net317),
    .S(net243),
    .X(_00836_));
 sky130_fd_sc_hd__mux2_1 _09848_ (.A0(\core_pipeline.pipeline_registers.registers[3][16] ),
    .A1(net315),
    .S(net243),
    .X(_00837_));
 sky130_fd_sc_hd__mux2_1 _09849_ (.A0(\core_pipeline.pipeline_registers.registers[3][17] ),
    .A1(net312),
    .S(net244),
    .X(_00838_));
 sky130_fd_sc_hd__mux2_1 _09850_ (.A0(\core_pipeline.pipeline_registers.registers[3][18] ),
    .A1(net311),
    .S(net244),
    .X(_00839_));
 sky130_fd_sc_hd__mux2_1 _09851_ (.A0(\core_pipeline.pipeline_registers.registers[3][19] ),
    .A1(net308),
    .S(net244),
    .X(_00840_));
 sky130_fd_sc_hd__mux2_1 _09852_ (.A0(\core_pipeline.pipeline_registers.registers[3][20] ),
    .A1(net305),
    .S(net244),
    .X(_00841_));
 sky130_fd_sc_hd__mux2_1 _09853_ (.A0(\core_pipeline.pipeline_registers.registers[3][21] ),
    .A1(net303),
    .S(net244),
    .X(_00842_));
 sky130_fd_sc_hd__mux2_1 _09854_ (.A0(\core_pipeline.pipeline_registers.registers[3][22] ),
    .A1(net301),
    .S(net244),
    .X(_00843_));
 sky130_fd_sc_hd__mux2_1 _09855_ (.A0(\core_pipeline.pipeline_registers.registers[3][23] ),
    .A1(net300),
    .S(net244),
    .X(_00844_));
 sky130_fd_sc_hd__mux2_1 _09856_ (.A0(\core_pipeline.pipeline_registers.registers[3][24] ),
    .A1(net298),
    .S(net243),
    .X(_00845_));
 sky130_fd_sc_hd__mux2_1 _09857_ (.A0(\core_pipeline.pipeline_registers.registers[3][25] ),
    .A1(net296),
    .S(net243),
    .X(_00846_));
 sky130_fd_sc_hd__mux2_1 _09858_ (.A0(\core_pipeline.pipeline_registers.registers[3][26] ),
    .A1(net293),
    .S(net243),
    .X(_00847_));
 sky130_fd_sc_hd__mux2_1 _09859_ (.A0(\core_pipeline.pipeline_registers.registers[3][27] ),
    .A1(net292),
    .S(net244),
    .X(_00848_));
 sky130_fd_sc_hd__mux2_1 _09860_ (.A0(\core_pipeline.pipeline_registers.registers[3][28] ),
    .A1(net289),
    .S(net244),
    .X(_00849_));
 sky130_fd_sc_hd__mux2_1 _09861_ (.A0(\core_pipeline.pipeline_registers.registers[3][29] ),
    .A1(net288),
    .S(net244),
    .X(_00850_));
 sky130_fd_sc_hd__mux2_1 _09862_ (.A0(\core_pipeline.pipeline_registers.registers[3][30] ),
    .A1(net284),
    .S(net244),
    .X(_00851_));
 sky130_fd_sc_hd__mux2_1 _09863_ (.A0(\core_pipeline.pipeline_registers.registers[3][31] ),
    .A1(net283),
    .S(net244),
    .X(_00852_));
 sky130_fd_sc_hd__and3b_4 _09864_ (.A_N(_04936_),
    .B(_04468_),
    .C(_03912_),
    .X(_05598_));
 sky130_fd_sc_hd__nand2b_4 _09865_ (.A_N(_04939_),
    .B(_05598_),
    .Y(_05599_));
 sky130_fd_sc_hd__mux2_1 _09866_ (.A0(net348),
    .A1(\core_pipeline.pipeline_registers.registers[4][0] ),
    .S(net197),
    .X(_00853_));
 sky130_fd_sc_hd__mux2_1 _09867_ (.A0(net346),
    .A1(\core_pipeline.pipeline_registers.registers[4][1] ),
    .S(net198),
    .X(_00854_));
 sky130_fd_sc_hd__mux2_1 _09868_ (.A0(net345),
    .A1(\core_pipeline.pipeline_registers.registers[4][2] ),
    .S(net198),
    .X(_00855_));
 sky130_fd_sc_hd__mux2_1 _09869_ (.A0(net342),
    .A1(\core_pipeline.pipeline_registers.registers[4][3] ),
    .S(net197),
    .X(_00856_));
 sky130_fd_sc_hd__mux2_1 _09870_ (.A0(net340),
    .A1(\core_pipeline.pipeline_registers.registers[4][4] ),
    .S(net197),
    .X(_00857_));
 sky130_fd_sc_hd__mux2_1 _09871_ (.A0(net337),
    .A1(\core_pipeline.pipeline_registers.registers[4][5] ),
    .S(net198),
    .X(_00858_));
 sky130_fd_sc_hd__mux2_1 _09872_ (.A0(net335),
    .A1(\core_pipeline.pipeline_registers.registers[4][6] ),
    .S(net197),
    .X(_00859_));
 sky130_fd_sc_hd__mux2_1 _09873_ (.A0(net334),
    .A1(\core_pipeline.pipeline_registers.registers[4][7] ),
    .S(net197),
    .X(_00860_));
 sky130_fd_sc_hd__mux2_1 _09874_ (.A0(net332),
    .A1(\core_pipeline.pipeline_registers.registers[4][8] ),
    .S(net197),
    .X(_00861_));
 sky130_fd_sc_hd__mux2_1 _09875_ (.A0(net329),
    .A1(\core_pipeline.pipeline_registers.registers[4][9] ),
    .S(net197),
    .X(_00862_));
 sky130_fd_sc_hd__mux2_1 _09876_ (.A0(net328),
    .A1(\core_pipeline.pipeline_registers.registers[4][10] ),
    .S(net197),
    .X(_00863_));
 sky130_fd_sc_hd__mux2_1 _09877_ (.A0(net325),
    .A1(\core_pipeline.pipeline_registers.registers[4][11] ),
    .S(net197),
    .X(_00864_));
 sky130_fd_sc_hd__mux2_1 _09878_ (.A0(net323),
    .A1(\core_pipeline.pipeline_registers.registers[4][12] ),
    .S(net197),
    .X(_00865_));
 sky130_fd_sc_hd__mux2_1 _09879_ (.A0(net322),
    .A1(\core_pipeline.pipeline_registers.registers[4][13] ),
    .S(net197),
    .X(_00866_));
 sky130_fd_sc_hd__mux2_1 _09880_ (.A0(net320),
    .A1(\core_pipeline.pipeline_registers.registers[4][14] ),
    .S(net197),
    .X(_00867_));
 sky130_fd_sc_hd__mux2_1 _09881_ (.A0(net317),
    .A1(\core_pipeline.pipeline_registers.registers[4][15] ),
    .S(net197),
    .X(_00868_));
 sky130_fd_sc_hd__mux2_1 _09882_ (.A0(net315),
    .A1(\core_pipeline.pipeline_registers.registers[4][16] ),
    .S(net197),
    .X(_00869_));
 sky130_fd_sc_hd__mux2_1 _09883_ (.A0(net312),
    .A1(\core_pipeline.pipeline_registers.registers[4][17] ),
    .S(net198),
    .X(_00870_));
 sky130_fd_sc_hd__mux2_1 _09884_ (.A0(_03976_),
    .A1(\core_pipeline.pipeline_registers.registers[4][18] ),
    .S(net198),
    .X(_00871_));
 sky130_fd_sc_hd__mux2_1 _09885_ (.A0(net309),
    .A1(\core_pipeline.pipeline_registers.registers[4][19] ),
    .S(net198),
    .X(_00872_));
 sky130_fd_sc_hd__mux2_1 _09886_ (.A0(net306),
    .A1(\core_pipeline.pipeline_registers.registers[4][20] ),
    .S(net198),
    .X(_00873_));
 sky130_fd_sc_hd__mux2_1 _09887_ (.A0(net303),
    .A1(\core_pipeline.pipeline_registers.registers[4][21] ),
    .S(net198),
    .X(_00874_));
 sky130_fd_sc_hd__mux2_1 _09888_ (.A0(net301),
    .A1(\core_pipeline.pipeline_registers.registers[4][22] ),
    .S(net198),
    .X(_00875_));
 sky130_fd_sc_hd__mux2_1 _09889_ (.A0(net300),
    .A1(\core_pipeline.pipeline_registers.registers[4][23] ),
    .S(net198),
    .X(_00876_));
 sky130_fd_sc_hd__mux2_1 _09890_ (.A0(net297),
    .A1(\core_pipeline.pipeline_registers.registers[4][24] ),
    .S(net197),
    .X(_00877_));
 sky130_fd_sc_hd__mux2_1 _09891_ (.A0(net295),
    .A1(\core_pipeline.pipeline_registers.registers[4][25] ),
    .S(net197),
    .X(_00878_));
 sky130_fd_sc_hd__mux2_1 _09892_ (.A0(net293),
    .A1(\core_pipeline.pipeline_registers.registers[4][26] ),
    .S(net197),
    .X(_00879_));
 sky130_fd_sc_hd__mux2_1 _09893_ (.A0(net291),
    .A1(\core_pipeline.pipeline_registers.registers[4][27] ),
    .S(net198),
    .X(_00880_));
 sky130_fd_sc_hd__mux2_1 _09894_ (.A0(net289),
    .A1(\core_pipeline.pipeline_registers.registers[4][28] ),
    .S(net198),
    .X(_00881_));
 sky130_fd_sc_hd__mux2_1 _09895_ (.A0(net288),
    .A1(\core_pipeline.pipeline_registers.registers[4][29] ),
    .S(net198),
    .X(_00882_));
 sky130_fd_sc_hd__mux2_1 _09896_ (.A0(net285),
    .A1(\core_pipeline.pipeline_registers.registers[4][30] ),
    .S(net198),
    .X(_00883_));
 sky130_fd_sc_hd__mux2_1 _09897_ (.A0(net282),
    .A1(\core_pipeline.pipeline_registers.registers[4][31] ),
    .S(net198),
    .X(_00884_));
 sky130_fd_sc_hd__nand2b_4 _09898_ (.A_N(_05589_),
    .B(_05598_),
    .Y(_05600_));
 sky130_fd_sc_hd__mux2_1 _09899_ (.A0(net348),
    .A1(\core_pipeline.pipeline_registers.registers[5][0] ),
    .S(net195),
    .X(_00885_));
 sky130_fd_sc_hd__mux2_1 _09900_ (.A0(net346),
    .A1(\core_pipeline.pipeline_registers.registers[5][1] ),
    .S(net196),
    .X(_00886_));
 sky130_fd_sc_hd__mux2_1 _09901_ (.A0(net345),
    .A1(\core_pipeline.pipeline_registers.registers[5][2] ),
    .S(net196),
    .X(_00887_));
 sky130_fd_sc_hd__mux2_1 _09902_ (.A0(net343),
    .A1(\core_pipeline.pipeline_registers.registers[5][3] ),
    .S(net195),
    .X(_00888_));
 sky130_fd_sc_hd__mux2_1 _09903_ (.A0(net341),
    .A1(\core_pipeline.pipeline_registers.registers[5][4] ),
    .S(net195),
    .X(_00889_));
 sky130_fd_sc_hd__mux2_1 _09904_ (.A0(net337),
    .A1(\core_pipeline.pipeline_registers.registers[5][5] ),
    .S(net196),
    .X(_00890_));
 sky130_fd_sc_hd__mux2_1 _09905_ (.A0(net335),
    .A1(\core_pipeline.pipeline_registers.registers[5][6] ),
    .S(net195),
    .X(_00891_));
 sky130_fd_sc_hd__mux2_1 _09906_ (.A0(net334),
    .A1(\core_pipeline.pipeline_registers.registers[5][7] ),
    .S(net195),
    .X(_00892_));
 sky130_fd_sc_hd__mux2_1 _09907_ (.A0(net332),
    .A1(\core_pipeline.pipeline_registers.registers[5][8] ),
    .S(net195),
    .X(_00893_));
 sky130_fd_sc_hd__mux2_1 _09908_ (.A0(net329),
    .A1(\core_pipeline.pipeline_registers.registers[5][9] ),
    .S(net195),
    .X(_00894_));
 sky130_fd_sc_hd__mux2_1 _09909_ (.A0(net328),
    .A1(\core_pipeline.pipeline_registers.registers[5][10] ),
    .S(net195),
    .X(_00895_));
 sky130_fd_sc_hd__mux2_1 _09910_ (.A0(net325),
    .A1(\core_pipeline.pipeline_registers.registers[5][11] ),
    .S(net195),
    .X(_00896_));
 sky130_fd_sc_hd__mux2_1 _09911_ (.A0(net323),
    .A1(\core_pipeline.pipeline_registers.registers[5][12] ),
    .S(net195),
    .X(_00897_));
 sky130_fd_sc_hd__mux2_1 _09912_ (.A0(net322),
    .A1(\core_pipeline.pipeline_registers.registers[5][13] ),
    .S(net195),
    .X(_00898_));
 sky130_fd_sc_hd__mux2_1 _09913_ (.A0(net320),
    .A1(\core_pipeline.pipeline_registers.registers[5][14] ),
    .S(net195),
    .X(_00899_));
 sky130_fd_sc_hd__mux2_1 _09914_ (.A0(net317),
    .A1(\core_pipeline.pipeline_registers.registers[5][15] ),
    .S(net195),
    .X(_00900_));
 sky130_fd_sc_hd__mux2_1 _09915_ (.A0(net315),
    .A1(\core_pipeline.pipeline_registers.registers[5][16] ),
    .S(net195),
    .X(_00901_));
 sky130_fd_sc_hd__mux2_1 _09916_ (.A0(net312),
    .A1(\core_pipeline.pipeline_registers.registers[5][17] ),
    .S(net196),
    .X(_00902_));
 sky130_fd_sc_hd__mux2_1 _09917_ (.A0(_03976_),
    .A1(\core_pipeline.pipeline_registers.registers[5][18] ),
    .S(net196),
    .X(_00903_));
 sky130_fd_sc_hd__mux2_1 _09918_ (.A0(net309),
    .A1(\core_pipeline.pipeline_registers.registers[5][19] ),
    .S(net196),
    .X(_00904_));
 sky130_fd_sc_hd__mux2_1 _09919_ (.A0(net306),
    .A1(\core_pipeline.pipeline_registers.registers[5][20] ),
    .S(net196),
    .X(_00905_));
 sky130_fd_sc_hd__mux2_1 _09920_ (.A0(net304),
    .A1(\core_pipeline.pipeline_registers.registers[5][21] ),
    .S(net196),
    .X(_00906_));
 sky130_fd_sc_hd__mux2_1 _09921_ (.A0(net301),
    .A1(\core_pipeline.pipeline_registers.registers[5][22] ),
    .S(net196),
    .X(_00907_));
 sky130_fd_sc_hd__mux2_1 _09922_ (.A0(net300),
    .A1(\core_pipeline.pipeline_registers.registers[5][23] ),
    .S(net196),
    .X(_00908_));
 sky130_fd_sc_hd__mux2_1 _09923_ (.A0(net297),
    .A1(\core_pipeline.pipeline_registers.registers[5][24] ),
    .S(net195),
    .X(_00909_));
 sky130_fd_sc_hd__mux2_1 _09924_ (.A0(net296),
    .A1(\core_pipeline.pipeline_registers.registers[5][25] ),
    .S(net195),
    .X(_00910_));
 sky130_fd_sc_hd__mux2_1 _09925_ (.A0(net294),
    .A1(\core_pipeline.pipeline_registers.registers[5][26] ),
    .S(net195),
    .X(_00911_));
 sky130_fd_sc_hd__mux2_1 _09926_ (.A0(net292),
    .A1(\core_pipeline.pipeline_registers.registers[5][27] ),
    .S(net196),
    .X(_00912_));
 sky130_fd_sc_hd__mux2_1 _09927_ (.A0(net289),
    .A1(\core_pipeline.pipeline_registers.registers[5][28] ),
    .S(net196),
    .X(_00913_));
 sky130_fd_sc_hd__mux2_1 _09928_ (.A0(net288),
    .A1(\core_pipeline.pipeline_registers.registers[5][29] ),
    .S(net196),
    .X(_00914_));
 sky130_fd_sc_hd__mux2_1 _09929_ (.A0(net285),
    .A1(\core_pipeline.pipeline_registers.registers[5][30] ),
    .S(net196),
    .X(_00915_));
 sky130_fd_sc_hd__mux2_1 _09930_ (.A0(net282),
    .A1(\core_pipeline.pipeline_registers.registers[5][31] ),
    .S(net196),
    .X(_00916_));
 sky130_fd_sc_hd__nand2b_4 _09931_ (.A_N(_04934_),
    .B(_05598_),
    .Y(_05601_));
 sky130_fd_sc_hd__mux2_1 _09932_ (.A0(net348),
    .A1(\core_pipeline.pipeline_registers.registers[6][0] ),
    .S(net193),
    .X(_00917_));
 sky130_fd_sc_hd__mux2_1 _09933_ (.A0(net347),
    .A1(\core_pipeline.pipeline_registers.registers[6][1] ),
    .S(net194),
    .X(_00918_));
 sky130_fd_sc_hd__mux2_1 _09934_ (.A0(net345),
    .A1(\core_pipeline.pipeline_registers.registers[6][2] ),
    .S(net194),
    .X(_00919_));
 sky130_fd_sc_hd__mux2_1 _09935_ (.A0(net343),
    .A1(\core_pipeline.pipeline_registers.registers[6][3] ),
    .S(net193),
    .X(_00920_));
 sky130_fd_sc_hd__mux2_1 _09936_ (.A0(net340),
    .A1(\core_pipeline.pipeline_registers.registers[6][4] ),
    .S(net193),
    .X(_00921_));
 sky130_fd_sc_hd__mux2_1 _09937_ (.A0(net337),
    .A1(\core_pipeline.pipeline_registers.registers[6][5] ),
    .S(net194),
    .X(_00922_));
 sky130_fd_sc_hd__mux2_1 _09938_ (.A0(net335),
    .A1(\core_pipeline.pipeline_registers.registers[6][6] ),
    .S(net193),
    .X(_00923_));
 sky130_fd_sc_hd__mux2_1 _09939_ (.A0(net334),
    .A1(\core_pipeline.pipeline_registers.registers[6][7] ),
    .S(net193),
    .X(_00924_));
 sky130_fd_sc_hd__mux2_1 _09940_ (.A0(net332),
    .A1(\core_pipeline.pipeline_registers.registers[6][8] ),
    .S(net193),
    .X(_00925_));
 sky130_fd_sc_hd__mux2_1 _09941_ (.A0(net329),
    .A1(\core_pipeline.pipeline_registers.registers[6][9] ),
    .S(net193),
    .X(_00926_));
 sky130_fd_sc_hd__mux2_1 _09942_ (.A0(net328),
    .A1(\core_pipeline.pipeline_registers.registers[6][10] ),
    .S(net193),
    .X(_00927_));
 sky130_fd_sc_hd__mux2_1 _09943_ (.A0(net325),
    .A1(\core_pipeline.pipeline_registers.registers[6][11] ),
    .S(net193),
    .X(_00928_));
 sky130_fd_sc_hd__mux2_1 _09944_ (.A0(net323),
    .A1(\core_pipeline.pipeline_registers.registers[6][12] ),
    .S(net193),
    .X(_00929_));
 sky130_fd_sc_hd__mux2_1 _09945_ (.A0(net322),
    .A1(\core_pipeline.pipeline_registers.registers[6][13] ),
    .S(net193),
    .X(_00930_));
 sky130_fd_sc_hd__mux2_1 _09946_ (.A0(net320),
    .A1(\core_pipeline.pipeline_registers.registers[6][14] ),
    .S(net193),
    .X(_00931_));
 sky130_fd_sc_hd__mux2_1 _09947_ (.A0(net317),
    .A1(\core_pipeline.pipeline_registers.registers[6][15] ),
    .S(net193),
    .X(_00932_));
 sky130_fd_sc_hd__mux2_1 _09948_ (.A0(net315),
    .A1(\core_pipeline.pipeline_registers.registers[6][16] ),
    .S(net193),
    .X(_00933_));
 sky130_fd_sc_hd__mux2_1 _09949_ (.A0(net312),
    .A1(\core_pipeline.pipeline_registers.registers[6][17] ),
    .S(net194),
    .X(_00934_));
 sky130_fd_sc_hd__mux2_1 _09950_ (.A0(net310),
    .A1(\core_pipeline.pipeline_registers.registers[6][18] ),
    .S(net194),
    .X(_00935_));
 sky130_fd_sc_hd__mux2_1 _09951_ (.A0(net308),
    .A1(\core_pipeline.pipeline_registers.registers[6][19] ),
    .S(net194),
    .X(_00936_));
 sky130_fd_sc_hd__mux2_1 _09952_ (.A0(net305),
    .A1(\core_pipeline.pipeline_registers.registers[6][20] ),
    .S(net194),
    .X(_00937_));
 sky130_fd_sc_hd__mux2_1 _09953_ (.A0(net303),
    .A1(\core_pipeline.pipeline_registers.registers[6][21] ),
    .S(net194),
    .X(_00938_));
 sky130_fd_sc_hd__mux2_1 _09954_ (.A0(net301),
    .A1(\core_pipeline.pipeline_registers.registers[6][22] ),
    .S(net194),
    .X(_00939_));
 sky130_fd_sc_hd__mux2_1 _09955_ (.A0(net300),
    .A1(\core_pipeline.pipeline_registers.registers[6][23] ),
    .S(net194),
    .X(_00940_));
 sky130_fd_sc_hd__mux2_1 _09956_ (.A0(net297),
    .A1(\core_pipeline.pipeline_registers.registers[6][24] ),
    .S(net193),
    .X(_00941_));
 sky130_fd_sc_hd__mux2_1 _09957_ (.A0(net295),
    .A1(\core_pipeline.pipeline_registers.registers[6][25] ),
    .S(net193),
    .X(_00942_));
 sky130_fd_sc_hd__mux2_1 _09958_ (.A0(net294),
    .A1(\core_pipeline.pipeline_registers.registers[6][26] ),
    .S(net193),
    .X(_00943_));
 sky130_fd_sc_hd__mux2_1 _09959_ (.A0(net292),
    .A1(\core_pipeline.pipeline_registers.registers[6][27] ),
    .S(net194),
    .X(_00944_));
 sky130_fd_sc_hd__mux2_1 _09960_ (.A0(net289),
    .A1(\core_pipeline.pipeline_registers.registers[6][28] ),
    .S(net194),
    .X(_00945_));
 sky130_fd_sc_hd__mux2_1 _09961_ (.A0(net288),
    .A1(\core_pipeline.pipeline_registers.registers[6][29] ),
    .S(net194),
    .X(_00946_));
 sky130_fd_sc_hd__mux2_1 _09962_ (.A0(net285),
    .A1(\core_pipeline.pipeline_registers.registers[6][30] ),
    .S(net194),
    .X(_00947_));
 sky130_fd_sc_hd__mux2_1 _09963_ (.A0(net282),
    .A1(\core_pipeline.pipeline_registers.registers[6][31] ),
    .S(net194),
    .X(_00948_));
 sky130_fd_sc_hd__nand2b_4 _09964_ (.A_N(_03915_),
    .B(_05598_),
    .Y(_05602_));
 sky130_fd_sc_hd__mux2_1 _09965_ (.A0(net348),
    .A1(\core_pipeline.pipeline_registers.registers[7][0] ),
    .S(net191),
    .X(_00949_));
 sky130_fd_sc_hd__mux2_1 _09966_ (.A0(net346),
    .A1(\core_pipeline.pipeline_registers.registers[7][1] ),
    .S(net192),
    .X(_00950_));
 sky130_fd_sc_hd__mux2_1 _09967_ (.A0(net345),
    .A1(\core_pipeline.pipeline_registers.registers[7][2] ),
    .S(net192),
    .X(_00951_));
 sky130_fd_sc_hd__mux2_1 _09968_ (.A0(net343),
    .A1(\core_pipeline.pipeline_registers.registers[7][3] ),
    .S(net191),
    .X(_00952_));
 sky130_fd_sc_hd__mux2_1 _09969_ (.A0(net341),
    .A1(\core_pipeline.pipeline_registers.registers[7][4] ),
    .S(net191),
    .X(_00953_));
 sky130_fd_sc_hd__mux2_1 _09970_ (.A0(net337),
    .A1(\core_pipeline.pipeline_registers.registers[7][5] ),
    .S(net192),
    .X(_00954_));
 sky130_fd_sc_hd__mux2_1 _09971_ (.A0(net335),
    .A1(\core_pipeline.pipeline_registers.registers[7][6] ),
    .S(net191),
    .X(_00955_));
 sky130_fd_sc_hd__mux2_1 _09972_ (.A0(net334),
    .A1(\core_pipeline.pipeline_registers.registers[7][7] ),
    .S(net191),
    .X(_00956_));
 sky130_fd_sc_hd__mux2_1 _09973_ (.A0(net332),
    .A1(\core_pipeline.pipeline_registers.registers[7][8] ),
    .S(net191),
    .X(_00957_));
 sky130_fd_sc_hd__mux2_1 _09974_ (.A0(net329),
    .A1(\core_pipeline.pipeline_registers.registers[7][9] ),
    .S(net191),
    .X(_00958_));
 sky130_fd_sc_hd__mux2_1 _09975_ (.A0(net327),
    .A1(\core_pipeline.pipeline_registers.registers[7][10] ),
    .S(net191),
    .X(_00959_));
 sky130_fd_sc_hd__mux2_1 _09976_ (.A0(net325),
    .A1(\core_pipeline.pipeline_registers.registers[7][11] ),
    .S(net191),
    .X(_00960_));
 sky130_fd_sc_hd__mux2_1 _09977_ (.A0(net323),
    .A1(\core_pipeline.pipeline_registers.registers[7][12] ),
    .S(net191),
    .X(_00961_));
 sky130_fd_sc_hd__mux2_1 _09978_ (.A0(net321),
    .A1(\core_pipeline.pipeline_registers.registers[7][13] ),
    .S(net191),
    .X(_00962_));
 sky130_fd_sc_hd__mux2_1 _09979_ (.A0(net320),
    .A1(\core_pipeline.pipeline_registers.registers[7][14] ),
    .S(net191),
    .X(_00963_));
 sky130_fd_sc_hd__mux2_1 _09980_ (.A0(net317),
    .A1(\core_pipeline.pipeline_registers.registers[7][15] ),
    .S(net191),
    .X(_00964_));
 sky130_fd_sc_hd__mux2_1 _09981_ (.A0(net315),
    .A1(\core_pipeline.pipeline_registers.registers[7][16] ),
    .S(net191),
    .X(_00965_));
 sky130_fd_sc_hd__mux2_1 _09982_ (.A0(net314),
    .A1(\core_pipeline.pipeline_registers.registers[7][17] ),
    .S(net192),
    .X(_00966_));
 sky130_fd_sc_hd__mux2_1 _09983_ (.A0(net311),
    .A1(\core_pipeline.pipeline_registers.registers[7][18] ),
    .S(net192),
    .X(_00967_));
 sky130_fd_sc_hd__mux2_1 _09984_ (.A0(net308),
    .A1(\core_pipeline.pipeline_registers.registers[7][19] ),
    .S(net192),
    .X(_00968_));
 sky130_fd_sc_hd__mux2_1 _09985_ (.A0(net305),
    .A1(\core_pipeline.pipeline_registers.registers[7][20] ),
    .S(net192),
    .X(_00969_));
 sky130_fd_sc_hd__mux2_1 _09986_ (.A0(net303),
    .A1(\core_pipeline.pipeline_registers.registers[7][21] ),
    .S(net192),
    .X(_00970_));
 sky130_fd_sc_hd__mux2_1 _09987_ (.A0(net301),
    .A1(\core_pipeline.pipeline_registers.registers[7][22] ),
    .S(net192),
    .X(_00971_));
 sky130_fd_sc_hd__mux2_1 _09988_ (.A0(net300),
    .A1(\core_pipeline.pipeline_registers.registers[7][23] ),
    .S(net192),
    .X(_00972_));
 sky130_fd_sc_hd__mux2_1 _09989_ (.A0(net297),
    .A1(\core_pipeline.pipeline_registers.registers[7][24] ),
    .S(net191),
    .X(_00973_));
 sky130_fd_sc_hd__mux2_1 _09990_ (.A0(net295),
    .A1(\core_pipeline.pipeline_registers.registers[7][25] ),
    .S(net191),
    .X(_00974_));
 sky130_fd_sc_hd__mux2_1 _09991_ (.A0(net294),
    .A1(\core_pipeline.pipeline_registers.registers[7][26] ),
    .S(net191),
    .X(_00975_));
 sky130_fd_sc_hd__mux2_1 _09992_ (.A0(net292),
    .A1(\core_pipeline.pipeline_registers.registers[7][27] ),
    .S(net192),
    .X(_00976_));
 sky130_fd_sc_hd__mux2_1 _09993_ (.A0(net289),
    .A1(\core_pipeline.pipeline_registers.registers[7][28] ),
    .S(net192),
    .X(_00977_));
 sky130_fd_sc_hd__mux2_1 _09994_ (.A0(net288),
    .A1(\core_pipeline.pipeline_registers.registers[7][29] ),
    .S(net192),
    .X(_00978_));
 sky130_fd_sc_hd__mux2_1 _09995_ (.A0(net285),
    .A1(\core_pipeline.pipeline_registers.registers[7][30] ),
    .S(net192),
    .X(_00979_));
 sky130_fd_sc_hd__mux2_1 _09996_ (.A0(net282),
    .A1(\core_pipeline.pipeline_registers.registers[7][31] ),
    .S(net192),
    .X(_00980_));
 sky130_fd_sc_hd__or4_4 _09997_ (.A(\core_pipeline.memory_to_writeback_rd_address[2] ),
    .B(\core_pipeline.memory_to_writeback_rd_address[4] ),
    .C(_04468_),
    .D(_04939_),
    .X(_05603_));
 sky130_fd_sc_hd__mux2_1 _09998_ (.A0(net348),
    .A1(\core_pipeline.pipeline_registers.registers[8][0] ),
    .S(net189),
    .X(_00981_));
 sky130_fd_sc_hd__mux2_1 _09999_ (.A0(net347),
    .A1(\core_pipeline.pipeline_registers.registers[8][1] ),
    .S(net190),
    .X(_00982_));
 sky130_fd_sc_hd__mux2_1 _10000_ (.A0(net344),
    .A1(\core_pipeline.pipeline_registers.registers[8][2] ),
    .S(net190),
    .X(_00983_));
 sky130_fd_sc_hd__mux2_1 _10001_ (.A0(net343),
    .A1(\core_pipeline.pipeline_registers.registers[8][3] ),
    .S(net189),
    .X(_00984_));
 sky130_fd_sc_hd__mux2_1 _10002_ (.A0(net340),
    .A1(\core_pipeline.pipeline_registers.registers[8][4] ),
    .S(net189),
    .X(_00985_));
 sky130_fd_sc_hd__mux2_1 _10003_ (.A0(net337),
    .A1(\core_pipeline.pipeline_registers.registers[8][5] ),
    .S(net190),
    .X(_00986_));
 sky130_fd_sc_hd__mux2_1 _10004_ (.A0(net336),
    .A1(\core_pipeline.pipeline_registers.registers[8][6] ),
    .S(net190),
    .X(_00987_));
 sky130_fd_sc_hd__mux2_1 _10005_ (.A0(net334),
    .A1(\core_pipeline.pipeline_registers.registers[8][7] ),
    .S(net189),
    .X(_00988_));
 sky130_fd_sc_hd__mux2_1 _10006_ (.A0(net332),
    .A1(\core_pipeline.pipeline_registers.registers[8][8] ),
    .S(net189),
    .X(_00989_));
 sky130_fd_sc_hd__mux2_1 _10007_ (.A0(net329),
    .A1(\core_pipeline.pipeline_registers.registers[8][9] ),
    .S(net189),
    .X(_00990_));
 sky130_fd_sc_hd__mux2_1 _10008_ (.A0(net328),
    .A1(\core_pipeline.pipeline_registers.registers[8][10] ),
    .S(net189),
    .X(_00991_));
 sky130_fd_sc_hd__mux2_1 _10009_ (.A0(net325),
    .A1(\core_pipeline.pipeline_registers.registers[8][11] ),
    .S(net189),
    .X(_00992_));
 sky130_fd_sc_hd__mux2_1 _10010_ (.A0(net323),
    .A1(\core_pipeline.pipeline_registers.registers[8][12] ),
    .S(net189),
    .X(_00993_));
 sky130_fd_sc_hd__mux2_1 _10011_ (.A0(net321),
    .A1(\core_pipeline.pipeline_registers.registers[8][13] ),
    .S(net189),
    .X(_00994_));
 sky130_fd_sc_hd__mux2_1 _10012_ (.A0(net320),
    .A1(\core_pipeline.pipeline_registers.registers[8][14] ),
    .S(net189),
    .X(_00995_));
 sky130_fd_sc_hd__mux2_1 _10013_ (.A0(net317),
    .A1(\core_pipeline.pipeline_registers.registers[8][15] ),
    .S(net189),
    .X(_00996_));
 sky130_fd_sc_hd__mux2_1 _10014_ (.A0(net315),
    .A1(\core_pipeline.pipeline_registers.registers[8][16] ),
    .S(net189),
    .X(_00997_));
 sky130_fd_sc_hd__mux2_1 _10015_ (.A0(net312),
    .A1(\core_pipeline.pipeline_registers.registers[8][17] ),
    .S(net190),
    .X(_00998_));
 sky130_fd_sc_hd__mux2_1 _10016_ (.A0(net311),
    .A1(\core_pipeline.pipeline_registers.registers[8][18] ),
    .S(net190),
    .X(_00999_));
 sky130_fd_sc_hd__mux2_1 _10017_ (.A0(net308),
    .A1(\core_pipeline.pipeline_registers.registers[8][19] ),
    .S(net190),
    .X(_01000_));
 sky130_fd_sc_hd__mux2_1 _10018_ (.A0(net306),
    .A1(\core_pipeline.pipeline_registers.registers[8][20] ),
    .S(net190),
    .X(_01001_));
 sky130_fd_sc_hd__mux2_1 _10019_ (.A0(net303),
    .A1(\core_pipeline.pipeline_registers.registers[8][21] ),
    .S(net190),
    .X(_01002_));
 sky130_fd_sc_hd__mux2_1 _10020_ (.A0(net301),
    .A1(\core_pipeline.pipeline_registers.registers[8][22] ),
    .S(net190),
    .X(_01003_));
 sky130_fd_sc_hd__mux2_1 _10021_ (.A0(net300),
    .A1(\core_pipeline.pipeline_registers.registers[8][23] ),
    .S(net190),
    .X(_01004_));
 sky130_fd_sc_hd__mux2_1 _10022_ (.A0(net297),
    .A1(\core_pipeline.pipeline_registers.registers[8][24] ),
    .S(net189),
    .X(_01005_));
 sky130_fd_sc_hd__mux2_1 _10023_ (.A0(net295),
    .A1(\core_pipeline.pipeline_registers.registers[8][25] ),
    .S(net189),
    .X(_01006_));
 sky130_fd_sc_hd__mux2_1 _10024_ (.A0(net293),
    .A1(\core_pipeline.pipeline_registers.registers[8][26] ),
    .S(net189),
    .X(_01007_));
 sky130_fd_sc_hd__mux2_1 _10025_ (.A0(net292),
    .A1(\core_pipeline.pipeline_registers.registers[8][27] ),
    .S(net190),
    .X(_01008_));
 sky130_fd_sc_hd__mux2_1 _10026_ (.A0(net289),
    .A1(\core_pipeline.pipeline_registers.registers[8][28] ),
    .S(net190),
    .X(_01009_));
 sky130_fd_sc_hd__mux2_1 _10027_ (.A0(net287),
    .A1(\core_pipeline.pipeline_registers.registers[8][29] ),
    .S(net190),
    .X(_01010_));
 sky130_fd_sc_hd__mux2_1 _10028_ (.A0(net284),
    .A1(\core_pipeline.pipeline_registers.registers[8][30] ),
    .S(net189),
    .X(_01011_));
 sky130_fd_sc_hd__mux2_1 _10029_ (.A0(net283),
    .A1(\core_pipeline.pipeline_registers.registers[8][31] ),
    .S(net190),
    .X(_01012_));
 sky130_fd_sc_hd__a32o_1 _10030_ (.A1(net638),
    .A2(\core_pipeline.csr_to_fetch_mret_vector[0] ),
    .A3(_04385_),
    .B1(_03517_),
    .B2(\core_pipeline.pipeline_fetch.pc[0] ),
    .X(_01013_));
 sky130_fd_sc_hd__a32o_1 _10031_ (.A1(net638),
    .A2(\core_pipeline.csr_to_fetch_mret_vector[1] ),
    .A3(_04385_),
    .B1(_03517_),
    .B2(\core_pipeline.pipeline_fetch.pc[1] ),
    .X(_01014_));
 sky130_fd_sc_hd__nor2_8 _10032_ (.A(_04469_),
    .B(_05589_),
    .Y(_05604_));
 sky130_fd_sc_hd__mux2_1 _10033_ (.A0(\core_pipeline.pipeline_registers.registers[29][0] ),
    .A1(net349),
    .S(net187),
    .X(_01015_));
 sky130_fd_sc_hd__mux2_1 _10034_ (.A0(\core_pipeline.pipeline_registers.registers[29][1] ),
    .A1(net346),
    .S(net188),
    .X(_01016_));
 sky130_fd_sc_hd__mux2_1 _10035_ (.A0(\core_pipeline.pipeline_registers.registers[29][2] ),
    .A1(net344),
    .S(net188),
    .X(_01017_));
 sky130_fd_sc_hd__mux2_1 _10036_ (.A0(\core_pipeline.pipeline_registers.registers[29][3] ),
    .A1(net342),
    .S(net187),
    .X(_01018_));
 sky130_fd_sc_hd__mux2_1 _10037_ (.A0(\core_pipeline.pipeline_registers.registers[29][4] ),
    .A1(net341),
    .S(net187),
    .X(_01019_));
 sky130_fd_sc_hd__mux2_1 _10038_ (.A0(\core_pipeline.pipeline_registers.registers[29][5] ),
    .A1(net338),
    .S(net188),
    .X(_01020_));
 sky130_fd_sc_hd__mux2_1 _10039_ (.A0(\core_pipeline.pipeline_registers.registers[29][6] ),
    .A1(net335),
    .S(net188),
    .X(_01021_));
 sky130_fd_sc_hd__mux2_1 _10040_ (.A0(\core_pipeline.pipeline_registers.registers[29][7] ),
    .A1(net333),
    .S(net187),
    .X(_01022_));
 sky130_fd_sc_hd__mux2_1 _10041_ (.A0(\core_pipeline.pipeline_registers.registers[29][8] ),
    .A1(net331),
    .S(net187),
    .X(_01023_));
 sky130_fd_sc_hd__mux2_1 _10042_ (.A0(\core_pipeline.pipeline_registers.registers[29][9] ),
    .A1(net330),
    .S(net187),
    .X(_01024_));
 sky130_fd_sc_hd__mux2_1 _10043_ (.A0(\core_pipeline.pipeline_registers.registers[29][10] ),
    .A1(net328),
    .S(net187),
    .X(_01025_));
 sky130_fd_sc_hd__mux2_1 _10044_ (.A0(\core_pipeline.pipeline_registers.registers[29][11] ),
    .A1(net326),
    .S(net187),
    .X(_01026_));
 sky130_fd_sc_hd__mux2_1 _10045_ (.A0(\core_pipeline.pipeline_registers.registers[29][12] ),
    .A1(net324),
    .S(net187),
    .X(_01027_));
 sky130_fd_sc_hd__mux2_1 _10046_ (.A0(\core_pipeline.pipeline_registers.registers[29][13] ),
    .A1(net322),
    .S(net187),
    .X(_01028_));
 sky130_fd_sc_hd__mux2_1 _10047_ (.A0(\core_pipeline.pipeline_registers.registers[29][14] ),
    .A1(net319),
    .S(net187),
    .X(_01029_));
 sky130_fd_sc_hd__mux2_1 _10048_ (.A0(\core_pipeline.pipeline_registers.registers[29][15] ),
    .A1(net318),
    .S(net187),
    .X(_01030_));
 sky130_fd_sc_hd__mux2_1 _10049_ (.A0(\core_pipeline.pipeline_registers.registers[29][16] ),
    .A1(net315),
    .S(net187),
    .X(_01031_));
 sky130_fd_sc_hd__mux2_1 _10050_ (.A0(\core_pipeline.pipeline_registers.registers[29][17] ),
    .A1(net312),
    .S(net188),
    .X(_01032_));
 sky130_fd_sc_hd__mux2_1 _10051_ (.A0(\core_pipeline.pipeline_registers.registers[29][18] ),
    .A1(net310),
    .S(net188),
    .X(_01033_));
 sky130_fd_sc_hd__mux2_1 _10052_ (.A0(\core_pipeline.pipeline_registers.registers[29][19] ),
    .A1(net309),
    .S(net188),
    .X(_01034_));
 sky130_fd_sc_hd__mux2_1 _10053_ (.A0(\core_pipeline.pipeline_registers.registers[29][20] ),
    .A1(net305),
    .S(net188),
    .X(_01035_));
 sky130_fd_sc_hd__mux2_1 _10054_ (.A0(\core_pipeline.pipeline_registers.registers[29][21] ),
    .A1(net303),
    .S(net188),
    .X(_01036_));
 sky130_fd_sc_hd__mux2_1 _10055_ (.A0(\core_pipeline.pipeline_registers.registers[29][22] ),
    .A1(net302),
    .S(net187),
    .X(_01037_));
 sky130_fd_sc_hd__mux2_1 _10056_ (.A0(\core_pipeline.pipeline_registers.registers[29][23] ),
    .A1(net300),
    .S(net188),
    .X(_01038_));
 sky130_fd_sc_hd__mux2_1 _10057_ (.A0(\core_pipeline.pipeline_registers.registers[29][24] ),
    .A1(net298),
    .S(net187),
    .X(_01039_));
 sky130_fd_sc_hd__mux2_1 _10058_ (.A0(\core_pipeline.pipeline_registers.registers[29][25] ),
    .A1(net296),
    .S(net187),
    .X(_01040_));
 sky130_fd_sc_hd__mux2_1 _10059_ (.A0(\core_pipeline.pipeline_registers.registers[29][26] ),
    .A1(net294),
    .S(net187),
    .X(_01041_));
 sky130_fd_sc_hd__mux2_1 _10060_ (.A0(\core_pipeline.pipeline_registers.registers[29][27] ),
    .A1(net291),
    .S(net188),
    .X(_01042_));
 sky130_fd_sc_hd__mux2_1 _10061_ (.A0(\core_pipeline.pipeline_registers.registers[29][28] ),
    .A1(net290),
    .S(net188),
    .X(_01043_));
 sky130_fd_sc_hd__mux2_1 _10062_ (.A0(\core_pipeline.pipeline_registers.registers[29][29] ),
    .A1(net286),
    .S(net188),
    .X(_01044_));
 sky130_fd_sc_hd__mux2_1 _10063_ (.A0(\core_pipeline.pipeline_registers.registers[29][30] ),
    .A1(net284),
    .S(net188),
    .X(_01045_));
 sky130_fd_sc_hd__mux2_1 _10064_ (.A0(\core_pipeline.pipeline_registers.registers[29][31] ),
    .A1(net282),
    .S(net188),
    .X(_01046_));
 sky130_fd_sc_hd__nor2_8 _10065_ (.A(_04937_),
    .B(_05589_),
    .Y(_05605_));
 sky130_fd_sc_hd__mux2_1 _10066_ (.A0(\core_pipeline.pipeline_registers.registers[1][0] ),
    .A1(net348),
    .S(net185),
    .X(_01047_));
 sky130_fd_sc_hd__mux2_1 _10067_ (.A0(\core_pipeline.pipeline_registers.registers[1][1] ),
    .A1(net347),
    .S(net186),
    .X(_01048_));
 sky130_fd_sc_hd__mux2_1 _10068_ (.A0(\core_pipeline.pipeline_registers.registers[1][2] ),
    .A1(net345),
    .S(net186),
    .X(_01049_));
 sky130_fd_sc_hd__mux2_1 _10069_ (.A0(\core_pipeline.pipeline_registers.registers[1][3] ),
    .A1(net342),
    .S(net185),
    .X(_01050_));
 sky130_fd_sc_hd__mux2_1 _10070_ (.A0(\core_pipeline.pipeline_registers.registers[1][4] ),
    .A1(net340),
    .S(net185),
    .X(_01051_));
 sky130_fd_sc_hd__mux2_1 _10071_ (.A0(\core_pipeline.pipeline_registers.registers[1][5] ),
    .A1(net338),
    .S(net186),
    .X(_01052_));
 sky130_fd_sc_hd__mux2_1 _10072_ (.A0(\core_pipeline.pipeline_registers.registers[1][6] ),
    .A1(net335),
    .S(net185),
    .X(_01053_));
 sky130_fd_sc_hd__mux2_1 _10073_ (.A0(\core_pipeline.pipeline_registers.registers[1][7] ),
    .A1(net334),
    .S(net185),
    .X(_01054_));
 sky130_fd_sc_hd__mux2_1 _10074_ (.A0(\core_pipeline.pipeline_registers.registers[1][8] ),
    .A1(net332),
    .S(net185),
    .X(_01055_));
 sky130_fd_sc_hd__mux2_1 _10075_ (.A0(\core_pipeline.pipeline_registers.registers[1][9] ),
    .A1(net329),
    .S(net185),
    .X(_01056_));
 sky130_fd_sc_hd__mux2_1 _10076_ (.A0(\core_pipeline.pipeline_registers.registers[1][10] ),
    .A1(net327),
    .S(net185),
    .X(_01057_));
 sky130_fd_sc_hd__mux2_1 _10077_ (.A0(\core_pipeline.pipeline_registers.registers[1][11] ),
    .A1(net325),
    .S(net185),
    .X(_01058_));
 sky130_fd_sc_hd__mux2_1 _10078_ (.A0(\core_pipeline.pipeline_registers.registers[1][12] ),
    .A1(net324),
    .S(net185),
    .X(_01059_));
 sky130_fd_sc_hd__mux2_1 _10079_ (.A0(\core_pipeline.pipeline_registers.registers[1][13] ),
    .A1(net322),
    .S(net185),
    .X(_01060_));
 sky130_fd_sc_hd__mux2_1 _10080_ (.A0(\core_pipeline.pipeline_registers.registers[1][14] ),
    .A1(net320),
    .S(net185),
    .X(_01061_));
 sky130_fd_sc_hd__mux2_1 _10081_ (.A0(\core_pipeline.pipeline_registers.registers[1][15] ),
    .A1(net317),
    .S(net185),
    .X(_01062_));
 sky130_fd_sc_hd__mux2_1 _10082_ (.A0(\core_pipeline.pipeline_registers.registers[1][16] ),
    .A1(net315),
    .S(net185),
    .X(_01063_));
 sky130_fd_sc_hd__mux2_1 _10083_ (.A0(\core_pipeline.pipeline_registers.registers[1][17] ),
    .A1(net313),
    .S(net186),
    .X(_01064_));
 sky130_fd_sc_hd__mux2_1 _10084_ (.A0(\core_pipeline.pipeline_registers.registers[1][18] ),
    .A1(net311),
    .S(net186),
    .X(_01065_));
 sky130_fd_sc_hd__mux2_1 _10085_ (.A0(\core_pipeline.pipeline_registers.registers[1][19] ),
    .A1(net308),
    .S(net186),
    .X(_01066_));
 sky130_fd_sc_hd__mux2_1 _10086_ (.A0(\core_pipeline.pipeline_registers.registers[1][20] ),
    .A1(net305),
    .S(net186),
    .X(_01067_));
 sky130_fd_sc_hd__mux2_1 _10087_ (.A0(\core_pipeline.pipeline_registers.registers[1][21] ),
    .A1(net304),
    .S(net186),
    .X(_01068_));
 sky130_fd_sc_hd__mux2_1 _10088_ (.A0(\core_pipeline.pipeline_registers.registers[1][22] ),
    .A1(net301),
    .S(net186),
    .X(_01069_));
 sky130_fd_sc_hd__mux2_1 _10089_ (.A0(\core_pipeline.pipeline_registers.registers[1][23] ),
    .A1(net300),
    .S(net186),
    .X(_01070_));
 sky130_fd_sc_hd__mux2_1 _10090_ (.A0(\core_pipeline.pipeline_registers.registers[1][24] ),
    .A1(net298),
    .S(net185),
    .X(_01071_));
 sky130_fd_sc_hd__mux2_1 _10091_ (.A0(\core_pipeline.pipeline_registers.registers[1][25] ),
    .A1(net295),
    .S(net185),
    .X(_01072_));
 sky130_fd_sc_hd__mux2_1 _10092_ (.A0(\core_pipeline.pipeline_registers.registers[1][26] ),
    .A1(net293),
    .S(net185),
    .X(_01073_));
 sky130_fd_sc_hd__mux2_1 _10093_ (.A0(\core_pipeline.pipeline_registers.registers[1][27] ),
    .A1(net292),
    .S(net186),
    .X(_01074_));
 sky130_fd_sc_hd__mux2_1 _10094_ (.A0(\core_pipeline.pipeline_registers.registers[1][28] ),
    .A1(net290),
    .S(net186),
    .X(_01075_));
 sky130_fd_sc_hd__mux2_1 _10095_ (.A0(\core_pipeline.pipeline_registers.registers[1][29] ),
    .A1(net288),
    .S(net186),
    .X(_01076_));
 sky130_fd_sc_hd__mux2_1 _10096_ (.A0(\core_pipeline.pipeline_registers.registers[1][30] ),
    .A1(net285),
    .S(net186),
    .X(_01077_));
 sky130_fd_sc_hd__mux2_1 _10097_ (.A0(\core_pipeline.pipeline_registers.registers[1][31] ),
    .A1(net283),
    .S(net186),
    .X(_01078_));
 sky130_fd_sc_hd__nor2_1 _10098_ (.A(_03644_),
    .B(_04110_),
    .Y(_05606_));
 sky130_fd_sc_hd__and3_4 _10099_ (.A(\core_pipeline.memory_to_writeback_csr_address[0] ),
    .B(_03647_),
    .C(_05606_),
    .X(_05607_));
 sky130_fd_sc_hd__mux2_1 _10100_ (.A0(\core_pipeline.pipeline_csr.mtimecmp[32] ),
    .A1(\core_pipeline.memory_to_writeback_alu_data[0] ),
    .S(net183),
    .X(_01111_));
 sky130_fd_sc_hd__mux2_1 _10101_ (.A0(\core_pipeline.pipeline_csr.mtimecmp[33] ),
    .A1(\core_pipeline.memory_to_writeback_alu_data[1] ),
    .S(net183),
    .X(_01112_));
 sky130_fd_sc_hd__mux2_1 _10102_ (.A0(\core_pipeline.pipeline_csr.mtimecmp[34] ),
    .A1(\core_pipeline.memory_to_writeback_alu_data[2] ),
    .S(net183),
    .X(_01113_));
 sky130_fd_sc_hd__mux2_1 _10103_ (.A0(\core_pipeline.pipeline_csr.mtimecmp[35] ),
    .A1(\core_pipeline.memory_to_writeback_alu_data[3] ),
    .S(net183),
    .X(_01114_));
 sky130_fd_sc_hd__mux2_1 _10104_ (.A0(\core_pipeline.pipeline_csr.mtimecmp[36] ),
    .A1(\core_pipeline.memory_to_writeback_alu_data[4] ),
    .S(net183),
    .X(_01115_));
 sky130_fd_sc_hd__mux2_1 _10105_ (.A0(\core_pipeline.pipeline_csr.mtimecmp[37] ),
    .A1(\core_pipeline.memory_to_writeback_alu_data[5] ),
    .S(net183),
    .X(_01116_));
 sky130_fd_sc_hd__mux2_1 _10106_ (.A0(\core_pipeline.pipeline_csr.mtimecmp[38] ),
    .A1(\core_pipeline.memory_to_writeback_alu_data[6] ),
    .S(net183),
    .X(_01117_));
 sky130_fd_sc_hd__mux2_1 _10107_ (.A0(\core_pipeline.pipeline_csr.mtimecmp[39] ),
    .A1(\core_pipeline.memory_to_writeback_alu_data[7] ),
    .S(net183),
    .X(_01118_));
 sky130_fd_sc_hd__mux2_1 _10108_ (.A0(\core_pipeline.pipeline_csr.mtimecmp[40] ),
    .A1(\core_pipeline.memory_to_writeback_alu_data[8] ),
    .S(net184),
    .X(_01119_));
 sky130_fd_sc_hd__mux2_1 _10109_ (.A0(\core_pipeline.pipeline_csr.mtimecmp[41] ),
    .A1(\core_pipeline.memory_to_writeback_alu_data[9] ),
    .S(net184),
    .X(_01120_));
 sky130_fd_sc_hd__mux2_1 _10110_ (.A0(\core_pipeline.pipeline_csr.mtimecmp[42] ),
    .A1(\core_pipeline.memory_to_writeback_alu_data[10] ),
    .S(net184),
    .X(_01121_));
 sky130_fd_sc_hd__mux2_1 _10111_ (.A0(\core_pipeline.pipeline_csr.mtimecmp[43] ),
    .A1(\core_pipeline.memory_to_writeback_alu_data[11] ),
    .S(net183),
    .X(_01122_));
 sky130_fd_sc_hd__mux2_1 _10112_ (.A0(\core_pipeline.pipeline_csr.mtimecmp[44] ),
    .A1(\core_pipeline.memory_to_writeback_alu_data[12] ),
    .S(net184),
    .X(_01123_));
 sky130_fd_sc_hd__mux2_1 _10113_ (.A0(\core_pipeline.pipeline_csr.mtimecmp[45] ),
    .A1(\core_pipeline.memory_to_writeback_alu_data[13] ),
    .S(net184),
    .X(_01124_));
 sky130_fd_sc_hd__mux2_1 _10114_ (.A0(\core_pipeline.pipeline_csr.mtimecmp[46] ),
    .A1(\core_pipeline.memory_to_writeback_alu_data[14] ),
    .S(net184),
    .X(_01125_));
 sky130_fd_sc_hd__mux2_1 _10115_ (.A0(\core_pipeline.pipeline_csr.mtimecmp[47] ),
    .A1(\core_pipeline.memory_to_writeback_alu_data[15] ),
    .S(net184),
    .X(_01126_));
 sky130_fd_sc_hd__mux2_1 _10116_ (.A0(\core_pipeline.pipeline_csr.mtimecmp[48] ),
    .A1(\core_pipeline.memory_to_writeback_alu_data[16] ),
    .S(net184),
    .X(_01127_));
 sky130_fd_sc_hd__mux2_1 _10117_ (.A0(\core_pipeline.pipeline_csr.mtimecmp[49] ),
    .A1(\core_pipeline.memory_to_writeback_alu_data[17] ),
    .S(net184),
    .X(_01128_));
 sky130_fd_sc_hd__mux2_1 _10118_ (.A0(\core_pipeline.pipeline_csr.mtimecmp[50] ),
    .A1(\core_pipeline.memory_to_writeback_alu_data[18] ),
    .S(net184),
    .X(_01129_));
 sky130_fd_sc_hd__mux2_1 _10119_ (.A0(\core_pipeline.pipeline_csr.mtimecmp[51] ),
    .A1(\core_pipeline.memory_to_writeback_alu_data[19] ),
    .S(net183),
    .X(_01130_));
 sky130_fd_sc_hd__mux2_1 _10120_ (.A0(\core_pipeline.pipeline_csr.mtimecmp[52] ),
    .A1(\core_pipeline.memory_to_writeback_alu_data[20] ),
    .S(net184),
    .X(_01131_));
 sky130_fd_sc_hd__mux2_1 _10121_ (.A0(\core_pipeline.pipeline_csr.mtimecmp[53] ),
    .A1(\core_pipeline.memory_to_writeback_alu_data[21] ),
    .S(net184),
    .X(_01132_));
 sky130_fd_sc_hd__mux2_1 _10122_ (.A0(\core_pipeline.pipeline_csr.mtimecmp[54] ),
    .A1(\core_pipeline.memory_to_writeback_alu_data[22] ),
    .S(net184),
    .X(_01133_));
 sky130_fd_sc_hd__mux2_1 _10123_ (.A0(\core_pipeline.pipeline_csr.mtimecmp[55] ),
    .A1(\core_pipeline.memory_to_writeback_alu_data[23] ),
    .S(net184),
    .X(_01134_));
 sky130_fd_sc_hd__mux2_1 _10124_ (.A0(\core_pipeline.pipeline_csr.mtimecmp[56] ),
    .A1(\core_pipeline.memory_to_writeback_alu_data[24] ),
    .S(net184),
    .X(_01135_));
 sky130_fd_sc_hd__mux2_1 _10125_ (.A0(\core_pipeline.pipeline_csr.mtimecmp[57] ),
    .A1(\core_pipeline.memory_to_writeback_alu_data[25] ),
    .S(net183),
    .X(_01136_));
 sky130_fd_sc_hd__mux2_1 _10126_ (.A0(\core_pipeline.pipeline_csr.mtimecmp[58] ),
    .A1(\core_pipeline.memory_to_writeback_alu_data[26] ),
    .S(net183),
    .X(_01137_));
 sky130_fd_sc_hd__mux2_1 _10127_ (.A0(\core_pipeline.pipeline_csr.mtimecmp[59] ),
    .A1(\core_pipeline.memory_to_writeback_alu_data[27] ),
    .S(net183),
    .X(_01138_));
 sky130_fd_sc_hd__mux2_1 _10128_ (.A0(\core_pipeline.pipeline_csr.mtimecmp[60] ),
    .A1(\core_pipeline.memory_to_writeback_alu_data[28] ),
    .S(net183),
    .X(_01139_));
 sky130_fd_sc_hd__mux2_1 _10129_ (.A0(\core_pipeline.pipeline_csr.mtimecmp[61] ),
    .A1(\core_pipeline.memory_to_writeback_alu_data[29] ),
    .S(net183),
    .X(_01140_));
 sky130_fd_sc_hd__mux2_1 _10130_ (.A0(\core_pipeline.pipeline_csr.mtimecmp[62] ),
    .A1(\core_pipeline.memory_to_writeback_alu_data[30] ),
    .S(net183),
    .X(_01141_));
 sky130_fd_sc_hd__mux2_1 _10131_ (.A0(\core_pipeline.pipeline_csr.mtimecmp[63] ),
    .A1(\core_pipeline.memory_to_writeback_alu_data[31] ),
    .S(net183),
    .X(_01142_));
 sky130_fd_sc_hd__nor2_8 _10132_ (.A(_04939_),
    .B(_05592_),
    .Y(_05608_));
 sky130_fd_sc_hd__mux2_1 _10133_ (.A0(\core_pipeline.pipeline_registers.registers[20][0] ),
    .A1(net348),
    .S(net181),
    .X(_01143_));
 sky130_fd_sc_hd__mux2_1 _10134_ (.A0(\core_pipeline.pipeline_registers.registers[20][1] ),
    .A1(net347),
    .S(net182),
    .X(_01144_));
 sky130_fd_sc_hd__mux2_1 _10135_ (.A0(\core_pipeline.pipeline_registers.registers[20][2] ),
    .A1(net345),
    .S(net182),
    .X(_01145_));
 sky130_fd_sc_hd__mux2_1 _10136_ (.A0(\core_pipeline.pipeline_registers.registers[20][3] ),
    .A1(net342),
    .S(net181),
    .X(_01146_));
 sky130_fd_sc_hd__mux2_1 _10137_ (.A0(\core_pipeline.pipeline_registers.registers[20][4] ),
    .A1(net341),
    .S(net181),
    .X(_01147_));
 sky130_fd_sc_hd__mux2_1 _10138_ (.A0(\core_pipeline.pipeline_registers.registers[20][5] ),
    .A1(net338),
    .S(net182),
    .X(_01148_));
 sky130_fd_sc_hd__mux2_1 _10139_ (.A0(\core_pipeline.pipeline_registers.registers[20][6] ),
    .A1(net336),
    .S(net181),
    .X(_01149_));
 sky130_fd_sc_hd__mux2_1 _10140_ (.A0(\core_pipeline.pipeline_registers.registers[20][7] ),
    .A1(net333),
    .S(net181),
    .X(_01150_));
 sky130_fd_sc_hd__mux2_1 _10141_ (.A0(\core_pipeline.pipeline_registers.registers[20][8] ),
    .A1(net331),
    .S(net181),
    .X(_01151_));
 sky130_fd_sc_hd__mux2_1 _10142_ (.A0(\core_pipeline.pipeline_registers.registers[20][9] ),
    .A1(net330),
    .S(net181),
    .X(_01152_));
 sky130_fd_sc_hd__mux2_1 _10143_ (.A0(\core_pipeline.pipeline_registers.registers[20][10] ),
    .A1(net327),
    .S(net181),
    .X(_01153_));
 sky130_fd_sc_hd__mux2_1 _10144_ (.A0(\core_pipeline.pipeline_registers.registers[20][11] ),
    .A1(net326),
    .S(net181),
    .X(_01154_));
 sky130_fd_sc_hd__mux2_1 _10145_ (.A0(\core_pipeline.pipeline_registers.registers[20][12] ),
    .A1(net324),
    .S(net181),
    .X(_01155_));
 sky130_fd_sc_hd__mux2_1 _10146_ (.A0(\core_pipeline.pipeline_registers.registers[20][13] ),
    .A1(net321),
    .S(net181),
    .X(_01156_));
 sky130_fd_sc_hd__mux2_1 _10147_ (.A0(\core_pipeline.pipeline_registers.registers[20][14] ),
    .A1(net319),
    .S(net181),
    .X(_01157_));
 sky130_fd_sc_hd__mux2_1 _10148_ (.A0(\core_pipeline.pipeline_registers.registers[20][15] ),
    .A1(net318),
    .S(net181),
    .X(_01158_));
 sky130_fd_sc_hd__mux2_1 _10149_ (.A0(\core_pipeline.pipeline_registers.registers[20][16] ),
    .A1(net316),
    .S(net181),
    .X(_01159_));
 sky130_fd_sc_hd__mux2_1 _10150_ (.A0(\core_pipeline.pipeline_registers.registers[20][17] ),
    .A1(net314),
    .S(net182),
    .X(_01160_));
 sky130_fd_sc_hd__mux2_1 _10151_ (.A0(\core_pipeline.pipeline_registers.registers[20][18] ),
    .A1(net310),
    .S(net182),
    .X(_01161_));
 sky130_fd_sc_hd__mux2_1 _10152_ (.A0(\core_pipeline.pipeline_registers.registers[20][19] ),
    .A1(net308),
    .S(net182),
    .X(_01162_));
 sky130_fd_sc_hd__mux2_1 _10153_ (.A0(\core_pipeline.pipeline_registers.registers[20][20] ),
    .A1(net306),
    .S(net182),
    .X(_01163_));
 sky130_fd_sc_hd__mux2_1 _10154_ (.A0(\core_pipeline.pipeline_registers.registers[20][21] ),
    .A1(net304),
    .S(net182),
    .X(_01164_));
 sky130_fd_sc_hd__mux2_1 _10155_ (.A0(\core_pipeline.pipeline_registers.registers[20][22] ),
    .A1(net302),
    .S(net182),
    .X(_01165_));
 sky130_fd_sc_hd__mux2_1 _10156_ (.A0(\core_pipeline.pipeline_registers.registers[20][23] ),
    .A1(net299),
    .S(net182),
    .X(_01166_));
 sky130_fd_sc_hd__mux2_1 _10157_ (.A0(\core_pipeline.pipeline_registers.registers[20][24] ),
    .A1(net297),
    .S(net181),
    .X(_01167_));
 sky130_fd_sc_hd__mux2_1 _10158_ (.A0(\core_pipeline.pipeline_registers.registers[20][25] ),
    .A1(net295),
    .S(net181),
    .X(_01168_));
 sky130_fd_sc_hd__mux2_1 _10159_ (.A0(\core_pipeline.pipeline_registers.registers[20][26] ),
    .A1(net293),
    .S(net181),
    .X(_01169_));
 sky130_fd_sc_hd__mux2_1 _10160_ (.A0(\core_pipeline.pipeline_registers.registers[20][27] ),
    .A1(net291),
    .S(net182),
    .X(_01170_));
 sky130_fd_sc_hd__mux2_1 _10161_ (.A0(\core_pipeline.pipeline_registers.registers[20][28] ),
    .A1(net290),
    .S(net182),
    .X(_01171_));
 sky130_fd_sc_hd__mux2_1 _10162_ (.A0(\core_pipeline.pipeline_registers.registers[20][29] ),
    .A1(net286),
    .S(net182),
    .X(_01172_));
 sky130_fd_sc_hd__mux2_1 _10163_ (.A0(\core_pipeline.pipeline_registers.registers[20][30] ),
    .A1(net285),
    .S(net182),
    .X(_01173_));
 sky130_fd_sc_hd__mux2_1 _10164_ (.A0(\core_pipeline.pipeline_registers.registers[20][31] ),
    .A1(net283),
    .S(net182),
    .X(_01174_));
 sky130_fd_sc_hd__or4_4 _10165_ (.A(\core_pipeline.memory_to_writeback_rd_address[2] ),
    .B(\core_pipeline.memory_to_writeback_rd_address[4] ),
    .C(_03915_),
    .D(_04468_),
    .X(_05609_));
 sky130_fd_sc_hd__mux2_1 _10166_ (.A0(net348),
    .A1(\core_pipeline.pipeline_registers.registers[11][0] ),
    .S(net241),
    .X(_01175_));
 sky130_fd_sc_hd__mux2_1 _10167_ (.A0(net346),
    .A1(\core_pipeline.pipeline_registers.registers[11][1] ),
    .S(net242),
    .X(_01176_));
 sky130_fd_sc_hd__mux2_1 _10168_ (.A0(net344),
    .A1(\core_pipeline.pipeline_registers.registers[11][2] ),
    .S(net242),
    .X(_01177_));
 sky130_fd_sc_hd__mux2_1 _10169_ (.A0(net343),
    .A1(\core_pipeline.pipeline_registers.registers[11][3] ),
    .S(net241),
    .X(_01178_));
 sky130_fd_sc_hd__mux2_1 _10170_ (.A0(net340),
    .A1(\core_pipeline.pipeline_registers.registers[11][4] ),
    .S(net241),
    .X(_01179_));
 sky130_fd_sc_hd__mux2_1 _10171_ (.A0(net337),
    .A1(\core_pipeline.pipeline_registers.registers[11][5] ),
    .S(net242),
    .X(_01180_));
 sky130_fd_sc_hd__mux2_1 _10172_ (.A0(net335),
    .A1(\core_pipeline.pipeline_registers.registers[11][6] ),
    .S(net241),
    .X(_01181_));
 sky130_fd_sc_hd__mux2_1 _10173_ (.A0(net334),
    .A1(\core_pipeline.pipeline_registers.registers[11][7] ),
    .S(net241),
    .X(_01182_));
 sky130_fd_sc_hd__mux2_1 _10174_ (.A0(net332),
    .A1(\core_pipeline.pipeline_registers.registers[11][8] ),
    .S(net241),
    .X(_01183_));
 sky130_fd_sc_hd__mux2_1 _10175_ (.A0(net329),
    .A1(\core_pipeline.pipeline_registers.registers[11][9] ),
    .S(net241),
    .X(_01184_));
 sky130_fd_sc_hd__mux2_1 _10176_ (.A0(net327),
    .A1(\core_pipeline.pipeline_registers.registers[11][10] ),
    .S(net241),
    .X(_01185_));
 sky130_fd_sc_hd__mux2_1 _10177_ (.A0(net325),
    .A1(\core_pipeline.pipeline_registers.registers[11][11] ),
    .S(net241),
    .X(_01186_));
 sky130_fd_sc_hd__mux2_1 _10178_ (.A0(net323),
    .A1(\core_pipeline.pipeline_registers.registers[11][12] ),
    .S(net241),
    .X(_01187_));
 sky130_fd_sc_hd__mux2_1 _10179_ (.A0(net321),
    .A1(\core_pipeline.pipeline_registers.registers[11][13] ),
    .S(net241),
    .X(_01188_));
 sky130_fd_sc_hd__mux2_1 _10180_ (.A0(net320),
    .A1(\core_pipeline.pipeline_registers.registers[11][14] ),
    .S(net241),
    .X(_01189_));
 sky130_fd_sc_hd__mux2_1 _10181_ (.A0(net317),
    .A1(\core_pipeline.pipeline_registers.registers[11][15] ),
    .S(net241),
    .X(_01190_));
 sky130_fd_sc_hd__mux2_1 _10182_ (.A0(net315),
    .A1(\core_pipeline.pipeline_registers.registers[11][16] ),
    .S(net241),
    .X(_01191_));
 sky130_fd_sc_hd__mux2_1 _10183_ (.A0(net312),
    .A1(\core_pipeline.pipeline_registers.registers[11][17] ),
    .S(net242),
    .X(_01192_));
 sky130_fd_sc_hd__mux2_1 _10184_ (.A0(net311),
    .A1(\core_pipeline.pipeline_registers.registers[11][18] ),
    .S(net242),
    .X(_01193_));
 sky130_fd_sc_hd__mux2_1 _10185_ (.A0(net308),
    .A1(\core_pipeline.pipeline_registers.registers[11][19] ),
    .S(net242),
    .X(_01194_));
 sky130_fd_sc_hd__mux2_1 _10186_ (.A0(net305),
    .A1(\core_pipeline.pipeline_registers.registers[11][20] ),
    .S(net242),
    .X(_01195_));
 sky130_fd_sc_hd__mux2_1 _10187_ (.A0(net303),
    .A1(\core_pipeline.pipeline_registers.registers[11][21] ),
    .S(net242),
    .X(_01196_));
 sky130_fd_sc_hd__mux2_1 _10188_ (.A0(net301),
    .A1(\core_pipeline.pipeline_registers.registers[11][22] ),
    .S(net242),
    .X(_01197_));
 sky130_fd_sc_hd__mux2_1 _10189_ (.A0(net300),
    .A1(\core_pipeline.pipeline_registers.registers[11][23] ),
    .S(net242),
    .X(_01198_));
 sky130_fd_sc_hd__mux2_1 _10190_ (.A0(net297),
    .A1(\core_pipeline.pipeline_registers.registers[11][24] ),
    .S(net241),
    .X(_01199_));
 sky130_fd_sc_hd__mux2_1 _10191_ (.A0(net295),
    .A1(\core_pipeline.pipeline_registers.registers[11][25] ),
    .S(net241),
    .X(_01200_));
 sky130_fd_sc_hd__mux2_1 _10192_ (.A0(net293),
    .A1(\core_pipeline.pipeline_registers.registers[11][26] ),
    .S(net241),
    .X(_01201_));
 sky130_fd_sc_hd__mux2_1 _10193_ (.A0(net292),
    .A1(\core_pipeline.pipeline_registers.registers[11][27] ),
    .S(net242),
    .X(_01202_));
 sky130_fd_sc_hd__mux2_1 _10194_ (.A0(net289),
    .A1(\core_pipeline.pipeline_registers.registers[11][28] ),
    .S(net242),
    .X(_01203_));
 sky130_fd_sc_hd__mux2_1 _10195_ (.A0(net286),
    .A1(\core_pipeline.pipeline_registers.registers[11][29] ),
    .S(net242),
    .X(_01204_));
 sky130_fd_sc_hd__mux2_1 _10196_ (.A0(net284),
    .A1(\core_pipeline.pipeline_registers.registers[11][30] ),
    .S(net242),
    .X(_01205_));
 sky130_fd_sc_hd__mux2_1 _10197_ (.A0(net282),
    .A1(\core_pipeline.pipeline_registers.registers[11][31] ),
    .S(net242),
    .X(_01206_));
 sky130_fd_sc_hd__mux2_1 _10198_ (.A0(net1),
    .A1(\core_pipeline.fetch_to_decode_instruction[0] ),
    .S(net107),
    .X(_01207_));
 sky130_fd_sc_hd__mux2_1 _10199_ (.A0(net12),
    .A1(\core_pipeline.fetch_to_decode_instruction[1] ),
    .S(net107),
    .X(_01208_));
 sky130_fd_sc_hd__mux2_1 _10200_ (.A0(net23),
    .A1(\core_pipeline.fetch_to_decode_instruction[2] ),
    .S(net107),
    .X(_01209_));
 sky130_fd_sc_hd__mux2_1 _10201_ (.A0(net26),
    .A1(\core_pipeline.fetch_to_decode_instruction[3] ),
    .S(net107),
    .X(_01210_));
 sky130_fd_sc_hd__mux2_1 _10202_ (.A0(net27),
    .A1(\core_pipeline.fetch_to_decode_instruction[4] ),
    .S(net107),
    .X(_01211_));
 sky130_fd_sc_hd__mux2_1 _10203_ (.A0(net28),
    .A1(\core_pipeline.fetch_to_decode_instruction[5] ),
    .S(net107),
    .X(_01212_));
 sky130_fd_sc_hd__mux2_1 _10204_ (.A0(net29),
    .A1(\core_pipeline.fetch_to_decode_instruction[6] ),
    .S(net107),
    .X(_01213_));
 sky130_fd_sc_hd__mux2_1 _10205_ (.A0(net30),
    .A1(\core_pipeline.fetch_to_decode_instruction[7] ),
    .S(net107),
    .X(_01214_));
 sky130_fd_sc_hd__mux2_1 _10206_ (.A0(net31),
    .A1(\core_pipeline.fetch_to_decode_instruction[8] ),
    .S(net107),
    .X(_01215_));
 sky130_fd_sc_hd__mux2_1 _10207_ (.A0(net32),
    .A1(\core_pipeline.fetch_to_decode_instruction[9] ),
    .S(net109),
    .X(_01216_));
 sky130_fd_sc_hd__mux2_1 _10208_ (.A0(net2),
    .A1(\core_pipeline.fetch_to_decode_instruction[10] ),
    .S(net107),
    .X(_01217_));
 sky130_fd_sc_hd__mux2_1 _10209_ (.A0(net3),
    .A1(\core_pipeline.fetch_to_decode_instruction[11] ),
    .S(net108),
    .X(_01218_));
 sky130_fd_sc_hd__mux2_1 _10210_ (.A0(net4),
    .A1(\core_pipeline.fetch_to_decode_instruction[12] ),
    .S(net107),
    .X(_01219_));
 sky130_fd_sc_hd__mux2_1 _10211_ (.A0(net5),
    .A1(\core_pipeline.fetch_to_decode_instruction[13] ),
    .S(net107),
    .X(_01220_));
 sky130_fd_sc_hd__mux2_1 _10212_ (.A0(net6),
    .A1(\core_pipeline.fetch_to_decode_instruction[14] ),
    .S(net107),
    .X(_01221_));
 sky130_fd_sc_hd__mux2_1 _10213_ (.A0(net7),
    .A1(net614),
    .S(net108),
    .X(_01222_));
 sky130_fd_sc_hd__mux2_1 _10214_ (.A0(net8),
    .A1(net602),
    .S(net111),
    .X(_01223_));
 sky130_fd_sc_hd__mux2_1 _10215_ (.A0(net9),
    .A1(net578),
    .S(net110),
    .X(_01224_));
 sky130_fd_sc_hd__mux2_1 _10216_ (.A0(net10),
    .A1(net572),
    .S(net107),
    .X(_01225_));
 sky130_fd_sc_hd__mux2_1 _10217_ (.A0(net11),
    .A1(net569),
    .S(net108),
    .X(_01226_));
 sky130_fd_sc_hd__mux2_1 _10218_ (.A0(net13),
    .A1(net565),
    .S(net109),
    .X(_01227_));
 sky130_fd_sc_hd__mux2_1 _10219_ (.A0(net14),
    .A1(net543),
    .S(net108),
    .X(_01228_));
 sky130_fd_sc_hd__mux2_1 _10220_ (.A0(net15),
    .A1(net521),
    .S(net108),
    .X(_01229_));
 sky130_fd_sc_hd__mux2_1 _10221_ (.A0(net16),
    .A1(net517),
    .S(net109),
    .X(_01230_));
 sky130_fd_sc_hd__mux2_1 _10222_ (.A0(net17),
    .A1(net513),
    .S(net111),
    .X(_01231_));
 sky130_fd_sc_hd__mux2_1 _10223_ (.A0(net18),
    .A1(\core_pipeline.decode_to_csr_read_address[5] ),
    .S(net109),
    .X(_01232_));
 sky130_fd_sc_hd__mux2_1 _10224_ (.A0(net19),
    .A1(\core_pipeline.decode_to_csr_read_address[6] ),
    .S(net109),
    .X(_01233_));
 sky130_fd_sc_hd__mux2_1 _10225_ (.A0(net20),
    .A1(\core_pipeline.decode_to_csr_read_address[7] ),
    .S(net107),
    .X(_01234_));
 sky130_fd_sc_hd__mux2_1 _10226_ (.A0(net21),
    .A1(\core_pipeline.decode_to_csr_read_address[8] ),
    .S(net109),
    .X(_01235_));
 sky130_fd_sc_hd__mux2_1 _10227_ (.A0(net22),
    .A1(\core_pipeline.decode_to_csr_read_address[9] ),
    .S(net107),
    .X(_01236_));
 sky130_fd_sc_hd__mux2_1 _10228_ (.A0(net24),
    .A1(\core_pipeline.decode_to_csr_read_address[10] ),
    .S(net109),
    .X(_01237_));
 sky130_fd_sc_hd__mux2_1 _10229_ (.A0(net25),
    .A1(\core_pipeline.decode_to_csr_read_address[11] ),
    .S(net108),
    .X(_01238_));
 sky130_fd_sc_hd__mux2_1 _10230_ (.A0(\core_pipeline.memory_to_writeback_pc[2] ),
    .A1(\core_pipeline.execute_to_memory_pc[2] ),
    .S(net454),
    .X(_01239_));
 sky130_fd_sc_hd__mux2_1 _10231_ (.A0(\core_pipeline.memory_to_writeback_pc[3] ),
    .A1(\core_pipeline.execute_to_memory_pc[3] ),
    .S(net454),
    .X(_01240_));
 sky130_fd_sc_hd__mux2_1 _10232_ (.A0(\core_pipeline.memory_to_writeback_pc[4] ),
    .A1(\core_pipeline.execute_to_memory_pc[4] ),
    .S(net448),
    .X(_01241_));
 sky130_fd_sc_hd__mux2_1 _10233_ (.A0(\core_pipeline.memory_to_writeback_pc[5] ),
    .A1(\core_pipeline.execute_to_memory_pc[5] ),
    .S(net448),
    .X(_01242_));
 sky130_fd_sc_hd__mux2_1 _10234_ (.A0(\core_pipeline.memory_to_writeback_pc[6] ),
    .A1(\core_pipeline.execute_to_memory_pc[6] ),
    .S(net447),
    .X(_01243_));
 sky130_fd_sc_hd__mux2_1 _10235_ (.A0(\core_pipeline.memory_to_writeback_pc[7] ),
    .A1(\core_pipeline.execute_to_memory_pc[7] ),
    .S(net455),
    .X(_01244_));
 sky130_fd_sc_hd__mux2_1 _10236_ (.A0(\core_pipeline.memory_to_writeback_pc[8] ),
    .A1(\core_pipeline.execute_to_memory_pc[8] ),
    .S(net451),
    .X(_01245_));
 sky130_fd_sc_hd__mux2_1 _10237_ (.A0(\core_pipeline.memory_to_writeback_pc[9] ),
    .A1(\core_pipeline.execute_to_memory_pc[9] ),
    .S(net449),
    .X(_01246_));
 sky130_fd_sc_hd__mux2_1 _10238_ (.A0(\core_pipeline.memory_to_writeback_pc[10] ),
    .A1(\core_pipeline.execute_to_memory_pc[10] ),
    .S(net453),
    .X(_01247_));
 sky130_fd_sc_hd__mux2_1 _10239_ (.A0(\core_pipeline.memory_to_writeback_pc[11] ),
    .A1(\core_pipeline.execute_to_memory_pc[11] ),
    .S(net449),
    .X(_01248_));
 sky130_fd_sc_hd__mux2_1 _10240_ (.A0(\core_pipeline.memory_to_writeback_pc[12] ),
    .A1(\core_pipeline.execute_to_memory_pc[12] ),
    .S(net449),
    .X(_01249_));
 sky130_fd_sc_hd__mux2_1 _10241_ (.A0(\core_pipeline.memory_to_writeback_pc[13] ),
    .A1(\core_pipeline.execute_to_memory_pc[13] ),
    .S(net449),
    .X(_01250_));
 sky130_fd_sc_hd__mux2_1 _10242_ (.A0(\core_pipeline.memory_to_writeback_pc[14] ),
    .A1(\core_pipeline.execute_to_memory_pc[14] ),
    .S(net453),
    .X(_01251_));
 sky130_fd_sc_hd__mux2_1 _10243_ (.A0(\core_pipeline.memory_to_writeback_pc[15] ),
    .A1(\core_pipeline.execute_to_memory_pc[15] ),
    .S(net449),
    .X(_01252_));
 sky130_fd_sc_hd__mux2_1 _10244_ (.A0(\core_pipeline.memory_to_writeback_pc[16] ),
    .A1(\core_pipeline.execute_to_memory_pc[16] ),
    .S(_03432_),
    .X(_01253_));
 sky130_fd_sc_hd__mux2_1 _10245_ (.A0(\core_pipeline.memory_to_writeback_pc[17] ),
    .A1(\core_pipeline.execute_to_memory_pc[17] ),
    .S(net457),
    .X(_01254_));
 sky130_fd_sc_hd__mux2_1 _10246_ (.A0(\core_pipeline.memory_to_writeback_pc[18] ),
    .A1(\core_pipeline.execute_to_memory_pc[18] ),
    .S(net457),
    .X(_01255_));
 sky130_fd_sc_hd__mux2_1 _10247_ (.A0(\core_pipeline.memory_to_writeback_pc[19] ),
    .A1(\core_pipeline.execute_to_memory_pc[19] ),
    .S(net453),
    .X(_01256_));
 sky130_fd_sc_hd__mux2_1 _10248_ (.A0(\core_pipeline.memory_to_writeback_pc[20] ),
    .A1(\core_pipeline.execute_to_memory_pc[20] ),
    .S(net457),
    .X(_01257_));
 sky130_fd_sc_hd__mux2_1 _10249_ (.A0(\core_pipeline.memory_to_writeback_pc[21] ),
    .A1(\core_pipeline.execute_to_memory_pc[21] ),
    .S(net456),
    .X(_01258_));
 sky130_fd_sc_hd__mux2_1 _10250_ (.A0(\core_pipeline.memory_to_writeback_pc[22] ),
    .A1(\core_pipeline.execute_to_memory_pc[22] ),
    .S(net456),
    .X(_01259_));
 sky130_fd_sc_hd__mux2_1 _10251_ (.A0(\core_pipeline.memory_to_writeback_pc[23] ),
    .A1(\core_pipeline.execute_to_memory_pc[23] ),
    .S(net452),
    .X(_01260_));
 sky130_fd_sc_hd__mux2_1 _10252_ (.A0(\core_pipeline.memory_to_writeback_pc[24] ),
    .A1(\core_pipeline.execute_to_memory_pc[24] ),
    .S(net450),
    .X(_01261_));
 sky130_fd_sc_hd__mux2_1 _10253_ (.A0(\core_pipeline.memory_to_writeback_pc[25] ),
    .A1(\core_pipeline.execute_to_memory_pc[25] ),
    .S(net451),
    .X(_01262_));
 sky130_fd_sc_hd__mux2_1 _10254_ (.A0(\core_pipeline.memory_to_writeback_pc[26] ),
    .A1(\core_pipeline.execute_to_memory_pc[26] ),
    .S(net452),
    .X(_01263_));
 sky130_fd_sc_hd__mux2_1 _10255_ (.A0(\core_pipeline.memory_to_writeback_pc[27] ),
    .A1(\core_pipeline.execute_to_memory_pc[27] ),
    .S(net456),
    .X(_01264_));
 sky130_fd_sc_hd__mux2_1 _10256_ (.A0(\core_pipeline.memory_to_writeback_pc[28] ),
    .A1(\core_pipeline.execute_to_memory_pc[28] ),
    .S(net455),
    .X(_01265_));
 sky130_fd_sc_hd__mux2_1 _10257_ (.A0(\core_pipeline.memory_to_writeback_pc[29] ),
    .A1(net656),
    .S(net447),
    .X(_01266_));
 sky130_fd_sc_hd__mux2_1 _10258_ (.A0(\core_pipeline.memory_to_writeback_pc[30] ),
    .A1(\core_pipeline.execute_to_memory_pc[30] ),
    .S(net448),
    .X(_01267_));
 sky130_fd_sc_hd__mux2_1 _10259_ (.A0(\core_pipeline.memory_to_writeback_pc[31] ),
    .A1(\core_pipeline.execute_to_memory_pc[31] ),
    .S(net455),
    .X(_01268_));
 sky130_fd_sc_hd__mux2_1 _10260_ (.A0(\core_pipeline.memory_to_writeback_next_pc[0] ),
    .A1(\core_pipeline.execute_to_memory_next_pc[0] ),
    .S(net446),
    .X(_01269_));
 sky130_fd_sc_hd__mux2_1 _10261_ (.A0(\core_pipeline.memory_to_writeback_next_pc[1] ),
    .A1(\core_pipeline.execute_to_memory_next_pc[1] ),
    .S(net446),
    .X(_01270_));
 sky130_fd_sc_hd__mux2_1 _10262_ (.A0(\core_pipeline.memory_to_writeback_next_pc[2] ),
    .A1(\core_pipeline.execute_to_memory_next_pc[2] ),
    .S(net454),
    .X(_01271_));
 sky130_fd_sc_hd__mux2_1 _10263_ (.A0(\core_pipeline.memory_to_writeback_next_pc[3] ),
    .A1(\core_pipeline.execute_to_memory_next_pc[3] ),
    .S(net454),
    .X(_01272_));
 sky130_fd_sc_hd__mux2_1 _10264_ (.A0(\core_pipeline.memory_to_writeback_next_pc[4] ),
    .A1(\core_pipeline.execute_to_memory_next_pc[4] ),
    .S(net448),
    .X(_01273_));
 sky130_fd_sc_hd__mux2_1 _10265_ (.A0(\core_pipeline.memory_to_writeback_next_pc[5] ),
    .A1(\core_pipeline.execute_to_memory_next_pc[5] ),
    .S(net446),
    .X(_01274_));
 sky130_fd_sc_hd__mux2_1 _10266_ (.A0(\core_pipeline.memory_to_writeback_next_pc[6] ),
    .A1(\core_pipeline.execute_to_memory_next_pc[6] ),
    .S(net447),
    .X(_01275_));
 sky130_fd_sc_hd__mux2_1 _10267_ (.A0(\core_pipeline.memory_to_writeback_next_pc[7] ),
    .A1(\core_pipeline.execute_to_memory_next_pc[7] ),
    .S(net455),
    .X(_01276_));
 sky130_fd_sc_hd__mux2_1 _10268_ (.A0(\core_pipeline.memory_to_writeback_next_pc[8] ),
    .A1(net657),
    .S(net451),
    .X(_01277_));
 sky130_fd_sc_hd__mux2_1 _10269_ (.A0(\core_pipeline.memory_to_writeback_next_pc[9] ),
    .A1(\core_pipeline.execute_to_memory_next_pc[9] ),
    .S(net453),
    .X(_01278_));
 sky130_fd_sc_hd__mux2_1 _10270_ (.A0(\core_pipeline.memory_to_writeback_next_pc[10] ),
    .A1(\core_pipeline.execute_to_memory_next_pc[10] ),
    .S(net453),
    .X(_01279_));
 sky130_fd_sc_hd__mux2_1 _10271_ (.A0(\core_pipeline.memory_to_writeback_next_pc[11] ),
    .A1(\core_pipeline.execute_to_memory_next_pc[11] ),
    .S(net449),
    .X(_01280_));
 sky130_fd_sc_hd__mux2_1 _10272_ (.A0(\core_pipeline.memory_to_writeback_next_pc[12] ),
    .A1(\core_pipeline.execute_to_memory_next_pc[12] ),
    .S(net449),
    .X(_01281_));
 sky130_fd_sc_hd__mux2_1 _10273_ (.A0(\core_pipeline.memory_to_writeback_next_pc[13] ),
    .A1(\core_pipeline.execute_to_memory_next_pc[13] ),
    .S(net449),
    .X(_01282_));
 sky130_fd_sc_hd__mux2_1 _10274_ (.A0(\core_pipeline.memory_to_writeback_next_pc[14] ),
    .A1(\core_pipeline.execute_to_memory_next_pc[14] ),
    .S(net453),
    .X(_01283_));
 sky130_fd_sc_hd__mux2_1 _10275_ (.A0(\core_pipeline.memory_to_writeback_next_pc[15] ),
    .A1(\core_pipeline.execute_to_memory_next_pc[15] ),
    .S(net450),
    .X(_01284_));
 sky130_fd_sc_hd__mux2_1 _10276_ (.A0(\core_pipeline.memory_to_writeback_next_pc[16] ),
    .A1(\core_pipeline.execute_to_memory_next_pc[16] ),
    .S(net449),
    .X(_01285_));
 sky130_fd_sc_hd__mux2_1 _10277_ (.A0(\core_pipeline.memory_to_writeback_next_pc[17] ),
    .A1(\core_pipeline.execute_to_memory_next_pc[17] ),
    .S(net457),
    .X(_01286_));
 sky130_fd_sc_hd__mux2_1 _10278_ (.A0(\core_pipeline.memory_to_writeback_next_pc[18] ),
    .A1(\core_pipeline.execute_to_memory_next_pc[18] ),
    .S(net457),
    .X(_01287_));
 sky130_fd_sc_hd__mux2_1 _10279_ (.A0(\core_pipeline.memory_to_writeback_next_pc[19] ),
    .A1(\core_pipeline.execute_to_memory_next_pc[19] ),
    .S(net457),
    .X(_01288_));
 sky130_fd_sc_hd__mux2_1 _10280_ (.A0(\core_pipeline.memory_to_writeback_next_pc[20] ),
    .A1(\core_pipeline.execute_to_memory_next_pc[20] ),
    .S(net457),
    .X(_01289_));
 sky130_fd_sc_hd__mux2_1 _10281_ (.A0(\core_pipeline.memory_to_writeback_next_pc[21] ),
    .A1(\core_pipeline.execute_to_memory_next_pc[21] ),
    .S(net456),
    .X(_01290_));
 sky130_fd_sc_hd__mux2_1 _10282_ (.A0(\core_pipeline.memory_to_writeback_next_pc[22] ),
    .A1(\core_pipeline.execute_to_memory_next_pc[22] ),
    .S(net456),
    .X(_01291_));
 sky130_fd_sc_hd__mux2_1 _10283_ (.A0(\core_pipeline.memory_to_writeback_next_pc[23] ),
    .A1(\core_pipeline.execute_to_memory_next_pc[23] ),
    .S(net453),
    .X(_01292_));
 sky130_fd_sc_hd__mux2_1 _10284_ (.A0(\core_pipeline.memory_to_writeback_next_pc[24] ),
    .A1(\core_pipeline.execute_to_memory_next_pc[24] ),
    .S(net451),
    .X(_01293_));
 sky130_fd_sc_hd__mux2_1 _10285_ (.A0(\core_pipeline.memory_to_writeback_next_pc[25] ),
    .A1(\core_pipeline.execute_to_memory_next_pc[25] ),
    .S(net451),
    .X(_01294_));
 sky130_fd_sc_hd__mux2_1 _10286_ (.A0(\core_pipeline.memory_to_writeback_next_pc[26] ),
    .A1(\core_pipeline.execute_to_memory_next_pc[26] ),
    .S(net453),
    .X(_01295_));
 sky130_fd_sc_hd__mux2_1 _10287_ (.A0(\core_pipeline.memory_to_writeback_next_pc[27] ),
    .A1(\core_pipeline.execute_to_memory_next_pc[27] ),
    .S(net456),
    .X(_01296_));
 sky130_fd_sc_hd__mux2_1 _10288_ (.A0(\core_pipeline.memory_to_writeback_next_pc[28] ),
    .A1(\core_pipeline.execute_to_memory_next_pc[28] ),
    .S(net454),
    .X(_01297_));
 sky130_fd_sc_hd__mux2_1 _10289_ (.A0(\core_pipeline.memory_to_writeback_next_pc[29] ),
    .A1(\core_pipeline.execute_to_memory_next_pc[29] ),
    .S(net452),
    .X(_01298_));
 sky130_fd_sc_hd__mux2_1 _10290_ (.A0(\core_pipeline.memory_to_writeback_next_pc[30] ),
    .A1(\core_pipeline.execute_to_memory_next_pc[30] ),
    .S(net447),
    .X(_01299_));
 sky130_fd_sc_hd__mux2_1 _10291_ (.A0(\core_pipeline.memory_to_writeback_next_pc[31] ),
    .A1(\core_pipeline.execute_to_memory_next_pc[31] ),
    .S(net454),
    .X(_01300_));
 sky130_fd_sc_hd__mux2_1 _10292_ (.A0(\core_pipeline.memory_to_writeback_csr_data[0] ),
    .A1(\core_pipeline.execute_to_memory_csr_data[0] ),
    .S(net448),
    .X(_01301_));
 sky130_fd_sc_hd__mux2_1 _10293_ (.A0(\core_pipeline.memory_to_writeback_csr_data[1] ),
    .A1(\core_pipeline.execute_to_memory_csr_data[1] ),
    .S(net446),
    .X(_01302_));
 sky130_fd_sc_hd__mux2_1 _10294_ (.A0(\core_pipeline.memory_to_writeback_csr_data[2] ),
    .A1(\core_pipeline.execute_to_memory_csr_data[2] ),
    .S(net454),
    .X(_01303_));
 sky130_fd_sc_hd__mux2_1 _10295_ (.A0(\core_pipeline.memory_to_writeback_csr_data[3] ),
    .A1(\core_pipeline.execute_to_memory_csr_data[3] ),
    .S(net448),
    .X(_01304_));
 sky130_fd_sc_hd__mux2_1 _10296_ (.A0(\core_pipeline.memory_to_writeback_csr_data[4] ),
    .A1(\core_pipeline.execute_to_memory_csr_data[4] ),
    .S(net448),
    .X(_01305_));
 sky130_fd_sc_hd__mux2_1 _10297_ (.A0(\core_pipeline.memory_to_writeback_csr_data[5] ),
    .A1(\core_pipeline.execute_to_memory_csr_data[5] ),
    .S(net446),
    .X(_01306_));
 sky130_fd_sc_hd__mux2_1 _10298_ (.A0(\core_pipeline.memory_to_writeback_csr_data[6] ),
    .A1(\core_pipeline.execute_to_memory_csr_data[6] ),
    .S(net447),
    .X(_01307_));
 sky130_fd_sc_hd__mux2_1 _10299_ (.A0(\core_pipeline.memory_to_writeback_csr_data[7] ),
    .A1(\core_pipeline.execute_to_memory_csr_data[7] ),
    .S(net448),
    .X(_01308_));
 sky130_fd_sc_hd__mux2_1 _10300_ (.A0(\core_pipeline.memory_to_writeback_csr_data[8] ),
    .A1(\core_pipeline.execute_to_memory_csr_data[8] ),
    .S(net450),
    .X(_01309_));
 sky130_fd_sc_hd__mux2_1 _10301_ (.A0(\core_pipeline.memory_to_writeback_csr_data[9] ),
    .A1(\core_pipeline.execute_to_memory_csr_data[9] ),
    .S(net450),
    .X(_01310_));
 sky130_fd_sc_hd__mux2_1 _10302_ (.A0(\core_pipeline.memory_to_writeback_csr_data[10] ),
    .A1(\core_pipeline.execute_to_memory_csr_data[10] ),
    .S(net450),
    .X(_01311_));
 sky130_fd_sc_hd__mux2_1 _10303_ (.A0(\core_pipeline.memory_to_writeback_csr_data[11] ),
    .A1(\core_pipeline.execute_to_memory_csr_data[11] ),
    .S(net448),
    .X(_01312_));
 sky130_fd_sc_hd__mux2_1 _10304_ (.A0(\core_pipeline.memory_to_writeback_csr_data[12] ),
    .A1(\core_pipeline.execute_to_memory_csr_data[12] ),
    .S(net449),
    .X(_01313_));
 sky130_fd_sc_hd__mux2_1 _10305_ (.A0(\core_pipeline.memory_to_writeback_csr_data[13] ),
    .A1(\core_pipeline.execute_to_memory_csr_data[13] ),
    .S(net449),
    .X(_01314_));
 sky130_fd_sc_hd__mux2_1 _10306_ (.A0(\core_pipeline.memory_to_writeback_csr_data[14] ),
    .A1(\core_pipeline.execute_to_memory_csr_data[14] ),
    .S(net449),
    .X(_01315_));
 sky130_fd_sc_hd__mux2_1 _10307_ (.A0(\core_pipeline.memory_to_writeback_csr_data[15] ),
    .A1(\core_pipeline.execute_to_memory_csr_data[15] ),
    .S(net450),
    .X(_01316_));
 sky130_fd_sc_hd__mux2_1 _10308_ (.A0(\core_pipeline.memory_to_writeback_csr_data[16] ),
    .A1(\core_pipeline.execute_to_memory_csr_data[16] ),
    .S(net449),
    .X(_01317_));
 sky130_fd_sc_hd__mux2_1 _10309_ (.A0(\core_pipeline.memory_to_writeback_csr_data[17] ),
    .A1(\core_pipeline.execute_to_memory_csr_data[17] ),
    .S(net457),
    .X(_01318_));
 sky130_fd_sc_hd__mux2_1 _10310_ (.A0(\core_pipeline.memory_to_writeback_csr_data[18] ),
    .A1(\core_pipeline.execute_to_memory_csr_data[18] ),
    .S(net456),
    .X(_01319_));
 sky130_fd_sc_hd__mux2_1 _10311_ (.A0(\core_pipeline.memory_to_writeback_csr_data[19] ),
    .A1(\core_pipeline.execute_to_memory_csr_data[19] ),
    .S(net456),
    .X(_01320_));
 sky130_fd_sc_hd__mux2_1 _10312_ (.A0(\core_pipeline.memory_to_writeback_csr_data[20] ),
    .A1(\core_pipeline.execute_to_memory_csr_data[20] ),
    .S(net456),
    .X(_01321_));
 sky130_fd_sc_hd__mux2_1 _10313_ (.A0(\core_pipeline.memory_to_writeback_csr_data[21] ),
    .A1(\core_pipeline.execute_to_memory_csr_data[21] ),
    .S(net456),
    .X(_01322_));
 sky130_fd_sc_hd__mux2_1 _10314_ (.A0(\core_pipeline.memory_to_writeback_csr_data[22] ),
    .A1(\core_pipeline.execute_to_memory_csr_data[22] ),
    .S(net452),
    .X(_01323_));
 sky130_fd_sc_hd__mux2_1 _10315_ (.A0(\core_pipeline.memory_to_writeback_csr_data[23] ),
    .A1(\core_pipeline.execute_to_memory_csr_data[23] ),
    .S(net452),
    .X(_01324_));
 sky130_fd_sc_hd__mux2_1 _10316_ (.A0(\core_pipeline.memory_to_writeback_csr_data[24] ),
    .A1(\core_pipeline.execute_to_memory_csr_data[24] ),
    .S(net452),
    .X(_01325_));
 sky130_fd_sc_hd__mux2_1 _10317_ (.A0(\core_pipeline.memory_to_writeback_csr_data[25] ),
    .A1(\core_pipeline.execute_to_memory_csr_data[25] ),
    .S(net450),
    .X(_01326_));
 sky130_fd_sc_hd__mux2_1 _10318_ (.A0(\core_pipeline.memory_to_writeback_csr_data[26] ),
    .A1(\core_pipeline.execute_to_memory_csr_data[26] ),
    .S(net450),
    .X(_01327_));
 sky130_fd_sc_hd__mux2_1 _10319_ (.A0(\core_pipeline.memory_to_writeback_csr_data[27] ),
    .A1(\core_pipeline.execute_to_memory_csr_data[27] ),
    .S(net456),
    .X(_01328_));
 sky130_fd_sc_hd__mux2_1 _10320_ (.A0(\core_pipeline.memory_to_writeback_csr_data[28] ),
    .A1(\core_pipeline.execute_to_memory_csr_data[28] ),
    .S(net454),
    .X(_01329_));
 sky130_fd_sc_hd__mux2_1 _10321_ (.A0(\core_pipeline.memory_to_writeback_csr_data[29] ),
    .A1(\core_pipeline.execute_to_memory_csr_data[29] ),
    .S(net446),
    .X(_01330_));
 sky130_fd_sc_hd__mux2_1 _10322_ (.A0(\core_pipeline.memory_to_writeback_csr_data[30] ),
    .A1(\core_pipeline.execute_to_memory_csr_data[30] ),
    .S(net446),
    .X(_01331_));
 sky130_fd_sc_hd__mux2_1 _10323_ (.A0(\core_pipeline.memory_to_writeback_csr_data[31] ),
    .A1(\core_pipeline.execute_to_memory_csr_data[31] ),
    .S(net454),
    .X(_01332_));
 sky130_fd_sc_hd__mux2_1 _10324_ (.A0(\core_pipeline.execute_to_memory_csr_write ),
    .A1(\core_pipeline.memory_to_writeback_csr_write ),
    .S(net458),
    .X(_01333_));
 sky130_fd_sc_hd__mux2_1 _10325_ (.A0(net510),
    .A1(net499),
    .S(net454),
    .X(_01334_));
 sky130_fd_sc_hd__mux2_1 _10326_ (.A0(net508),
    .A1(\core_pipeline.execute_to_memory_write_select[1] ),
    .S(net446),
    .X(_01335_));
 sky130_fd_sc_hd__mux2_1 _10327_ (.A0(\core_pipeline.execute_to_memory_rd_address[0] ),
    .A1(\core_pipeline.memory_to_writeback_rd_address[0] ),
    .S(_03431_),
    .X(_01336_));
 sky130_fd_sc_hd__mux2_1 _10328_ (.A0(\core_pipeline.execute_to_memory_rd_address[1] ),
    .A1(\core_pipeline.memory_to_writeback_rd_address[1] ),
    .S(_03431_),
    .X(_01337_));
 sky130_fd_sc_hd__mux2_1 _10329_ (.A0(\core_pipeline.execute_to_memory_rd_address[2] ),
    .A1(\core_pipeline.memory_to_writeback_rd_address[2] ),
    .S(_03431_),
    .X(_01338_));
 sky130_fd_sc_hd__mux2_1 _10330_ (.A0(\core_pipeline.execute_to_memory_rd_address[3] ),
    .A1(\core_pipeline.memory_to_writeback_rd_address[3] ),
    .S(_03431_),
    .X(_01339_));
 sky130_fd_sc_hd__mux2_1 _10331_ (.A0(\core_pipeline.execute_to_memory_rd_address[4] ),
    .A1(\core_pipeline.memory_to_writeback_rd_address[4] ),
    .S(net458),
    .X(_01340_));
 sky130_fd_sc_hd__mux2_1 _10332_ (.A0(\core_pipeline.memory_to_writeback_csr_address[0] ),
    .A1(\core_pipeline.execute_to_memory_csr_address[0] ),
    .S(net455),
    .X(_01341_));
 sky130_fd_sc_hd__mux2_1 _10333_ (.A0(\core_pipeline.memory_to_writeback_csr_address[1] ),
    .A1(\core_pipeline.execute_to_memory_csr_address[1] ),
    .S(net455),
    .X(_01342_));
 sky130_fd_sc_hd__mux2_1 _10334_ (.A0(\core_pipeline.memory_to_writeback_csr_address[2] ),
    .A1(\core_pipeline.execute_to_memory_csr_address[2] ),
    .S(net455),
    .X(_01343_));
 sky130_fd_sc_hd__mux2_1 _10335_ (.A0(\core_pipeline.memory_to_writeback_csr_address[3] ),
    .A1(\core_pipeline.execute_to_memory_csr_address[3] ),
    .S(net455),
    .X(_01344_));
 sky130_fd_sc_hd__mux2_1 _10336_ (.A0(\core_pipeline.memory_to_writeback_csr_address[4] ),
    .A1(\core_pipeline.execute_to_memory_csr_address[4] ),
    .S(net455),
    .X(_01345_));
 sky130_fd_sc_hd__mux2_1 _10337_ (.A0(\core_pipeline.memory_to_writeback_csr_address[5] ),
    .A1(\core_pipeline.execute_to_memory_csr_address[5] ),
    .S(net455),
    .X(_01346_));
 sky130_fd_sc_hd__mux2_1 _10338_ (.A0(\core_pipeline.memory_to_writeback_csr_address[6] ),
    .A1(\core_pipeline.execute_to_memory_csr_address[6] ),
    .S(net455),
    .X(_01347_));
 sky130_fd_sc_hd__mux2_1 _10339_ (.A0(\core_pipeline.memory_to_writeback_csr_address[7] ),
    .A1(\core_pipeline.execute_to_memory_csr_address[7] ),
    .S(net455),
    .X(_01348_));
 sky130_fd_sc_hd__mux2_1 _10340_ (.A0(\core_pipeline.memory_to_writeback_csr_address[8] ),
    .A1(\core_pipeline.execute_to_memory_csr_address[8] ),
    .S(net455),
    .X(_01349_));
 sky130_fd_sc_hd__mux2_1 _10341_ (.A0(\core_pipeline.memory_to_writeback_csr_address[9] ),
    .A1(\core_pipeline.execute_to_memory_csr_address[9] ),
    .S(net455),
    .X(_01350_));
 sky130_fd_sc_hd__mux2_1 _10342_ (.A0(\core_pipeline.memory_to_writeback_csr_address[10] ),
    .A1(\core_pipeline.execute_to_memory_csr_address[10] ),
    .S(net455),
    .X(_01351_));
 sky130_fd_sc_hd__mux2_1 _10343_ (.A0(\core_pipeline.memory_to_writeback_csr_address[11] ),
    .A1(\core_pipeline.execute_to_memory_csr_address[11] ),
    .S(net455),
    .X(_01352_));
 sky130_fd_sc_hd__mux2_1 _10344_ (.A0(\core_pipeline.execute_to_memory_mret ),
    .A1(\core_pipeline.memory_to_writeback_mret ),
    .S(net458),
    .X(_01353_));
 sky130_fd_sc_hd__and3b_1 _10345_ (.A_N(\core_pipeline.decode_to_execute_alu_function[2] ),
    .B(\core_pipeline.decode_to_execute_alu_function[1] ),
    .C(\core_pipeline.decode_to_execute_alu_function[0] ),
    .X(_05610_));
 sky130_fd_sc_hd__a22o_1 _10346_ (.A1(net501),
    .A2(\core_pipeline.decode_to_execute_csr_data[31] ),
    .B1(\core_pipeline.decode_to_execute_imm_data[31] ),
    .B2(net503),
    .X(_05611_));
 sky130_fd_sc_hd__a21oi_4 _10347_ (.A1(_03741_),
    .A2(net434),
    .B1(_05611_),
    .Y(_05612_));
 sky130_fd_sc_hd__a22o_1 _10348_ (.A1(net628),
    .A2(\core_pipeline.decode_to_execute_imm_data[31] ),
    .B1(\core_pipeline.decode_to_execute_pc[31] ),
    .B2(net630),
    .X(_05613_));
 sky130_fd_sc_hd__a21o_4 _10349_ (.A1(_03743_),
    .A2(net432),
    .B1(_05613_),
    .X(_05614_));
 sky130_fd_sc_hd__inv_2 _10350_ (.A(_05614_),
    .Y(_05615_));
 sky130_fd_sc_hd__or2_2 _10351_ (.A(_05612_),
    .B(_05614_),
    .X(_05616_));
 sky130_fd_sc_hd__a22o_2 _10352_ (.A1(net500),
    .A2(\core_pipeline.decode_to_execute_csr_data[14] ),
    .B1(\core_pipeline.decode_to_execute_imm_data[14] ),
    .B2(net502),
    .X(_05617_));
 sky130_fd_sc_hd__a21oi_4 _10353_ (.A1(_03826_),
    .A2(net433),
    .B1(_05617_),
    .Y(_05618_));
 sky130_fd_sc_hd__nand2_1 _10354_ (.A(_04608_),
    .B(_05618_),
    .Y(_05619_));
 sky130_fd_sc_hd__or2_1 _10355_ (.A(_04608_),
    .B(_05618_),
    .X(_05620_));
 sky130_fd_sc_hd__and2_1 _10356_ (.A(_05619_),
    .B(_05620_),
    .X(_05621_));
 sky130_fd_sc_hd__a22o_1 _10357_ (.A1(net501),
    .A2(\core_pipeline.decode_to_execute_csr_data[13] ),
    .B1(\core_pipeline.decode_to_execute_imm_data[13] ),
    .B2(net503),
    .X(_05622_));
 sky130_fd_sc_hd__a21o_4 _10358_ (.A1(_03830_),
    .A2(net433),
    .B1(_05622_),
    .X(_05623_));
 sky130_fd_sc_hd__nor2_1 _10359_ (.A(_04599_),
    .B(_05623_),
    .Y(_05624_));
 sky130_fd_sc_hd__and2_2 _10360_ (.A(_03822_),
    .B(net433),
    .X(_05625_));
 sky130_fd_sc_hd__a221oi_4 _10361_ (.A1(net501),
    .A2(\core_pipeline.decode_to_execute_csr_data[15] ),
    .B1(\core_pipeline.decode_to_execute_imm_data[15] ),
    .B2(net503),
    .C1(_05625_),
    .Y(_05626_));
 sky130_fd_sc_hd__a221o_4 _10362_ (.A1(\core_pipeline.pipeline_decode.alu_select_b_out[2] ),
    .A2(\core_pipeline.decode_to_execute_csr_data[15] ),
    .B1(\core_pipeline.decode_to_execute_imm_data[15] ),
    .B2(\core_pipeline.pipeline_decode.alu_select_b_out[1] ),
    .C1(_05625_),
    .X(_05627_));
 sky130_fd_sc_hd__nand2_1 _10363_ (.A(_04618_),
    .B(_05626_),
    .Y(_05628_));
 sky130_fd_sc_hd__or2_1 _10364_ (.A(_04618_),
    .B(_05626_),
    .X(_05629_));
 sky130_fd_sc_hd__nand2_1 _10365_ (.A(_05628_),
    .B(_05629_),
    .Y(_05630_));
 sky130_fd_sc_hd__or3_2 _10366_ (.A(_05621_),
    .B(_05624_),
    .C(_05630_),
    .X(_05631_));
 sky130_fd_sc_hd__a22o_1 _10367_ (.A1(net500),
    .A2(\core_pipeline.decode_to_execute_csr_data[8] ),
    .B1(\core_pipeline.decode_to_execute_imm_data[8] ),
    .B2(net502),
    .X(_05632_));
 sky130_fd_sc_hd__a21oi_4 _10368_ (.A1(_03852_),
    .A2(net433),
    .B1(_05632_),
    .Y(_05633_));
 sky130_fd_sc_hd__xor2_1 _10369_ (.A(_04553_),
    .B(_05633_),
    .X(_05634_));
 sky130_fd_sc_hd__a22o_2 _10370_ (.A1(net500),
    .A2(\core_pipeline.decode_to_execute_csr_data[9] ),
    .B1(\core_pipeline.decode_to_execute_imm_data[9] ),
    .B2(net502),
    .X(_05635_));
 sky130_fd_sc_hd__a21oi_4 _10371_ (.A1(_03847_),
    .A2(net433),
    .B1(_05635_),
    .Y(_05636_));
 sky130_fd_sc_hd__xor2_2 _10372_ (.A(_04565_),
    .B(_05636_),
    .X(_05637_));
 sky130_fd_sc_hd__a22o_2 _10373_ (.A1(\core_pipeline.pipeline_decode.alu_select_b_out[2] ),
    .A2(\core_pipeline.decode_to_execute_csr_data[11] ),
    .B1(\core_pipeline.decode_to_execute_imm_data[11] ),
    .B2(\core_pipeline.pipeline_decode.alu_select_b_out[1] ),
    .X(_05638_));
 sky130_fd_sc_hd__a21oi_4 _10374_ (.A1(_03843_),
    .A2(net433),
    .B1(_05638_),
    .Y(_05639_));
 sky130_fd_sc_hd__xor2_1 _10375_ (.A(_04581_),
    .B(_05639_),
    .X(_05640_));
 sky130_fd_sc_hd__a22o_1 _10376_ (.A1(\core_pipeline.pipeline_decode.alu_select_b_out[2] ),
    .A2(\core_pipeline.decode_to_execute_csr_data[12] ),
    .B1(\core_pipeline.decode_to_execute_imm_data[12] ),
    .B2(\core_pipeline.pipeline_decode.alu_select_b_out[1] ),
    .X(_05641_));
 sky130_fd_sc_hd__a21o_4 _10377_ (.A1(_03836_),
    .A2(net433),
    .B1(_05641_),
    .X(_05642_));
 sky130_fd_sc_hd__nand2_1 _10378_ (.A(net371),
    .B(_05642_),
    .Y(_05643_));
 sky130_fd_sc_hd__nor2_1 _10379_ (.A(net371),
    .B(_05642_),
    .Y(_05644_));
 sky130_fd_sc_hd__or2_1 _10380_ (.A(net371),
    .B(_05642_),
    .X(_05645_));
 sky130_fd_sc_hd__nand2_1 _10381_ (.A(_05643_),
    .B(_05645_),
    .Y(_05646_));
 sky130_fd_sc_hd__or4_1 _10382_ (.A(_05634_),
    .B(_05637_),
    .C(_05640_),
    .D(_05646_),
    .X(_05647_));
 sky130_fd_sc_hd__nand2_1 _10383_ (.A(_04599_),
    .B(_05623_),
    .Y(_05648_));
 sky130_fd_sc_hd__inv_2 _10384_ (.A(_05648_),
    .Y(_05649_));
 sky130_fd_sc_hd__a22o_2 _10385_ (.A1(net500),
    .A2(\core_pipeline.decode_to_execute_csr_data[10] ),
    .B1(\core_pipeline.decode_to_execute_imm_data[10] ),
    .B2(net502),
    .X(_05650_));
 sky130_fd_sc_hd__a21oi_4 _10386_ (.A1(_03840_),
    .A2(net433),
    .B1(_05650_),
    .Y(_05651_));
 sky130_fd_sc_hd__and2_1 _10387_ (.A(_04574_),
    .B(_05651_),
    .X(_05652_));
 sky130_fd_sc_hd__or2_1 _10388_ (.A(_04574_),
    .B(_05651_),
    .X(_05653_));
 sky130_fd_sc_hd__nand2b_1 _10389_ (.A_N(_05652_),
    .B(_05653_),
    .Y(_05654_));
 sky130_fd_sc_hd__or3_4 _10390_ (.A(_05647_),
    .B(_05649_),
    .C(_05654_),
    .X(_05655_));
 sky130_fd_sc_hd__a22o_1 _10391_ (.A1(net501),
    .A2(\core_pipeline.decode_to_execute_csr_data[7] ),
    .B1(\core_pipeline.decode_to_execute_imm_data[7] ),
    .B2(net503),
    .X(_05656_));
 sky130_fd_sc_hd__a21oi_4 _10392_ (.A1(_03862_),
    .A2(net434),
    .B1(_05656_),
    .Y(_05657_));
 sky130_fd_sc_hd__nand2b_1 _10393_ (.A_N(_04545_),
    .B(_05657_),
    .Y(_05658_));
 sky130_fd_sc_hd__nand2b_1 _10394_ (.A_N(_05657_),
    .B(_04545_),
    .Y(_05659_));
 sky130_fd_sc_hd__nand2_1 _10395_ (.A(_05658_),
    .B(_05659_),
    .Y(_05660_));
 sky130_fd_sc_hd__a22o_1 _10396_ (.A1(net501),
    .A2(\core_pipeline.decode_to_execute_csr_data[6] ),
    .B1(\core_pipeline.decode_to_execute_imm_data[6] ),
    .B2(net503),
    .X(_05661_));
 sky130_fd_sc_hd__a21oi_4 _10397_ (.A1(_03859_),
    .A2(net434),
    .B1(_05661_),
    .Y(_05662_));
 sky130_fd_sc_hd__xnor2_1 _10398_ (.A(_04538_),
    .B(_05662_),
    .Y(_05663_));
 sky130_fd_sc_hd__or2_1 _10399_ (.A(_05660_),
    .B(_05663_),
    .X(_05664_));
 sky130_fd_sc_hd__a22o_1 _10400_ (.A1(net501),
    .A2(\core_pipeline.decode_to_execute_csr_data[5] ),
    .B1(\core_pipeline.decode_to_execute_imm_data[5] ),
    .B2(net503),
    .X(_05665_));
 sky130_fd_sc_hd__a21oi_4 _10401_ (.A1(_03866_),
    .A2(net434),
    .B1(_05665_),
    .Y(_05666_));
 sky130_fd_sc_hd__or2_1 _10402_ (.A(_04530_),
    .B(_05666_),
    .X(_05667_));
 sky130_fd_sc_hd__nor2_1 _10403_ (.A(_04497_),
    .B(_04502_),
    .Y(_05668_));
 sky130_fd_sc_hd__a211o_1 _10404_ (.A1(net384),
    .A2(_04511_),
    .B1(_05668_),
    .C1(_04508_),
    .X(_05669_));
 sky130_fd_sc_hd__o221a_1 _10405_ (.A1(net384),
    .A2(_04511_),
    .B1(_04517_),
    .B2(net395),
    .C1(_05669_),
    .X(_05670_));
 sky130_fd_sc_hd__a221o_1 _10406_ (.A1(net395),
    .A2(_04517_),
    .B1(_04523_),
    .B2(net391),
    .C1(_05670_),
    .X(_05671_));
 sky130_fd_sc_hd__nand2_1 _10407_ (.A(_04530_),
    .B(_05666_),
    .Y(_05672_));
 sky130_fd_sc_hd__o211ai_1 _10408_ (.A1(net391),
    .A2(_04523_),
    .B1(_05671_),
    .C1(_05672_),
    .Y(_05673_));
 sky130_fd_sc_hd__xnor2_1 _10409_ (.A(net393),
    .B(_04522_),
    .Y(_05674_));
 sky130_fd_sc_hd__nand2_1 _10410_ (.A(_05667_),
    .B(_05672_),
    .Y(_05675_));
 sky130_fd_sc_hd__a21o_1 _10411_ (.A1(_05667_),
    .A2(_05673_),
    .B1(_05664_),
    .X(_05676_));
 sky130_fd_sc_hd__or3b_1 _10412_ (.A(_05662_),
    .B(_04538_),
    .C_N(_05658_),
    .X(_05677_));
 sky130_fd_sc_hd__a31o_2 _10413_ (.A1(_05659_),
    .A2(_05676_),
    .A3(_05677_),
    .B1(_05655_),
    .X(_05678_));
 sky130_fd_sc_hd__o32a_1 _10414_ (.A1(_04554_),
    .A2(_05633_),
    .A3(_05637_),
    .B1(_05636_),
    .B2(_04566_),
    .X(_05679_));
 sky130_fd_sc_hd__o221a_1 _10415_ (.A1(_04582_),
    .A2(_05639_),
    .B1(_05652_),
    .B2(_05679_),
    .C1(_05653_),
    .X(_05680_));
 sky130_fd_sc_hd__a211o_1 _10416_ (.A1(_04582_),
    .A2(_05639_),
    .B1(_05644_),
    .C1(_05680_),
    .X(_05681_));
 sky130_fd_sc_hd__a41o_1 _10417_ (.A1(_05643_),
    .A2(_05648_),
    .A3(_05678_),
    .A4(_05681_),
    .B1(_05631_),
    .X(_05682_));
 sky130_fd_sc_hd__nand3b_1 _10418_ (.A_N(_05618_),
    .B(_05628_),
    .C(_04608_),
    .Y(_05683_));
 sky130_fd_sc_hd__nand2_1 _10419_ (.A(_05612_),
    .B(_05614_),
    .Y(_05684_));
 sky130_fd_sc_hd__nand2_2 _10420_ (.A(_05616_),
    .B(_05684_),
    .Y(_05685_));
 sky130_fd_sc_hd__a22o_1 _10421_ (.A1(net628),
    .A2(\core_pipeline.decode_to_execute_imm_data[30] ),
    .B1(\core_pipeline.decode_to_execute_pc[30] ),
    .B2(net630),
    .X(_05686_));
 sky130_fd_sc_hd__a21o_4 _10422_ (.A1(_03770_),
    .A2(net432),
    .B1(_05686_),
    .X(_05687_));
 sky130_fd_sc_hd__clkinv_4 _10423_ (.A(_05687_),
    .Y(_05688_));
 sky130_fd_sc_hd__a22o_1 _10424_ (.A1(net501),
    .A2(\core_pipeline.decode_to_execute_csr_data[30] ),
    .B1(\core_pipeline.decode_to_execute_imm_data[30] ),
    .B2(net503),
    .X(_05689_));
 sky130_fd_sc_hd__a21o_4 _10425_ (.A1(_03771_),
    .A2(net434),
    .B1(_05689_),
    .X(_05690_));
 sky130_fd_sc_hd__inv_2 _10426_ (.A(_05690_),
    .Y(_05691_));
 sky130_fd_sc_hd__or2_1 _10427_ (.A(_05687_),
    .B(_05690_),
    .X(_05692_));
 sky130_fd_sc_hd__nand2_1 _10428_ (.A(_05687_),
    .B(_05690_),
    .Y(_05693_));
 sky130_fd_sc_hd__and2_1 _10429_ (.A(_05692_),
    .B(_05693_),
    .X(_05694_));
 sky130_fd_sc_hd__or2_1 _10430_ (.A(_05685_),
    .B(_05694_),
    .X(_05695_));
 sky130_fd_sc_hd__a22o_1 _10431_ (.A1(net500),
    .A2(\core_pipeline.decode_to_execute_csr_data[28] ),
    .B1(\core_pipeline.decode_to_execute_imm_data[28] ),
    .B2(net502),
    .X(_05696_));
 sky130_fd_sc_hd__a21oi_4 _10432_ (.A1(_03749_),
    .A2(_04474_),
    .B1(_05696_),
    .Y(_05697_));
 sky130_fd_sc_hd__a22o_1 _10433_ (.A1(net627),
    .A2(\core_pipeline.decode_to_execute_imm_data[28] ),
    .B1(\core_pipeline.decode_to_execute_pc[28] ),
    .B2(net629),
    .X(_05698_));
 sky130_fd_sc_hd__a21o_4 _10434_ (.A1(_03750_),
    .A2(net431),
    .B1(_05698_),
    .X(_05699_));
 sky130_fd_sc_hd__xnor2_2 _10435_ (.A(_05697_),
    .B(_05699_),
    .Y(_05700_));
 sky130_fd_sc_hd__a22o_1 _10436_ (.A1(net500),
    .A2(\core_pipeline.decode_to_execute_csr_data[29] ),
    .B1(\core_pipeline.decode_to_execute_imm_data[29] ),
    .B2(net502),
    .X(_05701_));
 sky130_fd_sc_hd__a21o_4 _10437_ (.A1(_03746_),
    .A2(net433),
    .B1(_05701_),
    .X(_05702_));
 sky130_fd_sc_hd__a22o_1 _10438_ (.A1(net627),
    .A2(\core_pipeline.decode_to_execute_imm_data[29] ),
    .B1(\core_pipeline.decode_to_execute_pc[29] ),
    .B2(\core_pipeline.pipeline_decode.alu_select_a_out[1] ),
    .X(_05703_));
 sky130_fd_sc_hd__a21oi_4 _10439_ (.A1(_03747_),
    .A2(net432),
    .B1(_05703_),
    .Y(_05704_));
 sky130_fd_sc_hd__nor2_1 _10440_ (.A(_05702_),
    .B(_05704_),
    .Y(_05705_));
 sky130_fd_sc_hd__and2_1 _10441_ (.A(_05702_),
    .B(_05704_),
    .X(_05706_));
 sky130_fd_sc_hd__inv_2 _10442_ (.A(_05706_),
    .Y(_05707_));
 sky130_fd_sc_hd__or2_1 _10443_ (.A(_05705_),
    .B(_05706_),
    .X(_05708_));
 sky130_fd_sc_hd__a22o_1 _10444_ (.A1(net501),
    .A2(\core_pipeline.decode_to_execute_csr_data[26] ),
    .B1(\core_pipeline.decode_to_execute_imm_data[26] ),
    .B2(net503),
    .X(_05709_));
 sky130_fd_sc_hd__a21oi_4 _10445_ (.A1(_03756_),
    .A2(net433),
    .B1(_05709_),
    .Y(_05710_));
 sky130_fd_sc_hd__a22o_1 _10446_ (.A1(net627),
    .A2(\core_pipeline.decode_to_execute_imm_data[26] ),
    .B1(\core_pipeline.decode_to_execute_pc[26] ),
    .B2(net629),
    .X(_05711_));
 sky130_fd_sc_hd__a21o_4 _10447_ (.A1(_03758_),
    .A2(net431),
    .B1(_05711_),
    .X(_05712_));
 sky130_fd_sc_hd__xnor2_2 _10448_ (.A(_05710_),
    .B(_05712_),
    .Y(_05713_));
 sky130_fd_sc_hd__a22o_1 _10449_ (.A1(net500),
    .A2(\core_pipeline.decode_to_execute_csr_data[24] ),
    .B1(\core_pipeline.decode_to_execute_imm_data[24] ),
    .B2(net502),
    .X(_05714_));
 sky130_fd_sc_hd__a21o_4 _10450_ (.A1(_03766_),
    .A2(net433),
    .B1(_05714_),
    .X(_05715_));
 sky130_fd_sc_hd__a22o_1 _10451_ (.A1(net627),
    .A2(\core_pipeline.decode_to_execute_imm_data[24] ),
    .B1(\core_pipeline.decode_to_execute_pc[24] ),
    .B2(net629),
    .X(_05716_));
 sky130_fd_sc_hd__a21o_4 _10452_ (.A1(_03767_),
    .A2(net432),
    .B1(_05716_),
    .X(_05717_));
 sky130_fd_sc_hd__or2_1 _10453_ (.A(_05715_),
    .B(_05717_),
    .X(_05718_));
 sky130_fd_sc_hd__nand2_1 _10454_ (.A(_05715_),
    .B(_05717_),
    .Y(_05719_));
 sky130_fd_sc_hd__and2_1 _10455_ (.A(_05718_),
    .B(_05719_),
    .X(_05720_));
 sky130_fd_sc_hd__a22o_1 _10456_ (.A1(net500),
    .A2(\core_pipeline.decode_to_execute_csr_data[27] ),
    .B1(\core_pipeline.decode_to_execute_imm_data[27] ),
    .B2(net502),
    .X(_05721_));
 sky130_fd_sc_hd__a21o_4 _10457_ (.A1(_03760_),
    .A2(net434),
    .B1(_05721_),
    .X(_05722_));
 sky130_fd_sc_hd__a22o_1 _10458_ (.A1(net627),
    .A2(\core_pipeline.decode_to_execute_imm_data[27] ),
    .B1(\core_pipeline.decode_to_execute_pc[27] ),
    .B2(net629),
    .X(_05723_));
 sky130_fd_sc_hd__a21oi_2 _10459_ (.A1(_03761_),
    .A2(net432),
    .B1(_05723_),
    .Y(_05724_));
 sky130_fd_sc_hd__nand2_1 _10460_ (.A(_05722_),
    .B(net360),
    .Y(_05725_));
 sky130_fd_sc_hd__or2_1 _10461_ (.A(_05722_),
    .B(net360),
    .X(_05726_));
 sky130_fd_sc_hd__nand2_1 _10462_ (.A(_05725_),
    .B(_05726_),
    .Y(_05727_));
 sky130_fd_sc_hd__a22o_1 _10463_ (.A1(net500),
    .A2(\core_pipeline.decode_to_execute_csr_data[25] ),
    .B1(\core_pipeline.decode_to_execute_imm_data[25] ),
    .B2(net502),
    .X(_05728_));
 sky130_fd_sc_hd__a21o_4 _10464_ (.A1(_03753_),
    .A2(net433),
    .B1(_05728_),
    .X(_05729_));
 sky130_fd_sc_hd__a22o_1 _10465_ (.A1(net627),
    .A2(\core_pipeline.decode_to_execute_imm_data[25] ),
    .B1(\core_pipeline.decode_to_execute_pc[25] ),
    .B2(net629),
    .X(_05730_));
 sky130_fd_sc_hd__a21o_4 _10466_ (.A1(_03754_),
    .A2(net431),
    .B1(_05730_),
    .X(_05731_));
 sky130_fd_sc_hd__and2b_1 _10467_ (.A_N(_05731_),
    .B(_05729_),
    .X(_05732_));
 sky130_fd_sc_hd__and2b_1 _10468_ (.A_N(_05729_),
    .B(_05731_),
    .X(_05733_));
 sky130_fd_sc_hd__or2_1 _10469_ (.A(_05732_),
    .B(_05733_),
    .X(_05734_));
 sky130_fd_sc_hd__or4_1 _10470_ (.A(_05713_),
    .B(_05720_),
    .C(_05727_),
    .D(_05734_),
    .X(_05735_));
 sky130_fd_sc_hd__or4_2 _10471_ (.A(_05695_),
    .B(_05700_),
    .C(_05708_),
    .D(_05735_),
    .X(_05736_));
 sky130_fd_sc_hd__a22o_1 _10472_ (.A1(net500),
    .A2(\core_pipeline.decode_to_execute_csr_data[23] ),
    .B1(\core_pipeline.decode_to_execute_imm_data[23] ),
    .B2(net502),
    .X(_05737_));
 sky130_fd_sc_hd__a21oi_4 _10473_ (.A1(_03779_),
    .A2(net433),
    .B1(_05737_),
    .Y(_05738_));
 sky130_fd_sc_hd__a22o_1 _10474_ (.A1(net628),
    .A2(\core_pipeline.decode_to_execute_imm_data[23] ),
    .B1(\core_pipeline.decode_to_execute_pc[23] ),
    .B2(net629),
    .X(_05739_));
 sky130_fd_sc_hd__a21o_4 _10475_ (.A1(_03781_),
    .A2(net432),
    .B1(_05739_),
    .X(_05740_));
 sky130_fd_sc_hd__nand2_1 _10476_ (.A(_05738_),
    .B(_05740_),
    .Y(_05741_));
 sky130_fd_sc_hd__or2_1 _10477_ (.A(_05738_),
    .B(_05740_),
    .X(_05742_));
 sky130_fd_sc_hd__nand2_1 _10478_ (.A(_05741_),
    .B(_05742_),
    .Y(_05743_));
 sky130_fd_sc_hd__a22o_1 _10479_ (.A1(net500),
    .A2(\core_pipeline.decode_to_execute_csr_data[17] ),
    .B1(\core_pipeline.decode_to_execute_imm_data[17] ),
    .B2(net502),
    .X(_05744_));
 sky130_fd_sc_hd__a21oi_4 _10480_ (.A1(_03800_),
    .A2(net433),
    .B1(_05744_),
    .Y(_05745_));
 sky130_fd_sc_hd__and2_2 _10481_ (.A(_03801_),
    .B(net432),
    .X(_05746_));
 sky130_fd_sc_hd__a22o_2 _10482_ (.A1(net628),
    .A2(\core_pipeline.decode_to_execute_imm_data[17] ),
    .B1(\core_pipeline.decode_to_execute_pc[17] ),
    .B2(net630),
    .X(_05747_));
 sky130_fd_sc_hd__or2_4 _10483_ (.A(_05746_),
    .B(_05747_),
    .X(_05748_));
 sky130_fd_sc_hd__xnor2_1 _10484_ (.A(_05745_),
    .B(_05748_),
    .Y(_05749_));
 sky130_fd_sc_hd__a22o_1 _10485_ (.A1(net500),
    .A2(\core_pipeline.decode_to_execute_csr_data[22] ),
    .B1(\core_pipeline.decode_to_execute_imm_data[22] ),
    .B2(net502),
    .X(_05750_));
 sky130_fd_sc_hd__a21o_4 _10486_ (.A1(_03783_),
    .A2(_04474_),
    .B1(_05750_),
    .X(_05751_));
 sky130_fd_sc_hd__a22o_1 _10487_ (.A1(net628),
    .A2(\core_pipeline.decode_to_execute_imm_data[22] ),
    .B1(\core_pipeline.decode_to_execute_pc[22] ),
    .B2(net630),
    .X(_05752_));
 sky130_fd_sc_hd__a21o_4 _10488_ (.A1(_03785_),
    .A2(net431),
    .B1(_05752_),
    .X(_05753_));
 sky130_fd_sc_hd__or2_1 _10489_ (.A(_05751_),
    .B(_05753_),
    .X(_05754_));
 sky130_fd_sc_hd__nand2_1 _10490_ (.A(_05751_),
    .B(_05753_),
    .Y(_05755_));
 sky130_fd_sc_hd__and2_1 _10491_ (.A(_05754_),
    .B(_05755_),
    .X(_05756_));
 sky130_fd_sc_hd__a22o_1 _10492_ (.A1(net500),
    .A2(\core_pipeline.decode_to_execute_csr_data[16] ),
    .B1(\core_pipeline.decode_to_execute_imm_data[16] ),
    .B2(net502),
    .X(_05757_));
 sky130_fd_sc_hd__a21oi_4 _10493_ (.A1(_03803_),
    .A2(_04474_),
    .B1(_05757_),
    .Y(_05758_));
 sky130_fd_sc_hd__a22o_1 _10494_ (.A1(net627),
    .A2(\core_pipeline.decode_to_execute_imm_data[16] ),
    .B1(\core_pipeline.decode_to_execute_pc[16] ),
    .B2(net629),
    .X(_05759_));
 sky130_fd_sc_hd__a21o_4 _10495_ (.A1(_03804_),
    .A2(net431),
    .B1(_05759_),
    .X(_05760_));
 sky130_fd_sc_hd__xnor2_1 _10496_ (.A(_05758_),
    .B(_05760_),
    .Y(_05761_));
 sky130_fd_sc_hd__a22o_1 _10497_ (.A1(net500),
    .A2(\core_pipeline.decode_to_execute_csr_data[21] ),
    .B1(\core_pipeline.decode_to_execute_imm_data[21] ),
    .B2(net502),
    .X(_05762_));
 sky130_fd_sc_hd__a21oi_4 _10498_ (.A1(_03789_),
    .A2(_04474_),
    .B1(_05762_),
    .Y(_05763_));
 sky130_fd_sc_hd__a22o_1 _10499_ (.A1(net628),
    .A2(\core_pipeline.decode_to_execute_imm_data[21] ),
    .B1(\core_pipeline.decode_to_execute_pc[21] ),
    .B2(net630),
    .X(_05764_));
 sky130_fd_sc_hd__a21o_4 _10500_ (.A1(_03790_),
    .A2(net431),
    .B1(_05764_),
    .X(_05765_));
 sky130_fd_sc_hd__inv_2 _10501_ (.A(_05765_),
    .Y(_05766_));
 sky130_fd_sc_hd__nand2_1 _10502_ (.A(_05763_),
    .B(_05765_),
    .Y(_05767_));
 sky130_fd_sc_hd__or2_1 _10503_ (.A(_05763_),
    .B(_05765_),
    .X(_05768_));
 sky130_fd_sc_hd__nand2_1 _10504_ (.A(_05767_),
    .B(_05768_),
    .Y(_05769_));
 sky130_fd_sc_hd__a22o_1 _10505_ (.A1(net500),
    .A2(\core_pipeline.decode_to_execute_csr_data[20] ),
    .B1(\core_pipeline.decode_to_execute_imm_data[20] ),
    .B2(net502),
    .X(_05770_));
 sky130_fd_sc_hd__a21oi_4 _10506_ (.A1(_03786_),
    .A2(net433),
    .B1(_05770_),
    .Y(_05771_));
 sky130_fd_sc_hd__a22o_1 _10507_ (.A1(net628),
    .A2(\core_pipeline.decode_to_execute_imm_data[20] ),
    .B1(\core_pipeline.decode_to_execute_pc[20] ),
    .B2(net630),
    .X(_05772_));
 sky130_fd_sc_hd__a21oi_4 _10508_ (.A1(_03787_),
    .A2(net431),
    .B1(_05772_),
    .Y(_05773_));
 sky130_fd_sc_hd__and2b_1 _10509_ (.A_N(_05771_),
    .B(_05773_),
    .X(_05774_));
 sky130_fd_sc_hd__nand2b_1 _10510_ (.A_N(_05773_),
    .B(_05771_),
    .Y(_05775_));
 sky130_fd_sc_hd__nand2_1 _10511_ (.A(_05771_),
    .B(_05773_),
    .Y(_05776_));
 sky130_fd_sc_hd__nand2b_1 _10512_ (.A_N(_05774_),
    .B(_05775_),
    .Y(_05777_));
 sky130_fd_sc_hd__a22o_1 _10513_ (.A1(net500),
    .A2(\core_pipeline.decode_to_execute_csr_data[18] ),
    .B1(\core_pipeline.decode_to_execute_imm_data[18] ),
    .B2(net502),
    .X(_05778_));
 sky130_fd_sc_hd__a21oi_4 _10514_ (.A1(_03793_),
    .A2(net433),
    .B1(_05778_),
    .Y(_05779_));
 sky130_fd_sc_hd__a22o_1 _10515_ (.A1(\core_pipeline.pipeline_decode.alu_select_a_out[2] ),
    .A2(\core_pipeline.decode_to_execute_imm_data[18] ),
    .B1(\core_pipeline.decode_to_execute_pc[18] ),
    .B2(net630),
    .X(_05780_));
 sky130_fd_sc_hd__a21o_4 _10516_ (.A1(_03794_),
    .A2(net431),
    .B1(_05780_),
    .X(_05781_));
 sky130_fd_sc_hd__nor2_1 _10517_ (.A(_05779_),
    .B(_05781_),
    .Y(_05782_));
 sky130_fd_sc_hd__and2_1 _10518_ (.A(_05779_),
    .B(_05781_),
    .X(_05783_));
 sky130_fd_sc_hd__or2_1 _10519_ (.A(_05782_),
    .B(_05783_),
    .X(_05784_));
 sky130_fd_sc_hd__a22o_1 _10520_ (.A1(net500),
    .A2(\core_pipeline.decode_to_execute_csr_data[19] ),
    .B1(\core_pipeline.decode_to_execute_imm_data[19] ),
    .B2(net502),
    .X(_05785_));
 sky130_fd_sc_hd__a21oi_4 _10521_ (.A1(_03796_),
    .A2(net433),
    .B1(_05785_),
    .Y(_05786_));
 sky130_fd_sc_hd__a22o_1 _10522_ (.A1(net627),
    .A2(\core_pipeline.decode_to_execute_imm_data[19] ),
    .B1(\core_pipeline.decode_to_execute_pc[19] ),
    .B2(net629),
    .X(_05787_));
 sky130_fd_sc_hd__a21oi_4 _10523_ (.A1(_03797_),
    .A2(net431),
    .B1(_05787_),
    .Y(_05788_));
 sky130_fd_sc_hd__and2b_1 _10524_ (.A_N(_05786_),
    .B(_05788_),
    .X(_05789_));
 sky130_fd_sc_hd__nand2b_1 _10525_ (.A_N(_05788_),
    .B(_05786_),
    .Y(_05790_));
 sky130_fd_sc_hd__nand2b_1 _10526_ (.A_N(_05789_),
    .B(_05790_),
    .Y(_05791_));
 sky130_fd_sc_hd__or4_1 _10527_ (.A(_05743_),
    .B(_05756_),
    .C(_05769_),
    .D(_05791_),
    .X(_05792_));
 sky130_fd_sc_hd__or4_1 _10528_ (.A(_05749_),
    .B(_05761_),
    .C(_05777_),
    .D(_05784_),
    .X(_05793_));
 sky130_fd_sc_hd__or2_2 _10529_ (.A(_05792_),
    .B(_05793_),
    .X(_05794_));
 sky130_fd_sc_hd__or3b_1 _10530_ (.A(_05687_),
    .B(_05691_),
    .C_N(_05684_),
    .X(_05795_));
 sky130_fd_sc_hd__and2b_1 _10531_ (.A_N(_05717_),
    .B(_05715_),
    .X(_05796_));
 sky130_fd_sc_hd__nor2_1 _10532_ (.A(_05732_),
    .B(_05796_),
    .Y(_05797_));
 sky130_fd_sc_hd__a21o_1 _10533_ (.A1(_05710_),
    .A2(_05712_),
    .B1(_05733_),
    .X(_05798_));
 sky130_fd_sc_hd__o221a_1 _10534_ (.A1(_05710_),
    .A2(_05712_),
    .B1(_05797_),
    .B2(_05798_),
    .C1(_05725_),
    .X(_05799_));
 sky130_fd_sc_hd__a21bo_1 _10535_ (.A1(_05697_),
    .A2(_05699_),
    .B1_N(_05726_),
    .X(_05800_));
 sky130_fd_sc_hd__o221a_1 _10536_ (.A1(_05697_),
    .A2(_05699_),
    .B1(_05799_),
    .B2(_05800_),
    .C1(_05707_),
    .X(_05801_));
 sky130_fd_sc_hd__or3_1 _10537_ (.A(_05695_),
    .B(_05705_),
    .C(_05801_),
    .X(_05802_));
 sky130_fd_sc_hd__o22a_1 _10538_ (.A1(_05745_),
    .A2(_05748_),
    .B1(_05758_),
    .B2(_05760_),
    .X(_05803_));
 sky130_fd_sc_hd__a211oi_1 _10539_ (.A1(_05745_),
    .A2(_05748_),
    .B1(_05783_),
    .C1(_05803_),
    .Y(_05804_));
 sky130_fd_sc_hd__o311a_1 _10540_ (.A1(_05782_),
    .A2(_05789_),
    .A3(_05804_),
    .B1(_05790_),
    .C1(_05775_),
    .X(_05805_));
 sky130_fd_sc_hd__nor2_1 _10541_ (.A(_05774_),
    .B(_05805_),
    .Y(_05806_));
 sky130_fd_sc_hd__nand2_1 _10542_ (.A(_05768_),
    .B(_05806_),
    .Y(_05807_));
 sky130_fd_sc_hd__and3b_1 _10543_ (.A_N(_05756_),
    .B(_05767_),
    .C(_05807_),
    .X(_05808_));
 sky130_fd_sc_hd__and2b_1 _10544_ (.A_N(_05753_),
    .B(_05751_),
    .X(_05809_));
 sky130_fd_sc_hd__a31o_1 _10545_ (.A1(_05629_),
    .A2(_05682_),
    .A3(_05683_),
    .B1(_05794_),
    .X(_05810_));
 sky130_fd_sc_hd__o21ai_1 _10546_ (.A1(_05808_),
    .A2(_05809_),
    .B1(_05741_),
    .Y(_05811_));
 sky130_fd_sc_hd__a31o_1 _10547_ (.A1(_05742_),
    .A2(_05810_),
    .A3(_05811_),
    .B1(_05736_),
    .X(_05812_));
 sky130_fd_sc_hd__and3_1 _10548_ (.A(_05795_),
    .B(_05802_),
    .C(_05812_),
    .X(_05813_));
 sky130_fd_sc_hd__xnor2_1 _10549_ (.A(net395),
    .B(_04517_),
    .Y(_05814_));
 sky130_fd_sc_hd__xnor2_1 _10550_ (.A(net384),
    .B(_04511_),
    .Y(_05815_));
 sky130_fd_sc_hd__nand2_1 _10551_ (.A(_04496_),
    .B(_04504_),
    .Y(_05816_));
 sky130_fd_sc_hd__or2_1 _10552_ (.A(net379),
    .B(_04502_),
    .X(_05817_));
 sky130_fd_sc_hd__nand2_1 _10553_ (.A(net379),
    .B(_04502_),
    .Y(_05818_));
 sky130_fd_sc_hd__and2_1 _10554_ (.A(_05817_),
    .B(_05818_),
    .X(_05819_));
 sky130_fd_sc_hd__or4_1 _10555_ (.A(_05674_),
    .B(_05675_),
    .C(_05816_),
    .D(_05819_),
    .X(_05820_));
 sky130_fd_sc_hd__or4_2 _10556_ (.A(_05664_),
    .B(_05814_),
    .C(_05815_),
    .D(_05820_),
    .X(_05821_));
 sky130_fd_sc_hd__or3_1 _10557_ (.A(_05631_),
    .B(_05736_),
    .C(_05821_),
    .X(_05822_));
 sky130_fd_sc_hd__nor3_2 _10558_ (.A(_05655_),
    .B(_05794_),
    .C(_05822_),
    .Y(_05823_));
 sky130_fd_sc_hd__a21oi_1 _10559_ (.A1(_05616_),
    .A2(_05813_),
    .B1(_05823_),
    .Y(_05824_));
 sky130_fd_sc_hd__mux2_1 _10560_ (.A0(\core_pipeline.pipeline_execute.ex_alu.result_sltu[0] ),
    .A1(_05824_),
    .S(_05610_),
    .X(_01354_));
 sky130_fd_sc_hd__nor3_4 _10561_ (.A(\core_pipeline.execute_to_memory_exception ),
    .B(_03426_),
    .C(_03428_),
    .Y(_05825_));
 sky130_fd_sc_hd__o31a_2 _10562_ (.A1(\core_pipeline.execute_to_memory_exception ),
    .A2(_03508_),
    .A3(_03509_),
    .B1(net446),
    .X(_05826_));
 sky130_fd_sc_hd__and2b_1 _10563_ (.A_N(_05825_),
    .B(_05826_),
    .X(_05827_));
 sky130_fd_sc_hd__inv_2 _10564_ (.A(_05827_),
    .Y(_05828_));
 sky130_fd_sc_hd__o22a_1 _10565_ (.A1(\core_pipeline.memory_to_writeback_exception ),
    .A2(net454),
    .B1(_05828_),
    .B2(\core_pipeline.execute_to_memory_exception ),
    .X(_01355_));
 sky130_fd_sc_hd__or2_1 _10566_ (.A(\core_pipeline.execute_to_memory_wfi ),
    .B(_03431_),
    .X(_01356_));
 sky130_fd_sc_hd__nor2_2 _10567_ (.A(\core_pipeline.pipeline_execute.ex_alu.old_function[1] ),
    .B(\core_pipeline.pipeline_execute.ex_alu.old_function[0] ),
    .Y(_05829_));
 sky130_fd_sc_hd__and2_2 _10568_ (.A(_03420_),
    .B(net423),
    .X(_05830_));
 sky130_fd_sc_hd__nand2_2 _10569_ (.A(_03420_),
    .B(net423),
    .Y(_05831_));
 sky130_fd_sc_hd__mux2_1 _10570_ (.A0(\core_pipeline.pipeline_execute.ex_alu.result_slt[0] ),
    .A1(\core_pipeline.pipeline_execute.ex_alu.result_sltu[0] ),
    .S(\core_pipeline.pipeline_execute.ex_alu.old_function[0] ),
    .X(_05832_));
 sky130_fd_sc_hd__or3b_1 _10571_ (.A(\core_pipeline.pipeline_execute.ex_alu.old_function[1] ),
    .B(\core_pipeline.pipeline_execute.ex_alu.result_sll[0] ),
    .C_N(\core_pipeline.pipeline_execute.ex_alu.old_function[0] ),
    .X(_05833_));
 sky130_fd_sc_hd__o211a_1 _10572_ (.A1(_03421_),
    .A2(_05832_),
    .B1(_05833_),
    .C1(_03420_),
    .X(_05834_));
 sky130_fd_sc_hd__and3_2 _10573_ (.A(\core_pipeline.pipeline_execute.ex_alu.old_function[2] ),
    .B(\core_pipeline.pipeline_execute.ex_alu.old_function[1] ),
    .C(\core_pipeline.pipeline_execute.ex_alu.old_function[0] ),
    .X(_05835_));
 sky130_fd_sc_hd__a32o_1 _10574_ (.A1(\core_pipeline.pipeline_execute.ex_alu.old_function[2] ),
    .A2(\core_pipeline.pipeline_execute.ex_alu.result_xor[0] ),
    .A3(net423),
    .B1(net421),
    .B2(\core_pipeline.pipeline_execute.ex_alu.result_and_clr[0] ),
    .X(_05836_));
 sky130_fd_sc_hd__and3_2 _10575_ (.A(\core_pipeline.pipeline_execute.ex_alu.old_function[2] ),
    .B(_03421_),
    .C(\core_pipeline.pipeline_execute.ex_alu.old_function[0] ),
    .X(_05837_));
 sky130_fd_sc_hd__and3b_2 _10576_ (.A_N(\core_pipeline.pipeline_execute.ex_alu.old_function[0] ),
    .B(\core_pipeline.pipeline_execute.ex_alu.old_function[1] ),
    .C(\core_pipeline.pipeline_execute.ex_alu.old_function[2] ),
    .X(_05838_));
 sky130_fd_sc_hd__a221o_1 _10577_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_srl_sra[0] ),
    .A2(net355),
    .B1(net419),
    .B2(\core_pipeline.pipeline_execute.ex_alu.result_or[0] ),
    .C1(_05836_),
    .X(_05839_));
 sky130_fd_sc_hd__o22a_1 _10578_ (.A1(net493),
    .A2(net357),
    .B1(_05834_),
    .B2(_05839_),
    .X(_05840_));
 sky130_fd_sc_hd__mux2_1 _10579_ (.A0(\core_pipeline.memory_to_writeback_alu_data[0] ),
    .A1(_05840_),
    .S(net448),
    .X(_01357_));
 sky130_fd_sc_hd__a221o_1 _10580_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_xor[1] ),
    .A2(net423),
    .B1(net355),
    .B2(\core_pipeline.pipeline_execute.ex_alu.result_srl_sra[1] ),
    .C1(net359),
    .X(_05841_));
 sky130_fd_sc_hd__and3_1 _10581_ (.A(_03420_),
    .B(_03421_),
    .C(\core_pipeline.pipeline_execute.ex_alu.old_function[0] ),
    .X(_05842_));
 sky130_fd_sc_hd__a22o_1 _10582_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_and_clr[1] ),
    .A2(net421),
    .B1(net419),
    .B2(\core_pipeline.pipeline_execute.ex_alu.result_or[1] ),
    .X(_05843_));
 sky130_fd_sc_hd__a21o_1 _10583_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_sll[1] ),
    .A2(net353),
    .B1(_05843_),
    .X(_05844_));
 sky130_fd_sc_hd__o22a_4 _10584_ (.A1(net492),
    .A2(net357),
    .B1(_05841_),
    .B2(_05844_),
    .X(_05845_));
 sky130_fd_sc_hd__mux2_1 _10585_ (.A0(\core_pipeline.memory_to_writeback_alu_data[1] ),
    .A1(_05845_),
    .S(net446),
    .X(_01358_));
 sky130_fd_sc_hd__a221o_1 _10586_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_xor[2] ),
    .A2(net423),
    .B1(net355),
    .B2(\core_pipeline.pipeline_execute.ex_alu.result_srl_sra[2] ),
    .C1(net359),
    .X(_05846_));
 sky130_fd_sc_hd__a22o_1 _10587_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_and_clr[2] ),
    .A2(net421),
    .B1(net419),
    .B2(\core_pipeline.pipeline_execute.ex_alu.result_or[2] ),
    .X(_05847_));
 sky130_fd_sc_hd__a21o_1 _10588_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_sll[2] ),
    .A2(net353),
    .B1(_05847_),
    .X(_05848_));
 sky130_fd_sc_hd__o22a_4 _10589_ (.A1(\core_busio.mem_address[2] ),
    .A2(net357),
    .B1(_05846_),
    .B2(_05848_),
    .X(_05849_));
 sky130_fd_sc_hd__mux2_1 _10590_ (.A0(\core_pipeline.memory_to_writeback_alu_data[2] ),
    .A1(_05849_),
    .S(net454),
    .X(_01359_));
 sky130_fd_sc_hd__a221o_1 _10591_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_xor[3] ),
    .A2(net423),
    .B1(net419),
    .B2(\core_pipeline.pipeline_execute.ex_alu.result_or[3] ),
    .C1(net359),
    .X(_05850_));
 sky130_fd_sc_hd__and2_1 _10592_ (.A(\core_pipeline.pipeline_execute.ex_alu.result_sll[3] ),
    .B(net353),
    .X(_05851_));
 sky130_fd_sc_hd__a22o_1 _10593_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_and_clr[3] ),
    .A2(net421),
    .B1(net355),
    .B2(\core_pipeline.pipeline_execute.ex_alu.result_srl_sra[3] ),
    .X(_05852_));
 sky130_fd_sc_hd__o32a_2 _10594_ (.A1(_05850_),
    .A2(_05851_),
    .A3(_05852_),
    .B1(net357),
    .B2(\core_busio.mem_address[3] ),
    .X(_05853_));
 sky130_fd_sc_hd__mux2_1 _10595_ (.A0(\core_pipeline.memory_to_writeback_alu_data[3] ),
    .A1(_05853_),
    .S(net448),
    .X(_01360_));
 sky130_fd_sc_hd__a221o_1 _10596_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_xor[4] ),
    .A2(net423),
    .B1(net355),
    .B2(\core_pipeline.pipeline_execute.ex_alu.result_srl_sra[4] ),
    .C1(net359),
    .X(_05854_));
 sky130_fd_sc_hd__a22o_1 _10597_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_and_clr[4] ),
    .A2(net421),
    .B1(net419),
    .B2(\core_pipeline.pipeline_execute.ex_alu.result_or[4] ),
    .X(_05855_));
 sky130_fd_sc_hd__a21o_1 _10598_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_sll[4] ),
    .A2(net353),
    .B1(_05855_),
    .X(_05856_));
 sky130_fd_sc_hd__o22a_2 _10599_ (.A1(\core_busio.mem_address[4] ),
    .A2(net357),
    .B1(_05854_),
    .B2(_05856_),
    .X(_05857_));
 sky130_fd_sc_hd__mux2_1 _10600_ (.A0(\core_pipeline.memory_to_writeback_alu_data[4] ),
    .A1(_05857_),
    .S(net448),
    .X(_01361_));
 sky130_fd_sc_hd__a221o_1 _10601_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_xor[5] ),
    .A2(net423),
    .B1(net419),
    .B2(\core_pipeline.pipeline_execute.ex_alu.result_or[5] ),
    .C1(net359),
    .X(_05858_));
 sky130_fd_sc_hd__and2_1 _10602_ (.A(\core_pipeline.pipeline_execute.ex_alu.result_sll[5] ),
    .B(net353),
    .X(_05859_));
 sky130_fd_sc_hd__a22o_1 _10603_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_and_clr[5] ),
    .A2(net421),
    .B1(net355),
    .B2(\core_pipeline.pipeline_execute.ex_alu.result_srl_sra[5] ),
    .X(_05860_));
 sky130_fd_sc_hd__o32a_4 _10604_ (.A1(_05858_),
    .A2(_05859_),
    .A3(_05860_),
    .B1(net357),
    .B2(\core_busio.mem_address[5] ),
    .X(_05861_));
 sky130_fd_sc_hd__mux2_1 _10605_ (.A0(\core_pipeline.memory_to_writeback_alu_data[5] ),
    .A1(_05861_),
    .S(net446),
    .X(_01362_));
 sky130_fd_sc_hd__and2_1 _10606_ (.A(\core_pipeline.pipeline_execute.ex_alu.result_and_clr[6] ),
    .B(net421),
    .X(_05862_));
 sky130_fd_sc_hd__a221o_1 _10607_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_xor[6] ),
    .A2(net423),
    .B1(net353),
    .B2(\core_pipeline.pipeline_execute.ex_alu.result_sll[6] ),
    .C1(net359),
    .X(_05863_));
 sky130_fd_sc_hd__a221o_2 _10608_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_srl_sra[6] ),
    .A2(net355),
    .B1(net419),
    .B2(\core_pipeline.pipeline_execute.ex_alu.result_or[6] ),
    .C1(_05863_),
    .X(_05864_));
 sky130_fd_sc_hd__o22a_2 _10609_ (.A1(\core_busio.mem_address[6] ),
    .A2(net357),
    .B1(_05862_),
    .B2(_05864_),
    .X(_05865_));
 sky130_fd_sc_hd__mux2_1 _10610_ (.A0(\core_pipeline.memory_to_writeback_alu_data[6] ),
    .A1(_05865_),
    .S(net447),
    .X(_01363_));
 sky130_fd_sc_hd__a221o_1 _10611_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_xor[7] ),
    .A2(net423),
    .B1(net355),
    .B2(\core_pipeline.pipeline_execute.ex_alu.result_srl_sra[7] ),
    .C1(net359),
    .X(_05866_));
 sky130_fd_sc_hd__a22o_1 _10612_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_and_clr[7] ),
    .A2(net421),
    .B1(net419),
    .B2(\core_pipeline.pipeline_execute.ex_alu.result_or[7] ),
    .X(_05867_));
 sky130_fd_sc_hd__a21o_1 _10613_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_sll[7] ),
    .A2(net353),
    .B1(_05867_),
    .X(_05868_));
 sky130_fd_sc_hd__o22a_1 _10614_ (.A1(\core_busio.mem_address[7] ),
    .A2(net357),
    .B1(_05866_),
    .B2(_05868_),
    .X(_05869_));
 sky130_fd_sc_hd__mux2_1 _10615_ (.A0(\core_pipeline.memory_to_writeback_alu_data[7] ),
    .A1(_05869_),
    .S(net448),
    .X(_01364_));
 sky130_fd_sc_hd__and2_1 _10616_ (.A(\core_pipeline.pipeline_execute.ex_alu.result_and_clr[8] ),
    .B(net420),
    .X(_05870_));
 sky130_fd_sc_hd__a221o_1 _10617_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_xor[8] ),
    .A2(net422),
    .B1(net352),
    .B2(\core_pipeline.pipeline_execute.ex_alu.result_sll[8] ),
    .C1(net358),
    .X(_05871_));
 sky130_fd_sc_hd__a221o_1 _10618_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_srl_sra[8] ),
    .A2(net354),
    .B1(net418),
    .B2(\core_pipeline.pipeline_execute.ex_alu.result_or[8] ),
    .C1(_05871_),
    .X(_05872_));
 sky130_fd_sc_hd__o22a_2 _10619_ (.A1(\core_busio.mem_address[8] ),
    .A2(net356),
    .B1(_05870_),
    .B2(_05872_),
    .X(_05873_));
 sky130_fd_sc_hd__mux2_1 _10620_ (.A0(\core_pipeline.memory_to_writeback_alu_data[8] ),
    .A1(_05873_),
    .S(net450),
    .X(_01365_));
 sky130_fd_sc_hd__and2_1 _10621_ (.A(\core_pipeline.pipeline_execute.ex_alu.result_and_clr[9] ),
    .B(net420),
    .X(_05874_));
 sky130_fd_sc_hd__a221o_1 _10622_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_xor[9] ),
    .A2(net422),
    .B1(net352),
    .B2(\core_pipeline.pipeline_execute.ex_alu.result_sll[9] ),
    .C1(net358),
    .X(_05875_));
 sky130_fd_sc_hd__a221o_1 _10623_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_srl_sra[9] ),
    .A2(net354),
    .B1(net418),
    .B2(\core_pipeline.pipeline_execute.ex_alu.result_or[9] ),
    .C1(_05875_),
    .X(_05876_));
 sky130_fd_sc_hd__o22a_4 _10624_ (.A1(\core_busio.mem_address[9] ),
    .A2(net356),
    .B1(_05874_),
    .B2(_05876_),
    .X(_05877_));
 sky130_fd_sc_hd__mux2_1 _10625_ (.A0(\core_pipeline.memory_to_writeback_alu_data[9] ),
    .A1(_05877_),
    .S(net450),
    .X(_01366_));
 sky130_fd_sc_hd__and2_1 _10626_ (.A(\core_pipeline.pipeline_execute.ex_alu.result_and_clr[10] ),
    .B(net420),
    .X(_05878_));
 sky130_fd_sc_hd__a221o_1 _10627_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_xor[10] ),
    .A2(net422),
    .B1(net352),
    .B2(\core_pipeline.pipeline_execute.ex_alu.result_sll[10] ),
    .C1(net358),
    .X(_05879_));
 sky130_fd_sc_hd__a221o_1 _10628_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_srl_sra[10] ),
    .A2(net354),
    .B1(net418),
    .B2(\core_pipeline.pipeline_execute.ex_alu.result_or[10] ),
    .C1(_05879_),
    .X(_05880_));
 sky130_fd_sc_hd__o22a_2 _10629_ (.A1(\core_busio.mem_address[10] ),
    .A2(net356),
    .B1(_05878_),
    .B2(_05880_),
    .X(_05881_));
 sky130_fd_sc_hd__mux2_1 _10630_ (.A0(\core_pipeline.memory_to_writeback_alu_data[10] ),
    .A1(_05881_),
    .S(net453),
    .X(_01367_));
 sky130_fd_sc_hd__a221o_1 _10631_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_xor[11] ),
    .A2(net422),
    .B1(net418),
    .B2(\core_pipeline.pipeline_execute.ex_alu.result_or[11] ),
    .C1(net358),
    .X(_05882_));
 sky130_fd_sc_hd__and2_1 _10632_ (.A(\core_pipeline.pipeline_execute.ex_alu.result_sll[11] ),
    .B(net352),
    .X(_05883_));
 sky130_fd_sc_hd__a22o_1 _10633_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_and_clr[11] ),
    .A2(net420),
    .B1(net354),
    .B2(\core_pipeline.pipeline_execute.ex_alu.result_srl_sra[11] ),
    .X(_05884_));
 sky130_fd_sc_hd__o32a_4 _10634_ (.A1(_05882_),
    .A2(_05883_),
    .A3(_05884_),
    .B1(net356),
    .B2(\core_busio.mem_address[11] ),
    .X(_05885_));
 sky130_fd_sc_hd__mux2_1 _10635_ (.A0(\core_pipeline.memory_to_writeback_alu_data[11] ),
    .A1(_05885_),
    .S(net449),
    .X(_01368_));
 sky130_fd_sc_hd__and2_1 _10636_ (.A(\core_pipeline.pipeline_execute.ex_alu.result_and_clr[12] ),
    .B(net420),
    .X(_05886_));
 sky130_fd_sc_hd__a221o_1 _10637_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_xor[12] ),
    .A2(net422),
    .B1(net352),
    .B2(\core_pipeline.pipeline_execute.ex_alu.result_sll[12] ),
    .C1(net358),
    .X(_05887_));
 sky130_fd_sc_hd__a221o_2 _10638_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_srl_sra[12] ),
    .A2(net354),
    .B1(net418),
    .B2(\core_pipeline.pipeline_execute.ex_alu.result_or[12] ),
    .C1(_05887_),
    .X(_05888_));
 sky130_fd_sc_hd__o22a_2 _10639_ (.A1(\core_busio.mem_address[12] ),
    .A2(net357),
    .B1(_05886_),
    .B2(_05888_),
    .X(_05889_));
 sky130_fd_sc_hd__mux2_1 _10640_ (.A0(\core_pipeline.memory_to_writeback_alu_data[12] ),
    .A1(_05889_),
    .S(net449),
    .X(_01369_));
 sky130_fd_sc_hd__and2_1 _10641_ (.A(\core_pipeline.pipeline_execute.ex_alu.result_and_clr[13] ),
    .B(net420),
    .X(_05890_));
 sky130_fd_sc_hd__a221o_1 _10642_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_xor[13] ),
    .A2(net422),
    .B1(net353),
    .B2(\core_pipeline.pipeline_execute.ex_alu.result_sll[13] ),
    .C1(net358),
    .X(_05891_));
 sky130_fd_sc_hd__a221o_1 _10643_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_srl_sra[13] ),
    .A2(net354),
    .B1(net418),
    .B2(\core_pipeline.pipeline_execute.ex_alu.result_or[13] ),
    .C1(_05891_),
    .X(_05892_));
 sky130_fd_sc_hd__o22a_2 _10644_ (.A1(\core_busio.mem_address[13] ),
    .A2(net356),
    .B1(_05890_),
    .B2(_05892_),
    .X(_05893_));
 sky130_fd_sc_hd__mux2_1 _10645_ (.A0(\core_pipeline.memory_to_writeback_alu_data[13] ),
    .A1(_05893_),
    .S(net449),
    .X(_01370_));
 sky130_fd_sc_hd__and2_1 _10646_ (.A(\core_pipeline.pipeline_execute.ex_alu.result_and_clr[14] ),
    .B(net420),
    .X(_05894_));
 sky130_fd_sc_hd__a221o_1 _10647_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_xor[14] ),
    .A2(net422),
    .B1(net352),
    .B2(\core_pipeline.pipeline_execute.ex_alu.result_sll[14] ),
    .C1(net358),
    .X(_05895_));
 sky130_fd_sc_hd__a221o_2 _10648_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_srl_sra[14] ),
    .A2(net354),
    .B1(net418),
    .B2(\core_pipeline.pipeline_execute.ex_alu.result_or[14] ),
    .C1(_05895_),
    .X(_05896_));
 sky130_fd_sc_hd__o22a_1 _10649_ (.A1(\core_busio.mem_address[14] ),
    .A2(net357),
    .B1(_05894_),
    .B2(_05896_),
    .X(_05897_));
 sky130_fd_sc_hd__mux2_1 _10650_ (.A0(\core_pipeline.memory_to_writeback_alu_data[14] ),
    .A1(_05897_),
    .S(net449),
    .X(_01371_));
 sky130_fd_sc_hd__a221o_1 _10651_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_xor[15] ),
    .A2(net422),
    .B1(net418),
    .B2(\core_pipeline.pipeline_execute.ex_alu.result_or[15] ),
    .C1(net359),
    .X(_05898_));
 sky130_fd_sc_hd__and2_1 _10652_ (.A(\core_pipeline.pipeline_execute.ex_alu.result_sll[15] ),
    .B(net352),
    .X(_05899_));
 sky130_fd_sc_hd__a22o_1 _10653_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_and_clr[15] ),
    .A2(net421),
    .B1(net354),
    .B2(\core_pipeline.pipeline_execute.ex_alu.result_srl_sra[15] ),
    .X(_05900_));
 sky130_fd_sc_hd__o32a_2 _10654_ (.A1(_05898_),
    .A2(_05899_),
    .A3(_05900_),
    .B1(net356),
    .B2(\core_busio.mem_address[15] ),
    .X(_05901_));
 sky130_fd_sc_hd__mux2_1 _10655_ (.A0(\core_pipeline.memory_to_writeback_alu_data[15] ),
    .A1(_05901_),
    .S(net450),
    .X(_01372_));
 sky130_fd_sc_hd__and2_1 _10656_ (.A(\core_pipeline.pipeline_execute.ex_alu.result_and_clr[16] ),
    .B(net420),
    .X(_05902_));
 sky130_fd_sc_hd__a221o_1 _10657_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_xor[16] ),
    .A2(net423),
    .B1(net352),
    .B2(\core_pipeline.pipeline_execute.ex_alu.result_sll[16] ),
    .C1(net359),
    .X(_05903_));
 sky130_fd_sc_hd__a221o_1 _10658_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_srl_sra[16] ),
    .A2(net355),
    .B1(net418),
    .B2(\core_pipeline.pipeline_execute.ex_alu.result_or[16] ),
    .C1(_05903_),
    .X(_05904_));
 sky130_fd_sc_hd__o22a_2 _10659_ (.A1(\core_busio.mem_address[16] ),
    .A2(net357),
    .B1(_05902_),
    .B2(_05904_),
    .X(_05905_));
 sky130_fd_sc_hd__mux2_1 _10660_ (.A0(\core_pipeline.memory_to_writeback_alu_data[16] ),
    .A1(_05905_),
    .S(net450),
    .X(_01373_));
 sky130_fd_sc_hd__a221o_1 _10661_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_xor[17] ),
    .A2(net423),
    .B1(net355),
    .B2(\core_pipeline.pipeline_execute.ex_alu.result_srl_sra[17] ),
    .C1(net359),
    .X(_05906_));
 sky130_fd_sc_hd__a22o_1 _10662_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_and_clr[17] ),
    .A2(net420),
    .B1(net418),
    .B2(\core_pipeline.pipeline_execute.ex_alu.result_or[17] ),
    .X(_05907_));
 sky130_fd_sc_hd__a21o_1 _10663_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_sll[17] ),
    .A2(net353),
    .B1(_05907_),
    .X(_05908_));
 sky130_fd_sc_hd__o22a_4 _10664_ (.A1(\core_busio.mem_address[17] ),
    .A2(net356),
    .B1(_05906_),
    .B2(_05908_),
    .X(_05909_));
 sky130_fd_sc_hd__mux2_1 _10665_ (.A0(\core_pipeline.memory_to_writeback_alu_data[17] ),
    .A1(_05909_),
    .S(net457),
    .X(_01374_));
 sky130_fd_sc_hd__and2_1 _10666_ (.A(\core_pipeline.pipeline_execute.ex_alu.result_and_clr[18] ),
    .B(net420),
    .X(_05910_));
 sky130_fd_sc_hd__a221o_1 _10667_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_xor[18] ),
    .A2(net422),
    .B1(net353),
    .B2(\core_pipeline.pipeline_execute.ex_alu.result_sll[18] ),
    .C1(net358),
    .X(_05911_));
 sky130_fd_sc_hd__a221o_1 _10668_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_srl_sra[18] ),
    .A2(net354),
    .B1(net418),
    .B2(\core_pipeline.pipeline_execute.ex_alu.result_or[18] ),
    .C1(_05911_),
    .X(_05912_));
 sky130_fd_sc_hd__o22a_4 _10669_ (.A1(\core_busio.mem_address[18] ),
    .A2(net356),
    .B1(_05910_),
    .B2(_05912_),
    .X(_05913_));
 sky130_fd_sc_hd__mux2_1 _10670_ (.A0(\core_pipeline.memory_to_writeback_alu_data[18] ),
    .A1(_05913_),
    .S(net456),
    .X(_01375_));
 sky130_fd_sc_hd__and2_1 _10671_ (.A(\core_pipeline.pipeline_execute.ex_alu.result_and_clr[19] ),
    .B(net420),
    .X(_05914_));
 sky130_fd_sc_hd__a221o_1 _10672_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_xor[19] ),
    .A2(net422),
    .B1(net352),
    .B2(\core_pipeline.pipeline_execute.ex_alu.result_sll[19] ),
    .C1(net358),
    .X(_05915_));
 sky130_fd_sc_hd__a221o_2 _10673_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_srl_sra[19] ),
    .A2(net354),
    .B1(net418),
    .B2(\core_pipeline.pipeline_execute.ex_alu.result_or[19] ),
    .C1(_05915_),
    .X(_05916_));
 sky130_fd_sc_hd__o22a_4 _10674_ (.A1(\core_busio.mem_address[19] ),
    .A2(net356),
    .B1(_05914_),
    .B2(_05916_),
    .X(_05917_));
 sky130_fd_sc_hd__mux2_1 _10675_ (.A0(\core_pipeline.memory_to_writeback_alu_data[19] ),
    .A1(_05917_),
    .S(net456),
    .X(_01376_));
 sky130_fd_sc_hd__and2_1 _10676_ (.A(\core_pipeline.pipeline_execute.ex_alu.result_and_clr[20] ),
    .B(net420),
    .X(_05918_));
 sky130_fd_sc_hd__a221o_1 _10677_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_xor[20] ),
    .A2(net422),
    .B1(net352),
    .B2(\core_pipeline.pipeline_execute.ex_alu.result_sll[20] ),
    .C1(net358),
    .X(_05919_));
 sky130_fd_sc_hd__a221o_2 _10678_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_srl_sra[20] ),
    .A2(net354),
    .B1(net418),
    .B2(\core_pipeline.pipeline_execute.ex_alu.result_or[20] ),
    .C1(_05919_),
    .X(_05920_));
 sky130_fd_sc_hd__o22a_4 _10679_ (.A1(\core_busio.mem_address[20] ),
    .A2(net356),
    .B1(_05918_),
    .B2(_05920_),
    .X(_05921_));
 sky130_fd_sc_hd__mux2_1 _10680_ (.A0(\core_pipeline.memory_to_writeback_alu_data[20] ),
    .A1(_05921_),
    .S(net456),
    .X(_01377_));
 sky130_fd_sc_hd__a221o_1 _10681_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_xor[21] ),
    .A2(_05829_),
    .B1(net354),
    .B2(\core_pipeline.pipeline_execute.ex_alu.result_srl_sra[21] ),
    .C1(net358),
    .X(_05922_));
 sky130_fd_sc_hd__a22o_1 _10682_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_and_clr[21] ),
    .A2(net421),
    .B1(net419),
    .B2(\core_pipeline.pipeline_execute.ex_alu.result_or[21] ),
    .X(_05923_));
 sky130_fd_sc_hd__a21o_1 _10683_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_sll[21] ),
    .A2(net352),
    .B1(_05923_),
    .X(_05924_));
 sky130_fd_sc_hd__o22a_4 _10684_ (.A1(\core_busio.mem_address[21] ),
    .A2(net356),
    .B1(_05922_),
    .B2(_05924_),
    .X(_05925_));
 sky130_fd_sc_hd__mux2_1 _10685_ (.A0(\core_pipeline.memory_to_writeback_alu_data[21] ),
    .A1(_05925_),
    .S(net456),
    .X(_01378_));
 sky130_fd_sc_hd__and2_1 _10686_ (.A(\core_pipeline.pipeline_execute.ex_alu.result_and_clr[22] ),
    .B(net420),
    .X(_05926_));
 sky130_fd_sc_hd__a221o_1 _10687_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_xor[22] ),
    .A2(net422),
    .B1(net352),
    .B2(\core_pipeline.pipeline_execute.ex_alu.result_sll[22] ),
    .C1(net358),
    .X(_05927_));
 sky130_fd_sc_hd__a221o_1 _10688_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_srl_sra[22] ),
    .A2(net354),
    .B1(net418),
    .B2(\core_pipeline.pipeline_execute.ex_alu.result_or[22] ),
    .C1(_05927_),
    .X(_05928_));
 sky130_fd_sc_hd__o22a_2 _10689_ (.A1(\core_busio.mem_address[22] ),
    .A2(net356),
    .B1(_05926_),
    .B2(_05928_),
    .X(_05929_));
 sky130_fd_sc_hd__mux2_1 _10690_ (.A0(\core_pipeline.memory_to_writeback_alu_data[22] ),
    .A1(_05929_),
    .S(net456),
    .X(_01379_));
 sky130_fd_sc_hd__a221o_1 _10691_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_xor[23] ),
    .A2(net422),
    .B1(net354),
    .B2(\core_pipeline.pipeline_execute.ex_alu.result_srl_sra[23] ),
    .C1(net358),
    .X(_05930_));
 sky130_fd_sc_hd__a22o_1 _10692_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_and_clr[23] ),
    .A2(net421),
    .B1(net419),
    .B2(\core_pipeline.pipeline_execute.ex_alu.result_or[23] ),
    .X(_05931_));
 sky130_fd_sc_hd__a21o_1 _10693_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_sll[23] ),
    .A2(net353),
    .B1(_05931_),
    .X(_05932_));
 sky130_fd_sc_hd__o22a_2 _10694_ (.A1(\core_busio.mem_address[23] ),
    .A2(net356),
    .B1(_05930_),
    .B2(_05932_),
    .X(_05933_));
 sky130_fd_sc_hd__mux2_1 _10695_ (.A0(\core_pipeline.memory_to_writeback_alu_data[23] ),
    .A1(_05933_),
    .S(net452),
    .X(_01380_));
 sky130_fd_sc_hd__and2_1 _10696_ (.A(\core_pipeline.pipeline_execute.ex_alu.result_and_clr[24] ),
    .B(net421),
    .X(_05934_));
 sky130_fd_sc_hd__a221o_1 _10697_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_xor[24] ),
    .A2(net422),
    .B1(net352),
    .B2(\core_pipeline.pipeline_execute.ex_alu.result_sll[24] ),
    .C1(net358),
    .X(_05935_));
 sky130_fd_sc_hd__a221o_1 _10698_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_srl_sra[24] ),
    .A2(net355),
    .B1(net419),
    .B2(\core_pipeline.pipeline_execute.ex_alu.result_or[24] ),
    .C1(_05935_),
    .X(_05936_));
 sky130_fd_sc_hd__o22a_2 _10699_ (.A1(\core_busio.mem_address[24] ),
    .A2(net356),
    .B1(_05934_),
    .B2(_05936_),
    .X(_05937_));
 sky130_fd_sc_hd__mux2_1 _10700_ (.A0(\core_pipeline.memory_to_writeback_alu_data[24] ),
    .A1(_05937_),
    .S(net450),
    .X(_01381_));
 sky130_fd_sc_hd__and2_1 _10701_ (.A(\core_pipeline.pipeline_execute.ex_alu.result_and_clr[25] ),
    .B(net420),
    .X(_05938_));
 sky130_fd_sc_hd__a221o_1 _10702_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_xor[25] ),
    .A2(net422),
    .B1(net352),
    .B2(\core_pipeline.pipeline_execute.ex_alu.result_sll[25] ),
    .C1(net358),
    .X(_05939_));
 sky130_fd_sc_hd__a221o_2 _10703_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_srl_sra[25] ),
    .A2(net355),
    .B1(net419),
    .B2(\core_pipeline.pipeline_execute.ex_alu.result_or[25] ),
    .C1(_05939_),
    .X(_05940_));
 sky130_fd_sc_hd__o22a_1 _10704_ (.A1(\core_busio.mem_address[25] ),
    .A2(net356),
    .B1(_05938_),
    .B2(_05940_),
    .X(_05941_));
 sky130_fd_sc_hd__mux2_1 _10705_ (.A0(\core_pipeline.memory_to_writeback_alu_data[25] ),
    .A1(_05941_),
    .S(net450),
    .X(_01382_));
 sky130_fd_sc_hd__and2_1 _10706_ (.A(\core_pipeline.pipeline_execute.ex_alu.result_and_clr[26] ),
    .B(net420),
    .X(_05942_));
 sky130_fd_sc_hd__a221o_1 _10707_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_xor[26] ),
    .A2(net422),
    .B1(net352),
    .B2(\core_pipeline.pipeline_execute.ex_alu.result_sll[26] ),
    .C1(net358),
    .X(_05943_));
 sky130_fd_sc_hd__a221o_1 _10708_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_srl_sra[26] ),
    .A2(net354),
    .B1(net418),
    .B2(\core_pipeline.pipeline_execute.ex_alu.result_or[26] ),
    .C1(_05943_),
    .X(_05944_));
 sky130_fd_sc_hd__o22a_1 _10709_ (.A1(\core_busio.mem_address[26] ),
    .A2(net356),
    .B1(_05942_),
    .B2(_05944_),
    .X(_05945_));
 sky130_fd_sc_hd__mux2_1 _10710_ (.A0(\core_pipeline.memory_to_writeback_alu_data[26] ),
    .A1(_05945_),
    .S(net450),
    .X(_01383_));
 sky130_fd_sc_hd__a221o_1 _10711_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_xor[27] ),
    .A2(net423),
    .B1(net354),
    .B2(\core_pipeline.pipeline_execute.ex_alu.result_srl_sra[27] ),
    .C1(net359),
    .X(_05946_));
 sky130_fd_sc_hd__a22o_1 _10712_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_and_clr[27] ),
    .A2(net420),
    .B1(net419),
    .B2(\core_pipeline.pipeline_execute.ex_alu.result_or[27] ),
    .X(_05947_));
 sky130_fd_sc_hd__a21o_1 _10713_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_sll[27] ),
    .A2(net352),
    .B1(_05947_),
    .X(_05948_));
 sky130_fd_sc_hd__o22a_4 _10714_ (.A1(\core_busio.mem_address[27] ),
    .A2(net356),
    .B1(_05946_),
    .B2(_05948_),
    .X(_05949_));
 sky130_fd_sc_hd__mux2_1 _10715_ (.A0(\core_pipeline.memory_to_writeback_alu_data[27] ),
    .A1(_05949_),
    .S(net456),
    .X(_01384_));
 sky130_fd_sc_hd__and2_1 _10716_ (.A(\core_pipeline.pipeline_execute.ex_alu.result_and_clr[28] ),
    .B(net421),
    .X(_05950_));
 sky130_fd_sc_hd__a221o_1 _10717_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_xor[28] ),
    .A2(net422),
    .B1(net352),
    .B2(\core_pipeline.pipeline_execute.ex_alu.result_sll[28] ),
    .C1(net358),
    .X(_05951_));
 sky130_fd_sc_hd__a221o_2 _10718_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_srl_sra[28] ),
    .A2(net354),
    .B1(net418),
    .B2(\core_pipeline.pipeline_execute.ex_alu.result_or[28] ),
    .C1(_05951_),
    .X(_05952_));
 sky130_fd_sc_hd__o22a_4 _10719_ (.A1(\core_busio.mem_address[28] ),
    .A2(net357),
    .B1(_05950_),
    .B2(_05952_),
    .X(_05953_));
 sky130_fd_sc_hd__mux2_1 _10720_ (.A0(\core_pipeline.memory_to_writeback_alu_data[28] ),
    .A1(_05953_),
    .S(net454),
    .X(_01385_));
 sky130_fd_sc_hd__a221o_1 _10721_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_xor[29] ),
    .A2(net423),
    .B1(net355),
    .B2(\core_pipeline.pipeline_execute.ex_alu.result_srl_sra[29] ),
    .C1(net359),
    .X(_05954_));
 sky130_fd_sc_hd__a22o_1 _10722_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_and_clr[29] ),
    .A2(net420),
    .B1(net418),
    .B2(\core_pipeline.pipeline_execute.ex_alu.result_or[29] ),
    .X(_05955_));
 sky130_fd_sc_hd__a21o_1 _10723_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_sll[29] ),
    .A2(net353),
    .B1(_05955_),
    .X(_05956_));
 sky130_fd_sc_hd__o22a_4 _10724_ (.A1(\core_busio.mem_address[29] ),
    .A2(net357),
    .B1(_05954_),
    .B2(_05956_),
    .X(_05957_));
 sky130_fd_sc_hd__mux2_1 _10725_ (.A0(\core_pipeline.memory_to_writeback_alu_data[29] ),
    .A1(_05957_),
    .S(net454),
    .X(_01386_));
 sky130_fd_sc_hd__and2_1 _10726_ (.A(\core_pipeline.pipeline_execute.ex_alu.result_and_clr[30] ),
    .B(net421),
    .X(_05958_));
 sky130_fd_sc_hd__a221o_1 _10727_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_xor[30] ),
    .A2(net423),
    .B1(net353),
    .B2(\core_pipeline.pipeline_execute.ex_alu.result_sll[30] ),
    .C1(net359),
    .X(_05959_));
 sky130_fd_sc_hd__a221o_1 _10728_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_srl_sra[30] ),
    .A2(net355),
    .B1(net419),
    .B2(\core_pipeline.pipeline_execute.ex_alu.result_or[30] ),
    .C1(_05959_),
    .X(_05960_));
 sky130_fd_sc_hd__o22a_2 _10729_ (.A1(\core_busio.mem_address[30] ),
    .A2(net357),
    .B1(_05958_),
    .B2(_05960_),
    .X(_05961_));
 sky130_fd_sc_hd__mux2_1 _10730_ (.A0(\core_pipeline.memory_to_writeback_alu_data[30] ),
    .A1(_05961_),
    .S(net446),
    .X(_01387_));
 sky130_fd_sc_hd__and2_1 _10731_ (.A(\core_pipeline.pipeline_execute.ex_alu.result_and_clr[31] ),
    .B(net421),
    .X(_05962_));
 sky130_fd_sc_hd__a221o_1 _10732_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_xor[31] ),
    .A2(net423),
    .B1(net353),
    .B2(\core_pipeline.pipeline_execute.ex_alu.result_sll[31] ),
    .C1(net359),
    .X(_05963_));
 sky130_fd_sc_hd__a221o_1 _10733_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_srl_sra[31] ),
    .A2(net355),
    .B1(net419),
    .B2(\core_pipeline.pipeline_execute.ex_alu.result_or[31] ),
    .C1(_05963_),
    .X(_05964_));
 sky130_fd_sc_hd__o22a_4 _10734_ (.A1(\core_busio.mem_address[31] ),
    .A2(net357),
    .B1(_05962_),
    .B2(_05964_),
    .X(_05965_));
 sky130_fd_sc_hd__mux2_1 _10735_ (.A0(\core_pipeline.memory_to_writeback_alu_data[31] ),
    .A1(_05965_),
    .S(net454),
    .X(_01388_));
 sky130_fd_sc_hd__mux2_1 _10736_ (.A0(\core_pipeline.decode_to_execute_pc[2] ),
    .A1(\core_pipeline.execute_to_memory_pc[2] ),
    .S(net132),
    .X(_01389_));
 sky130_fd_sc_hd__mux2_1 _10737_ (.A0(\core_pipeline.decode_to_execute_pc[3] ),
    .A1(\core_pipeline.execute_to_memory_pc[3] ),
    .S(net132),
    .X(_01390_));
 sky130_fd_sc_hd__mux2_1 _10738_ (.A0(\core_pipeline.decode_to_execute_pc[4] ),
    .A1(\core_pipeline.execute_to_memory_pc[4] ),
    .S(net123),
    .X(_01391_));
 sky130_fd_sc_hd__mux2_1 _10739_ (.A0(\core_pipeline.decode_to_execute_pc[5] ),
    .A1(\core_pipeline.execute_to_memory_pc[5] ),
    .S(net127),
    .X(_01392_));
 sky130_fd_sc_hd__mux2_1 _10740_ (.A0(\core_pipeline.decode_to_execute_pc[6] ),
    .A1(\core_pipeline.execute_to_memory_pc[6] ),
    .S(net129),
    .X(_01393_));
 sky130_fd_sc_hd__mux2_1 _10741_ (.A0(\core_pipeline.decode_to_execute_pc[7] ),
    .A1(\core_pipeline.execute_to_memory_pc[7] ),
    .S(net137),
    .X(_01394_));
 sky130_fd_sc_hd__mux2_1 _10742_ (.A0(\core_pipeline.decode_to_execute_pc[8] ),
    .A1(\core_pipeline.execute_to_memory_pc[8] ),
    .S(net128),
    .X(_01395_));
 sky130_fd_sc_hd__mux2_1 _10743_ (.A0(\core_pipeline.decode_to_execute_pc[9] ),
    .A1(\core_pipeline.execute_to_memory_pc[9] ),
    .S(net129),
    .X(_01396_));
 sky130_fd_sc_hd__mux2_1 _10744_ (.A0(\core_pipeline.decode_to_execute_pc[10] ),
    .A1(\core_pipeline.execute_to_memory_pc[10] ),
    .S(net129),
    .X(_01397_));
 sky130_fd_sc_hd__mux2_1 _10745_ (.A0(\core_pipeline.decode_to_execute_pc[11] ),
    .A1(\core_pipeline.execute_to_memory_pc[11] ),
    .S(net129),
    .X(_01398_));
 sky130_fd_sc_hd__mux2_1 _10746_ (.A0(\core_pipeline.decode_to_execute_pc[12] ),
    .A1(\core_pipeline.execute_to_memory_pc[12] ),
    .S(net129),
    .X(_01399_));
 sky130_fd_sc_hd__mux2_1 _10747_ (.A0(\core_pipeline.decode_to_execute_pc[13] ),
    .A1(\core_pipeline.execute_to_memory_pc[13] ),
    .S(net129),
    .X(_01400_));
 sky130_fd_sc_hd__mux2_1 _10748_ (.A0(\core_pipeline.decode_to_execute_pc[14] ),
    .A1(\core_pipeline.execute_to_memory_pc[14] ),
    .S(net129),
    .X(_01401_));
 sky130_fd_sc_hd__mux2_1 _10749_ (.A0(\core_pipeline.decode_to_execute_pc[15] ),
    .A1(\core_pipeline.execute_to_memory_pc[15] ),
    .S(net129),
    .X(_01402_));
 sky130_fd_sc_hd__mux2_1 _10750_ (.A0(\core_pipeline.decode_to_execute_pc[16] ),
    .A1(\core_pipeline.execute_to_memory_pc[16] ),
    .S(net128),
    .X(_01403_));
 sky130_fd_sc_hd__mux2_1 _10751_ (.A0(\core_pipeline.decode_to_execute_pc[17] ),
    .A1(\core_pipeline.execute_to_memory_pc[17] ),
    .S(net137),
    .X(_01404_));
 sky130_fd_sc_hd__mux2_1 _10752_ (.A0(\core_pipeline.decode_to_execute_pc[18] ),
    .A1(\core_pipeline.execute_to_memory_pc[18] ),
    .S(net137),
    .X(_01405_));
 sky130_fd_sc_hd__mux2_1 _10753_ (.A0(\core_pipeline.decode_to_execute_pc[19] ),
    .A1(\core_pipeline.execute_to_memory_pc[19] ),
    .S(net137),
    .X(_01406_));
 sky130_fd_sc_hd__mux2_1 _10754_ (.A0(\core_pipeline.decode_to_execute_pc[20] ),
    .A1(\core_pipeline.execute_to_memory_pc[20] ),
    .S(net137),
    .X(_01407_));
 sky130_fd_sc_hd__mux2_1 _10755_ (.A0(\core_pipeline.decode_to_execute_pc[21] ),
    .A1(\core_pipeline.execute_to_memory_pc[21] ),
    .S(net137),
    .X(_01408_));
 sky130_fd_sc_hd__mux2_1 _10756_ (.A0(\core_pipeline.decode_to_execute_pc[22] ),
    .A1(\core_pipeline.execute_to_memory_pc[22] ),
    .S(net137),
    .X(_01409_));
 sky130_fd_sc_hd__mux2_1 _10757_ (.A0(\core_pipeline.decode_to_execute_pc[23] ),
    .A1(\core_pipeline.execute_to_memory_pc[23] ),
    .S(net129),
    .X(_01410_));
 sky130_fd_sc_hd__mux2_1 _10758_ (.A0(\core_pipeline.decode_to_execute_pc[24] ),
    .A1(\core_pipeline.execute_to_memory_pc[24] ),
    .S(net129),
    .X(_01411_));
 sky130_fd_sc_hd__mux2_1 _10759_ (.A0(\core_pipeline.decode_to_execute_pc[25] ),
    .A1(\core_pipeline.execute_to_memory_pc[25] ),
    .S(net129),
    .X(_01412_));
 sky130_fd_sc_hd__mux2_1 _10760_ (.A0(\core_pipeline.decode_to_execute_pc[26] ),
    .A1(\core_pipeline.execute_to_memory_pc[26] ),
    .S(net137),
    .X(_01413_));
 sky130_fd_sc_hd__mux2_1 _10761_ (.A0(\core_pipeline.decode_to_execute_pc[27] ),
    .A1(\core_pipeline.execute_to_memory_pc[27] ),
    .S(net137),
    .X(_01414_));
 sky130_fd_sc_hd__mux2_1 _10762_ (.A0(\core_pipeline.decode_to_execute_pc[28] ),
    .A1(\core_pipeline.execute_to_memory_pc[28] ),
    .S(net137),
    .X(_01415_));
 sky130_fd_sc_hd__mux2_1 _10763_ (.A0(\core_pipeline.decode_to_execute_pc[29] ),
    .A1(\core_pipeline.execute_to_memory_pc[29] ),
    .S(net128),
    .X(_01416_));
 sky130_fd_sc_hd__mux2_1 _10764_ (.A0(\core_pipeline.decode_to_execute_pc[30] ),
    .A1(\core_pipeline.execute_to_memory_pc[30] ),
    .S(net128),
    .X(_01417_));
 sky130_fd_sc_hd__mux2_1 _10765_ (.A0(\core_pipeline.decode_to_execute_pc[31] ),
    .A1(\core_pipeline.execute_to_memory_pc[31] ),
    .S(net137),
    .X(_01418_));
 sky130_fd_sc_hd__mux2_1 _10766_ (.A0(\core_pipeline.decode_to_execute_next_pc[0] ),
    .A1(\core_pipeline.execute_to_memory_next_pc[0] ),
    .S(net126),
    .X(_01419_));
 sky130_fd_sc_hd__mux2_1 _10767_ (.A0(\core_pipeline.decode_to_execute_next_pc[1] ),
    .A1(\core_pipeline.execute_to_memory_next_pc[1] ),
    .S(net132),
    .X(_01420_));
 sky130_fd_sc_hd__mux2_1 _10768_ (.A0(\core_pipeline.execute_to_memory_next_pc[2] ),
    .A1(\core_pipeline.decode_to_execute_next_pc[2] ),
    .S(net157),
    .X(_01421_));
 sky130_fd_sc_hd__mux2_1 _10769_ (.A0(\core_pipeline.execute_to_memory_next_pc[3] ),
    .A1(\core_pipeline.decode_to_execute_next_pc[3] ),
    .S(net157),
    .X(_01422_));
 sky130_fd_sc_hd__mux2_1 _10770_ (.A0(\core_pipeline.execute_to_memory_next_pc[4] ),
    .A1(\core_pipeline.decode_to_execute_next_pc[4] ),
    .S(net149),
    .X(_01423_));
 sky130_fd_sc_hd__mux2_1 _10771_ (.A0(\core_pipeline.execute_to_memory_next_pc[5] ),
    .A1(\core_pipeline.decode_to_execute_next_pc[5] ),
    .S(net157),
    .X(_01424_));
 sky130_fd_sc_hd__mux2_1 _10772_ (.A0(\core_pipeline.execute_to_memory_next_pc[6] ),
    .A1(\core_pipeline.decode_to_execute_next_pc[6] ),
    .S(net151),
    .X(_01425_));
 sky130_fd_sc_hd__mux2_1 _10773_ (.A0(\core_pipeline.execute_to_memory_next_pc[7] ),
    .A1(\core_pipeline.decode_to_execute_next_pc[7] ),
    .S(net158),
    .X(_01426_));
 sky130_fd_sc_hd__mux2_1 _10774_ (.A0(\core_pipeline.execute_to_memory_next_pc[8] ),
    .A1(\core_pipeline.decode_to_execute_next_pc[8] ),
    .S(net151),
    .X(_01427_));
 sky130_fd_sc_hd__mux2_1 _10775_ (.A0(\core_pipeline.execute_to_memory_next_pc[9] ),
    .A1(\core_pipeline.decode_to_execute_next_pc[9] ),
    .S(net154),
    .X(_01428_));
 sky130_fd_sc_hd__mux2_1 _10776_ (.A0(\core_pipeline.execute_to_memory_next_pc[10] ),
    .A1(\core_pipeline.decode_to_execute_next_pc[10] ),
    .S(net154),
    .X(_01429_));
 sky130_fd_sc_hd__mux2_1 _10777_ (.A0(\core_pipeline.execute_to_memory_next_pc[11] ),
    .A1(\core_pipeline.decode_to_execute_next_pc[11] ),
    .S(net154),
    .X(_01430_));
 sky130_fd_sc_hd__mux2_1 _10778_ (.A0(\core_pipeline.execute_to_memory_next_pc[12] ),
    .A1(\core_pipeline.decode_to_execute_next_pc[12] ),
    .S(net153),
    .X(_01431_));
 sky130_fd_sc_hd__mux2_1 _10779_ (.A0(\core_pipeline.execute_to_memory_next_pc[13] ),
    .A1(\core_pipeline.decode_to_execute_next_pc[13] ),
    .S(net154),
    .X(_01432_));
 sky130_fd_sc_hd__mux2_1 _10780_ (.A0(\core_pipeline.execute_to_memory_next_pc[14] ),
    .A1(\core_pipeline.decode_to_execute_next_pc[14] ),
    .S(net153),
    .X(_01433_));
 sky130_fd_sc_hd__mux2_1 _10781_ (.A0(\core_pipeline.execute_to_memory_next_pc[15] ),
    .A1(\core_pipeline.decode_to_execute_next_pc[15] ),
    .S(net153),
    .X(_01434_));
 sky130_fd_sc_hd__mux2_1 _10782_ (.A0(\core_pipeline.execute_to_memory_next_pc[16] ),
    .A1(\core_pipeline.decode_to_execute_next_pc[16] ),
    .S(net153),
    .X(_01435_));
 sky130_fd_sc_hd__mux2_1 _10783_ (.A0(\core_pipeline.execute_to_memory_next_pc[17] ),
    .A1(net652),
    .S(net161),
    .X(_01436_));
 sky130_fd_sc_hd__mux2_1 _10784_ (.A0(\core_pipeline.execute_to_memory_next_pc[18] ),
    .A1(\core_pipeline.decode_to_execute_next_pc[18] ),
    .S(net161),
    .X(_01437_));
 sky130_fd_sc_hd__mux2_1 _10785_ (.A0(\core_pipeline.execute_to_memory_next_pc[19] ),
    .A1(\core_pipeline.decode_to_execute_next_pc[19] ),
    .S(net161),
    .X(_01438_));
 sky130_fd_sc_hd__mux2_1 _10786_ (.A0(\core_pipeline.execute_to_memory_next_pc[20] ),
    .A1(\core_pipeline.decode_to_execute_next_pc[20] ),
    .S(net160),
    .X(_01439_));
 sky130_fd_sc_hd__mux2_1 _10787_ (.A0(\core_pipeline.execute_to_memory_next_pc[21] ),
    .A1(\core_pipeline.decode_to_execute_next_pc[21] ),
    .S(net160),
    .X(_01440_));
 sky130_fd_sc_hd__mux2_1 _10788_ (.A0(\core_pipeline.execute_to_memory_next_pc[22] ),
    .A1(\core_pipeline.decode_to_execute_next_pc[22] ),
    .S(net160),
    .X(_01441_));
 sky130_fd_sc_hd__mux2_1 _10789_ (.A0(\core_pipeline.execute_to_memory_next_pc[23] ),
    .A1(\core_pipeline.decode_to_execute_next_pc[23] ),
    .S(net160),
    .X(_01442_));
 sky130_fd_sc_hd__mux2_1 _10790_ (.A0(\core_pipeline.execute_to_memory_next_pc[24] ),
    .A1(\core_pipeline.decode_to_execute_next_pc[24] ),
    .S(net155),
    .X(_01443_));
 sky130_fd_sc_hd__mux2_1 _10791_ (.A0(\core_pipeline.execute_to_memory_next_pc[25] ),
    .A1(net659),
    .S(net155),
    .X(_01444_));
 sky130_fd_sc_hd__mux2_1 _10792_ (.A0(\core_pipeline.execute_to_memory_next_pc[26] ),
    .A1(\core_pipeline.decode_to_execute_next_pc[26] ),
    .S(net161),
    .X(_01445_));
 sky130_fd_sc_hd__mux2_1 _10793_ (.A0(\core_pipeline.execute_to_memory_next_pc[27] ),
    .A1(\core_pipeline.decode_to_execute_next_pc[27] ),
    .S(net160),
    .X(_01446_));
 sky130_fd_sc_hd__mux2_1 _10794_ (.A0(\core_pipeline.execute_to_memory_next_pc[28] ),
    .A1(\core_pipeline.decode_to_execute_next_pc[28] ),
    .S(net158),
    .X(_01447_));
 sky130_fd_sc_hd__mux2_1 _10795_ (.A0(\core_pipeline.execute_to_memory_next_pc[29] ),
    .A1(\core_pipeline.decode_to_execute_next_pc[29] ),
    .S(net158),
    .X(_01448_));
 sky130_fd_sc_hd__mux2_1 _10796_ (.A0(\core_pipeline.execute_to_memory_next_pc[30] ),
    .A1(\core_pipeline.decode_to_execute_next_pc[30] ),
    .S(net157),
    .X(_01449_));
 sky130_fd_sc_hd__mux2_1 _10797_ (.A0(\core_pipeline.execute_to_memory_next_pc[31] ),
    .A1(\core_pipeline.decode_to_execute_next_pc[31] ),
    .S(net158),
    .X(_01450_));
 sky130_fd_sc_hd__mux2_1 _10798_ (.A0(\core_busio.mem_store_data[0] ),
    .A1(_03877_),
    .S(net140),
    .X(_01451_));
 sky130_fd_sc_hd__mux2_1 _10799_ (.A0(\core_busio.mem_store_data[1] ),
    .A1(_03873_),
    .S(net141),
    .X(_01452_));
 sky130_fd_sc_hd__mux2_1 _10800_ (.A0(\core_busio.mem_store_data[2] ),
    .A1(_03881_),
    .S(net143),
    .X(_01453_));
 sky130_fd_sc_hd__mux2_1 _10801_ (.A0(\core_busio.mem_store_data[3] ),
    .A1(_03886_),
    .S(net139),
    .X(_01454_));
 sky130_fd_sc_hd__mux2_1 _10802_ (.A0(\core_busio.mem_store_data[4] ),
    .A1(_03869_),
    .S(net141),
    .X(_01455_));
 sky130_fd_sc_hd__mux2_1 _10803_ (.A0(\core_busio.mem_store_data[5] ),
    .A1(_03866_),
    .S(net141),
    .X(_01456_));
 sky130_fd_sc_hd__mux2_1 _10804_ (.A0(\core_busio.mem_store_data[6] ),
    .A1(_03859_),
    .S(net143),
    .X(_01457_));
 sky130_fd_sc_hd__mux2_1 _10805_ (.A0(\core_busio.mem_store_data[7] ),
    .A1(_03862_),
    .S(net142),
    .X(_01458_));
 sky130_fd_sc_hd__mux2_1 _10806_ (.A0(\core_busio.mem_store_data[8] ),
    .A1(_03852_),
    .S(net139),
    .X(_01459_));
 sky130_fd_sc_hd__mux2_1 _10807_ (.A0(\core_busio.mem_store_data[9] ),
    .A1(_03847_),
    .S(net139),
    .X(_01460_));
 sky130_fd_sc_hd__mux2_1 _10808_ (.A0(\core_busio.mem_store_data[10] ),
    .A1(_03840_),
    .S(net140),
    .X(_01461_));
 sky130_fd_sc_hd__mux2_1 _10809_ (.A0(\core_busio.mem_store_data[11] ),
    .A1(_03843_),
    .S(net139),
    .X(_01462_));
 sky130_fd_sc_hd__mux2_1 _10810_ (.A0(\core_busio.mem_store_data[12] ),
    .A1(_03836_),
    .S(net139),
    .X(_01463_));
 sky130_fd_sc_hd__mux2_1 _10811_ (.A0(\core_busio.mem_store_data[13] ),
    .A1(_03830_),
    .S(net152),
    .X(_01464_));
 sky130_fd_sc_hd__mux2_1 _10812_ (.A0(\core_busio.mem_store_data[14] ),
    .A1(_03826_),
    .S(net139),
    .X(_01465_));
 sky130_fd_sc_hd__mux2_1 _10813_ (.A0(\core_busio.mem_store_data[15] ),
    .A1(_03822_),
    .S(net152),
    .X(_01466_));
 sky130_fd_sc_hd__mux2_1 _10814_ (.A0(\core_busio.mem_store_data[16] ),
    .A1(_03803_),
    .S(net141),
    .X(_01467_));
 sky130_fd_sc_hd__mux2_1 _10815_ (.A0(\core_busio.mem_store_data[17] ),
    .A1(_03800_),
    .S(net141),
    .X(_01468_));
 sky130_fd_sc_hd__mux2_1 _10816_ (.A0(\core_busio.mem_store_data[18] ),
    .A1(_03793_),
    .S(net142),
    .X(_01469_));
 sky130_fd_sc_hd__mux2_1 _10817_ (.A0(\core_busio.mem_store_data[19] ),
    .A1(_03796_),
    .S(net141),
    .X(_01470_));
 sky130_fd_sc_hd__mux2_1 _10818_ (.A0(\core_busio.mem_store_data[20] ),
    .A1(_03786_),
    .S(net141),
    .X(_01471_));
 sky130_fd_sc_hd__mux2_1 _10819_ (.A0(\core_busio.mem_store_data[21] ),
    .A1(_03789_),
    .S(net156),
    .X(_01472_));
 sky130_fd_sc_hd__mux2_1 _10820_ (.A0(\core_busio.mem_store_data[22] ),
    .A1(_03783_),
    .S(net141),
    .X(_01473_));
 sky130_fd_sc_hd__mux2_1 _10821_ (.A0(\core_busio.mem_store_data[23] ),
    .A1(_03779_),
    .S(net149),
    .X(_01474_));
 sky130_fd_sc_hd__mux2_1 _10822_ (.A0(\core_busio.mem_store_data[24] ),
    .A1(_03766_),
    .S(net141),
    .X(_01475_));
 sky130_fd_sc_hd__mux2_1 _10823_ (.A0(\core_busio.mem_store_data[25] ),
    .A1(_03753_),
    .S(net141),
    .X(_01476_));
 sky130_fd_sc_hd__mux2_1 _10824_ (.A0(\core_busio.mem_store_data[26] ),
    .A1(_03756_),
    .S(net142),
    .X(_01477_));
 sky130_fd_sc_hd__mux2_1 _10825_ (.A0(\core_busio.mem_store_data[27] ),
    .A1(_03760_),
    .S(net141),
    .X(_01478_));
 sky130_fd_sc_hd__mux2_1 _10826_ (.A0(\core_busio.mem_store_data[28] ),
    .A1(_03749_),
    .S(net141),
    .X(_01479_));
 sky130_fd_sc_hd__mux2_1 _10827_ (.A0(\core_busio.mem_store_data[29] ),
    .A1(_03746_),
    .S(net149),
    .X(_01480_));
 sky130_fd_sc_hd__mux2_1 _10828_ (.A0(\core_busio.mem_store_data[30] ),
    .A1(_03771_),
    .S(net141),
    .X(_01481_));
 sky130_fd_sc_hd__mux2_1 _10829_ (.A0(\core_busio.mem_store_data[31] ),
    .A1(_03741_),
    .S(net149),
    .X(_01482_));
 sky130_fd_sc_hd__mux2_1 _10830_ (.A0(\core_pipeline.decode_to_execute_csr_data[0] ),
    .A1(\core_pipeline.execute_to_memory_csr_data[0] ),
    .S(net123),
    .X(_01483_));
 sky130_fd_sc_hd__mux2_1 _10831_ (.A0(\core_pipeline.execute_to_memory_csr_data[1] ),
    .A1(\core_pipeline.decode_to_execute_csr_data[1] ),
    .S(net152),
    .X(_01484_));
 sky130_fd_sc_hd__mux2_1 _10832_ (.A0(\core_pipeline.execute_to_memory_csr_data[2] ),
    .A1(\core_pipeline.decode_to_execute_csr_data[2] ),
    .S(net157),
    .X(_01485_));
 sky130_fd_sc_hd__mux2_1 _10833_ (.A0(\core_pipeline.execute_to_memory_csr_data[3] ),
    .A1(\core_pipeline.decode_to_execute_csr_data[3] ),
    .S(net149),
    .X(_01486_));
 sky130_fd_sc_hd__mux2_1 _10834_ (.A0(\core_pipeline.decode_to_execute_csr_data[4] ),
    .A1(\core_pipeline.execute_to_memory_csr_data[4] ),
    .S(net123),
    .X(_01487_));
 sky130_fd_sc_hd__mux2_1 _10835_ (.A0(\core_pipeline.execute_to_memory_csr_data[5] ),
    .A1(\core_pipeline.decode_to_execute_csr_data[5] ),
    .S(net157),
    .X(_01488_));
 sky130_fd_sc_hd__mux2_1 _10836_ (.A0(\core_pipeline.execute_to_memory_csr_data[6] ),
    .A1(\core_pipeline.decode_to_execute_csr_data[6] ),
    .S(net150),
    .X(_01489_));
 sky130_fd_sc_hd__mux2_1 _10837_ (.A0(\core_pipeline.execute_to_memory_csr_data[7] ),
    .A1(\core_pipeline.decode_to_execute_csr_data[7] ),
    .S(net149),
    .X(_01490_));
 sky130_fd_sc_hd__mux2_1 _10838_ (.A0(\core_pipeline.execute_to_memory_csr_data[8] ),
    .A1(\core_pipeline.decode_to_execute_csr_data[8] ),
    .S(net151),
    .X(_01491_));
 sky130_fd_sc_hd__mux2_1 _10839_ (.A0(\core_pipeline.execute_to_memory_csr_data[9] ),
    .A1(\core_pipeline.decode_to_execute_csr_data[9] ),
    .S(net155),
    .X(_01492_));
 sky130_fd_sc_hd__mux2_1 _10840_ (.A0(\core_pipeline.execute_to_memory_csr_data[10] ),
    .A1(\core_pipeline.decode_to_execute_csr_data[10] ),
    .S(net155),
    .X(_01493_));
 sky130_fd_sc_hd__mux2_1 _10841_ (.A0(\core_pipeline.execute_to_memory_csr_data[11] ),
    .A1(\core_pipeline.decode_to_execute_csr_data[11] ),
    .S(net152),
    .X(_01494_));
 sky130_fd_sc_hd__mux2_1 _10842_ (.A0(\core_pipeline.execute_to_memory_csr_data[12] ),
    .A1(\core_pipeline.decode_to_execute_csr_data[12] ),
    .S(net153),
    .X(_01495_));
 sky130_fd_sc_hd__mux2_1 _10843_ (.A0(\core_pipeline.execute_to_memory_csr_data[13] ),
    .A1(\core_pipeline.decode_to_execute_csr_data[13] ),
    .S(net153),
    .X(_01496_));
 sky130_fd_sc_hd__mux2_1 _10844_ (.A0(\core_pipeline.execute_to_memory_csr_data[14] ),
    .A1(\core_pipeline.decode_to_execute_csr_data[14] ),
    .S(net153),
    .X(_01497_));
 sky130_fd_sc_hd__mux2_1 _10845_ (.A0(\core_pipeline.execute_to_memory_csr_data[15] ),
    .A1(\core_pipeline.decode_to_execute_csr_data[15] ),
    .S(net155),
    .X(_01498_));
 sky130_fd_sc_hd__mux2_1 _10846_ (.A0(\core_pipeline.execute_to_memory_csr_data[16] ),
    .A1(\core_pipeline.decode_to_execute_csr_data[16] ),
    .S(net155),
    .X(_01499_));
 sky130_fd_sc_hd__mux2_1 _10847_ (.A0(\core_pipeline.execute_to_memory_csr_data[17] ),
    .A1(\core_pipeline.decode_to_execute_csr_data[17] ),
    .S(net161),
    .X(_01500_));
 sky130_fd_sc_hd__mux2_1 _10848_ (.A0(\core_pipeline.execute_to_memory_csr_data[18] ),
    .A1(\core_pipeline.decode_to_execute_csr_data[18] ),
    .S(net160),
    .X(_01501_));
 sky130_fd_sc_hd__mux2_1 _10849_ (.A0(\core_pipeline.execute_to_memory_csr_data[19] ),
    .A1(\core_pipeline.decode_to_execute_csr_data[19] ),
    .S(net160),
    .X(_01502_));
 sky130_fd_sc_hd__mux2_1 _10850_ (.A0(\core_pipeline.execute_to_memory_csr_data[20] ),
    .A1(\core_pipeline.decode_to_execute_csr_data[20] ),
    .S(net160),
    .X(_01503_));
 sky130_fd_sc_hd__mux2_1 _10851_ (.A0(\core_pipeline.execute_to_memory_csr_data[21] ),
    .A1(\core_pipeline.decode_to_execute_csr_data[21] ),
    .S(net158),
    .X(_01504_));
 sky130_fd_sc_hd__mux2_1 _10852_ (.A0(\core_pipeline.execute_to_memory_csr_data[22] ),
    .A1(\core_pipeline.decode_to_execute_csr_data[22] ),
    .S(net160),
    .X(_01505_));
 sky130_fd_sc_hd__mux2_1 _10853_ (.A0(\core_pipeline.execute_to_memory_csr_data[23] ),
    .A1(\core_pipeline.decode_to_execute_csr_data[23] ),
    .S(net155),
    .X(_01506_));
 sky130_fd_sc_hd__mux2_1 _10854_ (.A0(\core_pipeline.execute_to_memory_csr_data[24] ),
    .A1(\core_pipeline.decode_to_execute_csr_data[24] ),
    .S(net155),
    .X(_01507_));
 sky130_fd_sc_hd__mux2_1 _10855_ (.A0(\core_pipeline.execute_to_memory_csr_data[25] ),
    .A1(\core_pipeline.decode_to_execute_csr_data[25] ),
    .S(net155),
    .X(_01508_));
 sky130_fd_sc_hd__mux2_1 _10856_ (.A0(\core_pipeline.execute_to_memory_csr_data[26] ),
    .A1(\core_pipeline.decode_to_execute_csr_data[26] ),
    .S(net150),
    .X(_01509_));
 sky130_fd_sc_hd__mux2_1 _10857_ (.A0(\core_pipeline.execute_to_memory_csr_data[27] ),
    .A1(\core_pipeline.decode_to_execute_csr_data[27] ),
    .S(net158),
    .X(_01510_));
 sky130_fd_sc_hd__mux2_1 _10858_ (.A0(\core_pipeline.execute_to_memory_csr_data[28] ),
    .A1(\core_pipeline.decode_to_execute_csr_data[28] ),
    .S(net158),
    .X(_01511_));
 sky130_fd_sc_hd__mux2_1 _10859_ (.A0(\core_pipeline.execute_to_memory_csr_data[29] ),
    .A1(\core_pipeline.decode_to_execute_csr_data[29] ),
    .S(net158),
    .X(_01512_));
 sky130_fd_sc_hd__mux2_1 _10860_ (.A0(\core_pipeline.execute_to_memory_csr_data[30] ),
    .A1(\core_pipeline.decode_to_execute_csr_data[30] ),
    .S(net156),
    .X(_01513_));
 sky130_fd_sc_hd__mux2_1 _10861_ (.A0(\core_pipeline.execute_to_memory_csr_data[31] ),
    .A1(\core_pipeline.decode_to_execute_csr_data[31] ),
    .S(net157),
    .X(_01514_));
 sky130_fd_sc_hd__mux2_1 _10862_ (.A0(\core_pipeline.execute_to_memory_jump ),
    .A1(\core_pipeline.decode_to_execute_jump ),
    .S(net143),
    .X(_01515_));
 sky130_fd_sc_hd__mux2_1 _10863_ (.A0(\core_pipeline.execute_to_memory_branch ),
    .A1(net651),
    .S(net143),
    .X(_01516_));
 sky130_fd_sc_hd__mux2_1 _10864_ (.A0(\core_pipeline.decode_to_execute_csr_write ),
    .A1(\core_pipeline.execute_to_memory_csr_write ),
    .S(net132),
    .X(_01517_));
 sky130_fd_sc_hd__mux2_1 _10865_ (.A0(\core_pipeline.execute_to_memory_load ),
    .A1(\core_pipeline.decode_to_execute_load ),
    .S(net147),
    .X(_01518_));
 sky130_fd_sc_hd__mux2_1 _10866_ (.A0(\core_pipeline.execute_to_memory_store ),
    .A1(\core_pipeline.decode_to_execute_store ),
    .S(net142),
    .X(_01519_));
 sky130_fd_sc_hd__mux2_1 _10867_ (.A0(\core_busio.mem_size[0] ),
    .A1(\core_pipeline.decode_to_execute_cmp_function[0] ),
    .S(net142),
    .X(_01520_));
 sky130_fd_sc_hd__mux2_1 _10868_ (.A0(\core_busio.mem_size[1] ),
    .A1(\core_pipeline.decode_to_execute_cmp_function[1] ),
    .S(net141),
    .X(_01521_));
 sky130_fd_sc_hd__mux2_1 _10869_ (.A0(\core_busio.mem_signed ),
    .A1(net653),
    .S(net149),
    .X(_01522_));
 sky130_fd_sc_hd__mux2_1 _10870_ (.A0(\core_pipeline.execute_to_memory_bypass_memory ),
    .A1(\core_pipeline.decode_to_execute_bypass_memory ),
    .S(net147),
    .X(_01523_));
 sky130_fd_sc_hd__mux2_1 _10871_ (.A0(net499),
    .A1(\core_pipeline.decode_to_execute_write_select[0] ),
    .S(net143),
    .X(_01524_));
 sky130_fd_sc_hd__mux2_1 _10872_ (.A0(\core_pipeline.decode_to_execute_write_select[1] ),
    .A1(\core_pipeline.execute_to_memory_write_select[1] ),
    .S(net127),
    .X(_01525_));
 sky130_fd_sc_hd__mux2_1 _10873_ (.A0(\core_pipeline.decode_to_execute_rd_address[0] ),
    .A1(\core_pipeline.execute_to_memory_rd_address[0] ),
    .S(net130),
    .X(_01526_));
 sky130_fd_sc_hd__mux2_1 _10874_ (.A0(\core_pipeline.decode_to_execute_rd_address[1] ),
    .A1(\core_pipeline.execute_to_memory_rd_address[1] ),
    .S(net132),
    .X(_01527_));
 sky130_fd_sc_hd__mux2_1 _10875_ (.A0(\core_pipeline.decode_to_execute_rd_address[2] ),
    .A1(\core_pipeline.execute_to_memory_rd_address[2] ),
    .S(net132),
    .X(_01528_));
 sky130_fd_sc_hd__mux2_1 _10876_ (.A0(\core_pipeline.decode_to_execute_rd_address[3] ),
    .A1(\core_pipeline.execute_to_memory_rd_address[3] ),
    .S(net130),
    .X(_01529_));
 sky130_fd_sc_hd__mux2_1 _10877_ (.A0(\core_pipeline.decode_to_execute_rd_address[4] ),
    .A1(\core_pipeline.execute_to_memory_rd_address[4] ),
    .S(net130),
    .X(_01530_));
 sky130_fd_sc_hd__mux2_1 _10878_ (.A0(\core_pipeline.execute_to_memory_csr_address[0] ),
    .A1(\core_pipeline.decode_to_execute_csr_address[0] ),
    .S(net146),
    .X(_01531_));
 sky130_fd_sc_hd__mux2_1 _10879_ (.A0(\core_pipeline.execute_to_memory_csr_address[1] ),
    .A1(\core_pipeline.decode_to_execute_csr_address[1] ),
    .S(net146),
    .X(_01532_));
 sky130_fd_sc_hd__mux2_1 _10880_ (.A0(\core_pipeline.execute_to_memory_csr_address[2] ),
    .A1(\core_pipeline.decode_to_execute_csr_address[2] ),
    .S(net146),
    .X(_01533_));
 sky130_fd_sc_hd__mux2_1 _10881_ (.A0(\core_pipeline.execute_to_memory_csr_address[3] ),
    .A1(\core_pipeline.decode_to_execute_csr_address[3] ),
    .S(net146),
    .X(_01534_));
 sky130_fd_sc_hd__mux2_1 _10882_ (.A0(\core_pipeline.execute_to_memory_csr_address[4] ),
    .A1(\core_pipeline.decode_to_execute_csr_address[4] ),
    .S(net146),
    .X(_01535_));
 sky130_fd_sc_hd__mux2_1 _10883_ (.A0(\core_pipeline.execute_to_memory_csr_address[5] ),
    .A1(\core_pipeline.decode_to_execute_csr_address[5] ),
    .S(net146),
    .X(_01536_));
 sky130_fd_sc_hd__mux2_1 _10884_ (.A0(\core_pipeline.execute_to_memory_csr_address[6] ),
    .A1(\core_pipeline.decode_to_execute_csr_address[6] ),
    .S(net146),
    .X(_01537_));
 sky130_fd_sc_hd__mux2_1 _10885_ (.A0(\core_pipeline.execute_to_memory_csr_address[7] ),
    .A1(\core_pipeline.decode_to_execute_csr_address[7] ),
    .S(net146),
    .X(_01538_));
 sky130_fd_sc_hd__mux2_1 _10886_ (.A0(\core_pipeline.execute_to_memory_csr_address[8] ),
    .A1(\core_pipeline.decode_to_execute_csr_address[8] ),
    .S(net148),
    .X(_01539_));
 sky130_fd_sc_hd__mux2_1 _10887_ (.A0(\core_pipeline.execute_to_memory_csr_address[9] ),
    .A1(\core_pipeline.decode_to_execute_csr_address[9] ),
    .S(net146),
    .X(_01540_));
 sky130_fd_sc_hd__mux2_1 _10888_ (.A0(\core_pipeline.execute_to_memory_csr_address[10] ),
    .A1(\core_pipeline.decode_to_execute_csr_address[10] ),
    .S(net148),
    .X(_01541_));
 sky130_fd_sc_hd__mux2_1 _10889_ (.A0(\core_pipeline.execute_to_memory_csr_address[11] ),
    .A1(\core_pipeline.decode_to_execute_csr_address[11] ),
    .S(net146),
    .X(_01542_));
 sky130_fd_sc_hd__mux2_1 _10890_ (.A0(\core_pipeline.execute_to_memory_mret ),
    .A1(\core_pipeline.decode_to_execute_mret ),
    .S(net147),
    .X(_01543_));
 sky130_fd_sc_hd__o22a_1 _10891_ (.A1(\core_pipeline.decode_to_execute_csr_readable ),
    .A2(_03412_),
    .B1(\core_pipeline.decode_to_execute_csr_writeable ),
    .B2(_03337_),
    .X(_05966_));
 sky130_fd_sc_hd__or3b_1 _10892_ (.A(\core_pipeline.decode_to_execute_exception ),
    .B(net133),
    .C_N(_05966_),
    .X(_05967_));
 sky130_fd_sc_hd__o21a_1 _10893_ (.A1(\core_pipeline.execute_to_memory_exception ),
    .A2(net147),
    .B1(_05967_),
    .X(_01544_));
 sky130_fd_sc_hd__and3b_4 _10894_ (.A_N(\core_pipeline.decode_to_execute_alu_function[0] ),
    .B(\core_pipeline.decode_to_execute_alu_function[1] ),
    .C(\core_pipeline.decode_to_execute_alu_function[2] ),
    .X(_05968_));
 sky130_fd_sc_hd__or2_1 _10895_ (.A(net374),
    .B(_04495_),
    .X(_05969_));
 sky130_fd_sc_hd__mux2_1 _10896_ (.A0(\core_pipeline.pipeline_execute.ex_alu.result_or[0] ),
    .A1(_05969_),
    .S(net414),
    .X(_01545_));
 sky130_fd_sc_hd__mux2_1 _10897_ (.A0(\core_pipeline.pipeline_execute.ex_alu.result_or[1] ),
    .A1(_05817_),
    .S(net414),
    .X(_01546_));
 sky130_fd_sc_hd__nand2_1 _10898_ (.A(_04511_),
    .B(net414),
    .Y(_05970_));
 sky130_fd_sc_hd__o22a_1 _10899_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_or[2] ),
    .A2(net414),
    .B1(_05970_),
    .B2(net384),
    .X(_01547_));
 sky130_fd_sc_hd__nand2_1 _10900_ (.A(_04517_),
    .B(net414),
    .Y(_05971_));
 sky130_fd_sc_hd__o22a_1 _10901_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_or[3] ),
    .A2(net414),
    .B1(_05971_),
    .B2(net395),
    .X(_01548_));
 sky130_fd_sc_hd__nand2_1 _10902_ (.A(net393),
    .B(net414),
    .Y(_05972_));
 sky130_fd_sc_hd__o22a_1 _10903_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_or[4] ),
    .A2(net414),
    .B1(_05972_),
    .B2(_04522_),
    .X(_01549_));
 sky130_fd_sc_hd__nand2_1 _10904_ (.A(_05666_),
    .B(net414),
    .Y(_05973_));
 sky130_fd_sc_hd__o22a_1 _10905_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_or[5] ),
    .A2(net414),
    .B1(_05973_),
    .B2(_04530_),
    .X(_01550_));
 sky130_fd_sc_hd__nand2_1 _10906_ (.A(_05662_),
    .B(net414),
    .Y(_05974_));
 sky130_fd_sc_hd__o22a_1 _10907_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_or[6] ),
    .A2(net414),
    .B1(_05974_),
    .B2(_04538_),
    .X(_01551_));
 sky130_fd_sc_hd__nand2_1 _10908_ (.A(_04545_),
    .B(_05657_),
    .Y(_05975_));
 sky130_fd_sc_hd__mux2_1 _10909_ (.A0(\core_pipeline.pipeline_execute.ex_alu.result_or[7] ),
    .A1(_05975_),
    .S(net414),
    .X(_01552_));
 sky130_fd_sc_hd__nand2_1 _10910_ (.A(_05633_),
    .B(net415),
    .Y(_05976_));
 sky130_fd_sc_hd__o22a_1 _10911_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_or[8] ),
    .A2(net415),
    .B1(_05976_),
    .B2(_04554_),
    .X(_01553_));
 sky130_fd_sc_hd__nand2_1 _10912_ (.A(_05636_),
    .B(net415),
    .Y(_05977_));
 sky130_fd_sc_hd__o22a_1 _10913_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_or[9] ),
    .A2(net415),
    .B1(_05977_),
    .B2(_04566_),
    .X(_01554_));
 sky130_fd_sc_hd__nand2_1 _10914_ (.A(_05651_),
    .B(net415),
    .Y(_05978_));
 sky130_fd_sc_hd__o22a_1 _10915_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_or[10] ),
    .A2(net415),
    .B1(_05978_),
    .B2(_04574_),
    .X(_01555_));
 sky130_fd_sc_hd__nand2_1 _10916_ (.A(_05639_),
    .B(net415),
    .Y(_05979_));
 sky130_fd_sc_hd__o22a_1 _10917_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_or[11] ),
    .A2(net415),
    .B1(_05979_),
    .B2(_04582_),
    .X(_01556_));
 sky130_fd_sc_hd__nand2_1 _10918_ (.A(net371),
    .B(net415),
    .Y(_05980_));
 sky130_fd_sc_hd__o22a_1 _10919_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_or[12] ),
    .A2(net415),
    .B1(_05980_),
    .B2(_05642_),
    .X(_01557_));
 sky130_fd_sc_hd__nand2_1 _10920_ (.A(_04599_),
    .B(net415),
    .Y(_05981_));
 sky130_fd_sc_hd__o22a_1 _10921_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_or[13] ),
    .A2(net416),
    .B1(_05981_),
    .B2(_05623_),
    .X(_01558_));
 sky130_fd_sc_hd__mux2_1 _10922_ (.A0(\core_pipeline.pipeline_execute.ex_alu.result_or[14] ),
    .A1(_05619_),
    .S(net415),
    .X(_01559_));
 sky130_fd_sc_hd__nand2_1 _10923_ (.A(_05626_),
    .B(net416),
    .Y(_05982_));
 sky130_fd_sc_hd__o22a_1 _10924_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_or[15] ),
    .A2(net416),
    .B1(_05982_),
    .B2(_04618_),
    .X(_01560_));
 sky130_fd_sc_hd__and2b_1 _10925_ (.A_N(_05760_),
    .B(net416),
    .X(_05983_));
 sky130_fd_sc_hd__o2bb2a_1 _10926_ (.A1_N(_05758_),
    .A2_N(_05983_),
    .B1(net416),
    .B2(\core_pipeline.pipeline_execute.ex_alu.result_or[16] ),
    .X(_01561_));
 sky130_fd_sc_hd__nand2_1 _10927_ (.A(_05745_),
    .B(net416),
    .Y(_05984_));
 sky130_fd_sc_hd__o22a_1 _10928_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_or[17] ),
    .A2(net416),
    .B1(_05984_),
    .B2(_05748_),
    .X(_01562_));
 sky130_fd_sc_hd__nand2_1 _10929_ (.A(_05779_),
    .B(net416),
    .Y(_05985_));
 sky130_fd_sc_hd__o22a_1 _10930_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_or[18] ),
    .A2(net416),
    .B1(_05985_),
    .B2(_05781_),
    .X(_01563_));
 sky130_fd_sc_hd__nand2_1 _10931_ (.A(_05786_),
    .B(_05788_),
    .Y(_05986_));
 sky130_fd_sc_hd__mux2_1 _10932_ (.A0(\core_pipeline.pipeline_execute.ex_alu.result_or[19] ),
    .A1(_05986_),
    .S(net415),
    .X(_01564_));
 sky130_fd_sc_hd__mux2_1 _10933_ (.A0(\core_pipeline.pipeline_execute.ex_alu.result_or[20] ),
    .A1(_05776_),
    .S(net417),
    .X(_01565_));
 sky130_fd_sc_hd__nand2_1 _10934_ (.A(_05763_),
    .B(net417),
    .Y(_05987_));
 sky130_fd_sc_hd__o22a_1 _10935_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_or[21] ),
    .A2(net417),
    .B1(_05987_),
    .B2(_05765_),
    .X(_01566_));
 sky130_fd_sc_hd__mux2_1 _10936_ (.A0(\core_pipeline.pipeline_execute.ex_alu.result_or[22] ),
    .A1(_05754_),
    .S(net417),
    .X(_01567_));
 sky130_fd_sc_hd__nand2_1 _10937_ (.A(_05738_),
    .B(net414),
    .Y(_05988_));
 sky130_fd_sc_hd__o22a_1 _10938_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_or[23] ),
    .A2(net414),
    .B1(_05988_),
    .B2(_05740_),
    .X(_01568_));
 sky130_fd_sc_hd__mux2_1 _10939_ (.A0(\core_pipeline.pipeline_execute.ex_alu.result_or[24] ),
    .A1(_05718_),
    .S(net415),
    .X(_01569_));
 sky130_fd_sc_hd__or2_1 _10940_ (.A(_05729_),
    .B(_05731_),
    .X(_05989_));
 sky130_fd_sc_hd__mux2_1 _10941_ (.A0(\core_pipeline.pipeline_execute.ex_alu.result_or[25] ),
    .A1(_05989_),
    .S(net415),
    .X(_01570_));
 sky130_fd_sc_hd__nand2_1 _10942_ (.A(_05710_),
    .B(net417),
    .Y(_05990_));
 sky130_fd_sc_hd__o22a_1 _10943_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_or[26] ),
    .A2(net417),
    .B1(_05990_),
    .B2(_05712_),
    .X(_01571_));
 sky130_fd_sc_hd__nand2_1 _10944_ (.A(net360),
    .B(net415),
    .Y(_05991_));
 sky130_fd_sc_hd__o22a_1 _10945_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_or[27] ),
    .A2(net415),
    .B1(_05991_),
    .B2(_05722_),
    .X(_01572_));
 sky130_fd_sc_hd__nand2_1 _10946_ (.A(_05697_),
    .B(net417),
    .Y(_05992_));
 sky130_fd_sc_hd__o22a_1 _10947_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_or[28] ),
    .A2(net417),
    .B1(_05992_),
    .B2(_05699_),
    .X(_01573_));
 sky130_fd_sc_hd__nand2_1 _10948_ (.A(_05704_),
    .B(net417),
    .Y(_05993_));
 sky130_fd_sc_hd__o22a_1 _10949_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_or[29] ),
    .A2(net417),
    .B1(_05993_),
    .B2(_05702_),
    .X(_01574_));
 sky130_fd_sc_hd__mux2_1 _10950_ (.A0(\core_pipeline.pipeline_execute.ex_alu.result_or[30] ),
    .A1(_05692_),
    .S(net414),
    .X(_01575_));
 sky130_fd_sc_hd__nand2_1 _10951_ (.A(_05612_),
    .B(net414),
    .Y(_05994_));
 sky130_fd_sc_hd__o22a_1 _10952_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_or[31] ),
    .A2(_05968_),
    .B1(_05994_),
    .B2(_05614_),
    .X(_01576_));
 sky130_fd_sc_hd__and2_1 _10953_ (.A(net376),
    .B(_05712_),
    .X(_05995_));
 sky130_fd_sc_hd__o21bai_1 _10954_ (.A1(net376),
    .A2(net360),
    .B1_N(_05995_),
    .Y(_05996_));
 sky130_fd_sc_hd__nor2_1 _10955_ (.A(net382),
    .B(_05996_),
    .Y(_05997_));
 sky130_fd_sc_hd__and2_1 _10956_ (.A(net373),
    .B(_05731_),
    .X(_05998_));
 sky130_fd_sc_hd__and2_1 _10957_ (.A(net376),
    .B(_05717_),
    .X(_05999_));
 sky130_fd_sc_hd__nor2_1 _10958_ (.A(_05998_),
    .B(_05999_),
    .Y(_06000_));
 sky130_fd_sc_hd__a21oi_1 _10959_ (.A1(net382),
    .A2(_06000_),
    .B1(_05997_),
    .Y(_06001_));
 sky130_fd_sc_hd__mux2_1 _10960_ (.A0(_05614_),
    .A1(_05687_),
    .S(net376),
    .X(_06002_));
 sky130_fd_sc_hd__or2_2 _10961_ (.A(net376),
    .B(_05704_),
    .X(_06003_));
 sky130_fd_sc_hd__nand2_1 _10962_ (.A(net376),
    .B(_05699_),
    .Y(_06004_));
 sky130_fd_sc_hd__nand2_1 _10963_ (.A(_06003_),
    .B(_06004_),
    .Y(_06005_));
 sky130_fd_sc_hd__mux2_1 _10964_ (.A0(_06002_),
    .A1(_06005_),
    .S(net382),
    .X(_06006_));
 sky130_fd_sc_hd__mux2_1 _10965_ (.A0(_06001_),
    .A1(_06006_),
    .S(net385),
    .X(_06007_));
 sky130_fd_sc_hd__nor2_1 _10966_ (.A(net375),
    .B(_05788_),
    .Y(_06008_));
 sky130_fd_sc_hd__and2_1 _10967_ (.A(net375),
    .B(_05781_),
    .X(_06009_));
 sky130_fd_sc_hd__nor2_1 _10968_ (.A(_06008_),
    .B(_06009_),
    .Y(_06010_));
 sky130_fd_sc_hd__and2_1 _10969_ (.A(net372),
    .B(_05748_),
    .X(_06011_));
 sky130_fd_sc_hd__and2_1 _10970_ (.A(net375),
    .B(_05760_),
    .X(_06012_));
 sky130_fd_sc_hd__nor2_1 _10971_ (.A(_06011_),
    .B(_06012_),
    .Y(_06013_));
 sky130_fd_sc_hd__or2_1 _10972_ (.A(net382),
    .B(_06010_),
    .X(_06014_));
 sky130_fd_sc_hd__o21ai_1 _10973_ (.A1(net378),
    .A2(_06013_),
    .B1(_06014_),
    .Y(_06015_));
 sky130_fd_sc_hd__nand2_1 _10974_ (.A(net375),
    .B(_05753_),
    .Y(_06016_));
 sky130_fd_sc_hd__a21boi_1 _10975_ (.A1(net373),
    .A2(_05740_),
    .B1_N(_06016_),
    .Y(_06017_));
 sky130_fd_sc_hd__nand2_1 _10976_ (.A(net372),
    .B(_05765_),
    .Y(_06018_));
 sky130_fd_sc_hd__nor2_1 _10977_ (.A(net372),
    .B(_05773_),
    .Y(_06019_));
 sky130_fd_sc_hd__o21a_1 _10978_ (.A1(net372),
    .A2(_05773_),
    .B1(_06018_),
    .X(_06020_));
 sky130_fd_sc_hd__or2_1 _10979_ (.A(net382),
    .B(_06017_),
    .X(_06021_));
 sky130_fd_sc_hd__o21ai_1 _10980_ (.A1(net379),
    .A2(_06020_),
    .B1(_06021_),
    .Y(_06022_));
 sky130_fd_sc_hd__mux2_1 _10981_ (.A0(_06015_),
    .A1(_06022_),
    .S(net385),
    .X(_06023_));
 sky130_fd_sc_hd__mux2_2 _10982_ (.A0(_06007_),
    .A1(_06023_),
    .S(net398),
    .X(_06024_));
 sky130_fd_sc_hd__and3b_4 _10983_ (.A_N(\core_pipeline.decode_to_execute_alu_function[1] ),
    .B(\core_pipeline.decode_to_execute_alu_function[0] ),
    .C(\core_pipeline.decode_to_execute_alu_function[2] ),
    .X(_06025_));
 sky130_fd_sc_hd__nand3b_4 _10984_ (.A_N(\core_pipeline.decode_to_execute_alu_function[1] ),
    .B(\core_pipeline.decode_to_execute_alu_function[0] ),
    .C(\core_pipeline.decode_to_execute_alu_function[2] ),
    .Y(_06026_));
 sky130_fd_sc_hd__a21oi_1 _10985_ (.A1(net375),
    .A2(_04574_),
    .B1(_04588_),
    .Y(_06027_));
 sky130_fd_sc_hd__nor2_1 _10986_ (.A(_04555_),
    .B(_04572_),
    .Y(_06028_));
 sky130_fd_sc_hd__or2_1 _10987_ (.A(net378),
    .B(_06028_),
    .X(_06029_));
 sky130_fd_sc_hd__o21ai_1 _10988_ (.A1(net381),
    .A2(_06027_),
    .B1(_06029_),
    .Y(_06030_));
 sky130_fd_sc_hd__and2_1 _10989_ (.A(net372),
    .B(_04618_),
    .X(_06031_));
 sky130_fd_sc_hd__nor2_1 _10990_ (.A(_04609_),
    .B(_06031_),
    .Y(_06032_));
 sky130_fd_sc_hd__nor2_1 _10991_ (.A(_04591_),
    .B(_04606_),
    .Y(_06033_));
 sky130_fd_sc_hd__or2_1 _10992_ (.A(net381),
    .B(_06032_),
    .X(_06034_));
 sky130_fd_sc_hd__o21ai_1 _10993_ (.A1(net378),
    .A2(_06033_),
    .B1(_06034_),
    .Y(_06035_));
 sky130_fd_sc_hd__mux2_2 _10994_ (.A0(_06030_),
    .A1(_06035_),
    .S(net385),
    .X(_06036_));
 sky130_fd_sc_hd__mux2_1 _10995_ (.A0(_04511_),
    .A1(_04517_),
    .S(net374),
    .X(_06037_));
 sky130_fd_sc_hd__nor2_1 _10996_ (.A(net380),
    .B(_06037_),
    .Y(_06038_));
 sky130_fd_sc_hd__a311o_1 _10997_ (.A1(net380),
    .A2(net374),
    .A3(_04502_),
    .B1(_04497_),
    .C1(net384),
    .X(_06039_));
 sky130_fd_sc_hd__a21oi_1 _10998_ (.A1(net377),
    .A2(_04538_),
    .B1(_04556_),
    .Y(_06040_));
 sky130_fd_sc_hd__nor2_1 _10999_ (.A(_04524_),
    .B(_04536_),
    .Y(_06041_));
 sky130_fd_sc_hd__mux2_1 _11000_ (.A0(_06040_),
    .A1(_06041_),
    .S(net380),
    .X(_06042_));
 sky130_fd_sc_hd__o2bb2a_1 _11001_ (.A1_N(net384),
    .A2_N(_06042_),
    .B1(_06039_),
    .B2(_06038_),
    .X(_06043_));
 sky130_fd_sc_hd__mux2_1 _11002_ (.A0(_06036_),
    .A1(_06043_),
    .S(net399),
    .X(_06044_));
 sky130_fd_sc_hd__mux2_1 _11003_ (.A0(_06024_),
    .A1(_06044_),
    .S(net393),
    .X(_06045_));
 sky130_fd_sc_hd__mux2_1 _11004_ (.A0(\core_pipeline.pipeline_execute.ex_alu.result_srl_sra[0] ),
    .A1(_06045_),
    .S(net412),
    .X(_01577_));
 sky130_fd_sc_hd__nand2_1 _11005_ (.A(net373),
    .B(_05699_),
    .Y(_06046_));
 sky130_fd_sc_hd__or2_1 _11006_ (.A(net373),
    .B(net360),
    .X(_06047_));
 sky130_fd_sc_hd__and3_1 _11007_ (.A(_04488_),
    .B(_06046_),
    .C(_06047_),
    .X(_06048_));
 sky130_fd_sc_hd__nand2_1 _11008_ (.A(net376),
    .B(_05731_),
    .Y(_06049_));
 sky130_fd_sc_hd__nand2_1 _11009_ (.A(net373),
    .B(_05712_),
    .Y(_06050_));
 sky130_fd_sc_hd__a31oi_2 _11010_ (.A1(net382),
    .A2(_06049_),
    .A3(_06050_),
    .B1(_06048_),
    .Y(_06051_));
 sky130_fd_sc_hd__nor2_1 _11011_ (.A(net631),
    .B(net377),
    .Y(_06052_));
 sky130_fd_sc_hd__a21o_1 _11012_ (.A1(net459),
    .A2(net373),
    .B1(net383),
    .X(_06053_));
 sky130_fd_sc_hd__or2_1 _11013_ (.A(net373),
    .B(_05704_),
    .X(_06054_));
 sky130_fd_sc_hd__o21ai_1 _11014_ (.A1(net376),
    .A2(_05688_),
    .B1(_06054_),
    .Y(_06055_));
 sky130_fd_sc_hd__a2bb2o_1 _11015_ (.A1_N(_05615_),
    .A2_N(_06053_),
    .B1(_06055_),
    .B2(net383),
    .X(_06056_));
 sky130_fd_sc_hd__mux2_1 _11016_ (.A0(_06051_),
    .A1(_06056_),
    .S(net384),
    .X(_06057_));
 sky130_fd_sc_hd__mux2_1 _11017_ (.A0(_05773_),
    .A1(_05788_),
    .S(net375),
    .X(_06058_));
 sky130_fd_sc_hd__and2_1 _11018_ (.A(net372),
    .B(_05781_),
    .X(_06059_));
 sky130_fd_sc_hd__and2_1 _11019_ (.A(net375),
    .B(_05748_),
    .X(_06060_));
 sky130_fd_sc_hd__nor2_1 _11020_ (.A(_06059_),
    .B(_06060_),
    .Y(_06061_));
 sky130_fd_sc_hd__mux2_1 _11021_ (.A0(_06058_),
    .A1(_06061_),
    .S(net381),
    .X(_06062_));
 sky130_fd_sc_hd__nand2_1 _11022_ (.A(net372),
    .B(_05717_),
    .Y(_06063_));
 sky130_fd_sc_hd__nand2_1 _11023_ (.A(net376),
    .B(_05740_),
    .Y(_06064_));
 sky130_fd_sc_hd__and2_1 _11024_ (.A(_06063_),
    .B(_06064_),
    .X(_06065_));
 sky130_fd_sc_hd__nand2_1 _11025_ (.A(net375),
    .B(_05765_),
    .Y(_06066_));
 sky130_fd_sc_hd__nand2_1 _11026_ (.A(net372),
    .B(_05753_),
    .Y(_06067_));
 sky130_fd_sc_hd__and2_1 _11027_ (.A(_06066_),
    .B(_06067_),
    .X(_06068_));
 sky130_fd_sc_hd__mux2_1 _11028_ (.A0(_06065_),
    .A1(_06068_),
    .S(net382),
    .X(_06069_));
 sky130_fd_sc_hd__inv_2 _11029_ (.A(_06069_),
    .Y(_06070_));
 sky130_fd_sc_hd__mux2_1 _11030_ (.A0(_06062_),
    .A1(_06069_),
    .S(net384),
    .X(_06071_));
 sky130_fd_sc_hd__inv_2 _11031_ (.A(_06071_),
    .Y(_06072_));
 sky130_fd_sc_hd__mux2_1 _11032_ (.A0(_06057_),
    .A1(_06072_),
    .S(net398),
    .X(_06073_));
 sky130_fd_sc_hd__nor2_1 _11033_ (.A(_04567_),
    .B(_04579_),
    .Y(_06074_));
 sky130_fd_sc_hd__nor2_1 _11034_ (.A(_04583_),
    .B(_04597_),
    .Y(_06075_));
 sky130_fd_sc_hd__mux2_1 _11035_ (.A0(_06074_),
    .A1(_06075_),
    .S(net378),
    .X(_06076_));
 sky130_fd_sc_hd__nor2_1 _11036_ (.A(_04600_),
    .B(_04616_),
    .Y(_06077_));
 sky130_fd_sc_hd__and2_1 _11037_ (.A(net372),
    .B(_05760_),
    .X(_06078_));
 sky130_fd_sc_hd__a21oi_1 _11038_ (.A1(net375),
    .A2(_04618_),
    .B1(_06078_),
    .Y(_06079_));
 sky130_fd_sc_hd__mux2_1 _11039_ (.A0(_06077_),
    .A1(_06079_),
    .S(net378),
    .X(_06080_));
 sky130_fd_sc_hd__mux2_1 _11040_ (.A0(_06076_),
    .A1(_06080_),
    .S(net384),
    .X(_06081_));
 sky130_fd_sc_hd__nor2_1 _11041_ (.A(_04518_),
    .B(_04528_),
    .Y(_06082_));
 sky130_fd_sc_hd__a211oi_1 _11042_ (.A1(net377),
    .A2(_04502_),
    .B1(_04515_),
    .C1(net379),
    .Y(_06083_));
 sky130_fd_sc_hd__a211o_1 _11043_ (.A1(net379),
    .A2(_06082_),
    .B1(_06083_),
    .C1(_04499_),
    .X(_06084_));
 sky130_fd_sc_hd__nor2_1 _11044_ (.A(_04531_),
    .B(_04543_),
    .Y(_06085_));
 sky130_fd_sc_hd__nor2_1 _11045_ (.A(_04546_),
    .B(_04563_),
    .Y(_06086_));
 sky130_fd_sc_hd__mux2_1 _11046_ (.A0(_06085_),
    .A1(_06086_),
    .S(net379),
    .X(_06087_));
 sky130_fd_sc_hd__nor2_4 _11047_ (.A(net395),
    .B(net388),
    .Y(_06088_));
 sky130_fd_sc_hd__nand2_8 _11048_ (.A(net399),
    .B(net384),
    .Y(_06089_));
 sky130_fd_sc_hd__o221a_1 _11049_ (.A1(net399),
    .A2(_06081_),
    .B1(_06087_),
    .B2(_06089_),
    .C1(_06084_),
    .X(_06090_));
 sky130_fd_sc_hd__nor2_1 _11050_ (.A(net391),
    .B(_06090_),
    .Y(_06091_));
 sky130_fd_sc_hd__a211o_1 _11051_ (.A1(net391),
    .A2(_06073_),
    .B1(_06091_),
    .C1(_06026_),
    .X(_06092_));
 sky130_fd_sc_hd__o21a_1 _11052_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_srl_sra[1] ),
    .A2(net412),
    .B1(_06092_),
    .X(_01578_));
 sky130_fd_sc_hd__mux2_1 _11053_ (.A0(_05996_),
    .A1(_06005_),
    .S(_04488_),
    .X(_06093_));
 sky130_fd_sc_hd__nand2_4 _11054_ (.A(net631),
    .B(_05614_),
    .Y(_06094_));
 sky130_fd_sc_hd__inv_2 _11055_ (.A(_06094_),
    .Y(_06095_));
 sky130_fd_sc_hd__mux2_1 _11056_ (.A0(_06002_),
    .A1(_06095_),
    .S(net378),
    .X(_06096_));
 sky130_fd_sc_hd__mux2_2 _11057_ (.A0(_06093_),
    .A1(_06096_),
    .S(net385),
    .X(_06097_));
 sky130_fd_sc_hd__inv_2 _11058_ (.A(_06097_),
    .Y(_06098_));
 sky130_fd_sc_hd__mux2_1 _11059_ (.A0(_06010_),
    .A1(_06020_),
    .S(net378),
    .X(_06099_));
 sky130_fd_sc_hd__mux2_1 _11060_ (.A0(_06000_),
    .A1(_06017_),
    .S(net383),
    .X(_06100_));
 sky130_fd_sc_hd__inv_2 _11061_ (.A(_06100_),
    .Y(_06101_));
 sky130_fd_sc_hd__mux2_1 _11062_ (.A0(_06099_),
    .A1(_06100_),
    .S(net385),
    .X(_06102_));
 sky130_fd_sc_hd__mux2_2 _11063_ (.A0(_06098_),
    .A1(_06102_),
    .S(net398),
    .X(_06103_));
 sky130_fd_sc_hd__nor2_1 _11064_ (.A(net393),
    .B(_06103_),
    .Y(_06104_));
 sky130_fd_sc_hd__mux2_1 _11065_ (.A0(_06027_),
    .A1(_06033_),
    .S(net378),
    .X(_06105_));
 sky130_fd_sc_hd__mux2_1 _11066_ (.A0(_06013_),
    .A1(_06032_),
    .S(net381),
    .X(_06106_));
 sky130_fd_sc_hd__mux2_2 _11067_ (.A0(_06105_),
    .A1(_06106_),
    .S(net385),
    .X(_06107_));
 sky130_fd_sc_hd__a21o_1 _11068_ (.A1(net380),
    .A2(_06037_),
    .B1(_04499_),
    .X(_06108_));
 sky130_fd_sc_hd__a21o_1 _11069_ (.A1(net379),
    .A2(_06041_),
    .B1(_06108_),
    .X(_06109_));
 sky130_fd_sc_hd__mux2_2 _11070_ (.A0(_06028_),
    .A1(_06040_),
    .S(net380),
    .X(_06110_));
 sky130_fd_sc_hd__o221a_1 _11071_ (.A1(net399),
    .A2(_06107_),
    .B1(_06110_),
    .B2(_06089_),
    .C1(_06109_),
    .X(_06111_));
 sky130_fd_sc_hd__o21ai_1 _11072_ (.A1(net391),
    .A2(_06111_),
    .B1(net412),
    .Y(_06112_));
 sky130_fd_sc_hd__o22a_1 _11073_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_srl_sra[2] ),
    .A2(net412),
    .B1(_06104_),
    .B2(_06112_),
    .X(_01579_));
 sky130_fd_sc_hd__mux2_1 _11074_ (.A0(_06058_),
    .A1(_06068_),
    .S(net378),
    .X(_06113_));
 sky130_fd_sc_hd__and3_1 _11075_ (.A(net378),
    .B(_06049_),
    .C(_06050_),
    .X(_06114_));
 sky130_fd_sc_hd__a21o_1 _11076_ (.A1(net382),
    .A2(_06065_),
    .B1(_06114_),
    .X(_06115_));
 sky130_fd_sc_hd__mux2_1 _11077_ (.A0(_06113_),
    .A1(_06115_),
    .S(net384),
    .X(_06116_));
 sky130_fd_sc_hd__o21ai_4 _11078_ (.A1(net631),
    .A2(_04492_),
    .B1(net384),
    .Y(_06117_));
 sky130_fd_sc_hd__nor2_1 _11079_ (.A(net382),
    .B(_06055_),
    .Y(_06118_));
 sky130_fd_sc_hd__a31o_2 _11080_ (.A1(net382),
    .A2(_06046_),
    .A3(_06047_),
    .B1(_06118_),
    .X(_06119_));
 sky130_fd_sc_hd__o22ai_4 _11081_ (.A1(_05615_),
    .A2(_06117_),
    .B1(_06119_),
    .B2(net384),
    .Y(_06120_));
 sky130_fd_sc_hd__inv_2 _11082_ (.A(_06120_),
    .Y(_06121_));
 sky130_fd_sc_hd__mux2_1 _11083_ (.A0(_06116_),
    .A1(_06121_),
    .S(net394),
    .X(_06122_));
 sky130_fd_sc_hd__mux2_1 _11084_ (.A0(_06061_),
    .A1(_06079_),
    .S(net381),
    .X(_06123_));
 sky130_fd_sc_hd__mux2_1 _11085_ (.A0(_06075_),
    .A1(_06077_),
    .S(net378),
    .X(_06124_));
 sky130_fd_sc_hd__mux2_1 _11086_ (.A0(_06123_),
    .A1(_06124_),
    .S(net386),
    .X(_06125_));
 sky130_fd_sc_hd__mux2_1 _11087_ (.A0(_06082_),
    .A1(_06085_),
    .S(net379),
    .X(_06126_));
 sky130_fd_sc_hd__mux2_1 _11088_ (.A0(_06074_),
    .A1(_06086_),
    .S(net380),
    .X(_06127_));
 sky130_fd_sc_hd__o221a_1 _11089_ (.A1(_04499_),
    .A2(_06126_),
    .B1(_06127_),
    .B2(_06089_),
    .C1(net393),
    .X(_06128_));
 sky130_fd_sc_hd__o21ai_1 _11090_ (.A1(net399),
    .A2(_06125_),
    .B1(_06128_),
    .Y(_06129_));
 sky130_fd_sc_hd__a21oi_1 _11091_ (.A1(net391),
    .A2(_06122_),
    .B1(_06026_),
    .Y(_06130_));
 sky130_fd_sc_hd__a22o_1 _11092_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_srl_sra[3] ),
    .A2(_06026_),
    .B1(_06129_),
    .B2(_06130_),
    .X(_01580_));
 sky130_fd_sc_hd__mux2_2 _11093_ (.A0(_06001_),
    .A1(_06022_),
    .S(net387),
    .X(_06131_));
 sky130_fd_sc_hd__nor2_2 _11094_ (.A(net387),
    .B(_06094_),
    .Y(_06132_));
 sky130_fd_sc_hd__a21o_1 _11095_ (.A1(net387),
    .A2(_06006_),
    .B1(_06132_),
    .X(_06133_));
 sky130_fd_sc_hd__or2_2 _11096_ (.A(net398),
    .B(_06133_),
    .X(_06134_));
 sky130_fd_sc_hd__o21ai_4 _11097_ (.A1(net395),
    .A2(_06131_),
    .B1(_06134_),
    .Y(_06135_));
 sky130_fd_sc_hd__mux2_1 _11098_ (.A0(_06015_),
    .A1(_06035_),
    .S(net386),
    .X(_06136_));
 sky130_fd_sc_hd__a21oi_1 _11099_ (.A1(_06030_),
    .A2(_06088_),
    .B1(net389),
    .Y(_06137_));
 sky130_fd_sc_hd__o2bb2a_1 _11100_ (.A1_N(net394),
    .A2_N(_06136_),
    .B1(_06042_),
    .B2(_04499_),
    .X(_06138_));
 sky130_fd_sc_hd__a221o_1 _11101_ (.A1(net389),
    .A2(_06135_),
    .B1(_06137_),
    .B2(_06138_),
    .C1(_06026_),
    .X(_06139_));
 sky130_fd_sc_hd__a21bo_1 _11102_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_srl_sra[4] ),
    .A2(_06026_),
    .B1_N(_06139_),
    .X(_01581_));
 sky130_fd_sc_hd__mux2_1 _11103_ (.A0(_06051_),
    .A1(_06070_),
    .S(net387),
    .X(_06140_));
 sky130_fd_sc_hd__a21o_1 _11104_ (.A1(net387),
    .A2(_06056_),
    .B1(_06132_),
    .X(_06141_));
 sky130_fd_sc_hd__or2_1 _11105_ (.A(net398),
    .B(_06141_),
    .X(_06142_));
 sky130_fd_sc_hd__o21ai_2 _11106_ (.A1(net394),
    .A2(_06140_),
    .B1(_06142_),
    .Y(_06143_));
 sky130_fd_sc_hd__mux2_2 _11107_ (.A0(_06062_),
    .A1(_06080_),
    .S(net387),
    .X(_06144_));
 sky130_fd_sc_hd__o221a_1 _11108_ (.A1(_04499_),
    .A2(_06087_),
    .B1(_06089_),
    .B2(_06076_),
    .C1(net393),
    .X(_06145_));
 sky130_fd_sc_hd__o21ai_1 _11109_ (.A1(net399),
    .A2(_06144_),
    .B1(_06145_),
    .Y(_06146_));
 sky130_fd_sc_hd__a21oi_1 _11110_ (.A1(net391),
    .A2(_06143_),
    .B1(_06026_),
    .Y(_06147_));
 sky130_fd_sc_hd__a22o_1 _11111_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_srl_sra[5] ),
    .A2(_06026_),
    .B1(_06146_),
    .B2(_06147_),
    .X(_01582_));
 sky130_fd_sc_hd__mux2_1 _11112_ (.A0(_06093_),
    .A1(_06101_),
    .S(net386),
    .X(_06148_));
 sky130_fd_sc_hd__a21o_1 _11113_ (.A1(net387),
    .A2(_06096_),
    .B1(_06132_),
    .X(_06149_));
 sky130_fd_sc_hd__mux2_1 _11114_ (.A0(_06148_),
    .A1(_06149_),
    .S(net395),
    .X(_06150_));
 sky130_fd_sc_hd__mux2_1 _11115_ (.A0(_06099_),
    .A1(_06106_),
    .S(net387),
    .X(_06151_));
 sky130_fd_sc_hd__o221a_1 _11116_ (.A1(_06089_),
    .A2(_06105_),
    .B1(_06110_),
    .B2(_04499_),
    .C1(net392),
    .X(_06152_));
 sky130_fd_sc_hd__o21ai_1 _11117_ (.A1(net398),
    .A2(_06151_),
    .B1(_06152_),
    .Y(_06153_));
 sky130_fd_sc_hd__o211a_1 _11118_ (.A1(net392),
    .A2(_06150_),
    .B1(_06153_),
    .C1(net412),
    .X(_06154_));
 sky130_fd_sc_hd__a21o_1 _11119_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_srl_sra[6] ),
    .A2(_06026_),
    .B1(_06154_),
    .X(_01583_));
 sky130_fd_sc_hd__a31o_1 _11120_ (.A1(net388),
    .A2(net380),
    .A3(net377),
    .B1(net631),
    .X(_06155_));
 sky130_fd_sc_hd__nand2_1 _11121_ (.A(net395),
    .B(_06155_),
    .Y(_06156_));
 sky130_fd_sc_hd__mux2_1 _11122_ (.A0(_06115_),
    .A1(_06119_),
    .S(net385),
    .X(_06157_));
 sky130_fd_sc_hd__o22a_1 _11123_ (.A1(_05615_),
    .A2(_06156_),
    .B1(_06157_),
    .B2(net395),
    .X(_06158_));
 sky130_fd_sc_hd__mux2_1 _11124_ (.A0(_06113_),
    .A1(_06123_),
    .S(net386),
    .X(_06159_));
 sky130_fd_sc_hd__a221o_1 _11125_ (.A1(_06088_),
    .A2(_06124_),
    .B1(_06127_),
    .B2(_04498_),
    .C1(net391),
    .X(_06160_));
 sky130_fd_sc_hd__a21o_1 _11126_ (.A1(net395),
    .A2(_06159_),
    .B1(_06160_),
    .X(_06161_));
 sky130_fd_sc_hd__o211a_1 _11127_ (.A1(net393),
    .A2(_06158_),
    .B1(_06161_),
    .C1(net412),
    .X(_06162_));
 sky130_fd_sc_hd__o21ba_1 _11128_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_srl_sra[7] ),
    .A2(net412),
    .B1_N(_06162_),
    .X(_01584_));
 sky130_fd_sc_hd__nor2_4 _11129_ (.A(net398),
    .B(_06094_),
    .Y(_06163_));
 sky130_fd_sc_hd__a21oi_1 _11130_ (.A1(net398),
    .A2(_06007_),
    .B1(_06163_),
    .Y(_06164_));
 sky130_fd_sc_hd__nand2_1 _11131_ (.A(net390),
    .B(_06164_),
    .Y(_06165_));
 sky130_fd_sc_hd__mux2_1 _11132_ (.A0(_06023_),
    .A1(_06036_),
    .S(net396),
    .X(_06166_));
 sky130_fd_sc_hd__o21a_1 _11133_ (.A1(net389),
    .A2(_06166_),
    .B1(net412),
    .X(_06167_));
 sky130_fd_sc_hd__a22o_1 _11134_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_srl_sra[8] ),
    .A2(_06026_),
    .B1(_06165_),
    .B2(_06167_),
    .X(_01585_));
 sky130_fd_sc_hd__a21oi_1 _11135_ (.A1(net398),
    .A2(_06057_),
    .B1(_06163_),
    .Y(_06168_));
 sky130_fd_sc_hd__or2_1 _11136_ (.A(net394),
    .B(_06081_),
    .X(_06169_));
 sky130_fd_sc_hd__o211a_1 _11137_ (.A1(net398),
    .A2(_06071_),
    .B1(_06169_),
    .C1(net392),
    .X(_06170_));
 sky130_fd_sc_hd__a21oi_1 _11138_ (.A1(net389),
    .A2(_06168_),
    .B1(_06170_),
    .Y(_06171_));
 sky130_fd_sc_hd__mux2_1 _11139_ (.A0(\core_pipeline.pipeline_execute.ex_alu.result_srl_sra[9] ),
    .A1(_06171_),
    .S(net413),
    .X(_01586_));
 sky130_fd_sc_hd__a21oi_2 _11140_ (.A1(net399),
    .A2(_06097_),
    .B1(_06163_),
    .Y(_06172_));
 sky130_fd_sc_hd__nand2_1 _11141_ (.A(net389),
    .B(_06172_),
    .Y(_06173_));
 sky130_fd_sc_hd__mux2_1 _11142_ (.A0(_06102_),
    .A1(_06107_),
    .S(net396),
    .X(_06174_));
 sky130_fd_sc_hd__a21oi_1 _11143_ (.A1(net392),
    .A2(_06174_),
    .B1(_06026_),
    .Y(_06175_));
 sky130_fd_sc_hd__a22o_1 _11144_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_srl_sra[10] ),
    .A2(_06026_),
    .B1(_06173_),
    .B2(_06175_),
    .X(_01587_));
 sky130_fd_sc_hd__a21oi_1 _11145_ (.A1(net398),
    .A2(_06120_),
    .B1(_06163_),
    .Y(_06176_));
 sky130_fd_sc_hd__nand2_1 _11146_ (.A(net390),
    .B(_06176_),
    .Y(_06177_));
 sky130_fd_sc_hd__mux2_1 _11147_ (.A0(_06116_),
    .A1(_06125_),
    .S(net399),
    .X(_06178_));
 sky130_fd_sc_hd__a21oi_1 _11148_ (.A1(net392),
    .A2(_06178_),
    .B1(_06026_),
    .Y(_06179_));
 sky130_fd_sc_hd__a22o_1 _11149_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_srl_sra[11] ),
    .A2(_06026_),
    .B1(_06177_),
    .B2(_06179_),
    .X(_01588_));
 sky130_fd_sc_hd__a21oi_1 _11150_ (.A1(net398),
    .A2(_06133_),
    .B1(_06163_),
    .Y(_06180_));
 sky130_fd_sc_hd__nand2_1 _11151_ (.A(net390),
    .B(_06180_),
    .Y(_06181_));
 sky130_fd_sc_hd__mux2_1 _11152_ (.A0(_06131_),
    .A1(_06136_),
    .S(net396),
    .X(_06182_));
 sky130_fd_sc_hd__o211a_1 _11153_ (.A1(net389),
    .A2(_06182_),
    .B1(_06181_),
    .C1(net412),
    .X(_06183_));
 sky130_fd_sc_hd__a21o_1 _11154_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_srl_sra[12] ),
    .A2(_06026_),
    .B1(_06183_),
    .X(_01589_));
 sky130_fd_sc_hd__a21oi_2 _11155_ (.A1(net398),
    .A2(_06141_),
    .B1(_06163_),
    .Y(_06184_));
 sky130_fd_sc_hd__nand2_1 _11156_ (.A(net394),
    .B(_06140_),
    .Y(_06185_));
 sky130_fd_sc_hd__o211a_1 _11157_ (.A1(net394),
    .A2(_06144_),
    .B1(_06185_),
    .C1(net393),
    .X(_06186_));
 sky130_fd_sc_hd__a21oi_2 _11158_ (.A1(net390),
    .A2(_06184_),
    .B1(_06186_),
    .Y(_06187_));
 sky130_fd_sc_hd__mux2_1 _11159_ (.A0(\core_pipeline.pipeline_execute.ex_alu.result_srl_sra[13] ),
    .A1(_06187_),
    .S(net413),
    .X(_01590_));
 sky130_fd_sc_hd__a21oi_2 _11160_ (.A1(net398),
    .A2(_06149_),
    .B1(_06163_),
    .Y(_06188_));
 sky130_fd_sc_hd__nor2_1 _11161_ (.A(net394),
    .B(_06151_),
    .Y(_06189_));
 sky130_fd_sc_hd__a21o_1 _11162_ (.A1(net395),
    .A2(_06148_),
    .B1(net390),
    .X(_06190_));
 sky130_fd_sc_hd__o2bb2a_1 _11163_ (.A1_N(net390),
    .A2_N(_06188_),
    .B1(_06189_),
    .B2(_06190_),
    .X(_06191_));
 sky130_fd_sc_hd__mux2_1 _11164_ (.A0(\core_pipeline.pipeline_execute.ex_alu.result_srl_sra[14] ),
    .A1(_06191_),
    .S(net413),
    .X(_01591_));
 sky130_fd_sc_hd__mux2_1 _11165_ (.A0(_06157_),
    .A1(_06159_),
    .S(net399),
    .X(_06192_));
 sky130_fd_sc_hd__a41o_4 _11166_ (.A1(net399),
    .A2(net388),
    .A3(net380),
    .A4(net377),
    .B1(net631),
    .X(_06193_));
 sky130_fd_sc_hd__a21oi_1 _11167_ (.A1(_05614_),
    .A2(_06193_),
    .B1(net393),
    .Y(_06194_));
 sky130_fd_sc_hd__a21oi_2 _11168_ (.A1(net393),
    .A2(_06192_),
    .B1(_06194_),
    .Y(_06195_));
 sky130_fd_sc_hd__mux2_1 _11169_ (.A0(\core_pipeline.pipeline_execute.ex_alu.result_srl_sra[15] ),
    .A1(_06195_),
    .S(net412),
    .X(_01592_));
 sky130_fd_sc_hd__a31o_4 _11170_ (.A1(net631),
    .A2(net391),
    .A3(_05614_),
    .B1(_06026_),
    .X(_06196_));
 sky130_fd_sc_hd__a21o_1 _11171_ (.A1(net392),
    .A2(_06024_),
    .B1(_06196_),
    .X(_06197_));
 sky130_fd_sc_hd__o21a_1 _11172_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_srl_sra[16] ),
    .A2(net413),
    .B1(_06197_),
    .X(_01593_));
 sky130_fd_sc_hd__a21o_1 _11173_ (.A1(net393),
    .A2(_06073_),
    .B1(_06196_),
    .X(_06198_));
 sky130_fd_sc_hd__o21a_1 _11174_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_srl_sra[17] ),
    .A2(net413),
    .B1(_06198_),
    .X(_01594_));
 sky130_fd_sc_hd__nor2_1 _11175_ (.A(net390),
    .B(_06103_),
    .Y(_06199_));
 sky130_fd_sc_hd__o22a_1 _11176_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_srl_sra[18] ),
    .A2(net413),
    .B1(_06196_),
    .B2(_06199_),
    .X(_01595_));
 sky130_fd_sc_hd__nor2_1 _11177_ (.A(net391),
    .B(_06122_),
    .Y(_06200_));
 sky130_fd_sc_hd__o22a_1 _11178_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_srl_sra[19] ),
    .A2(net412),
    .B1(_06196_),
    .B2(_06200_),
    .X(_01596_));
 sky130_fd_sc_hd__nor2_1 _11179_ (.A(net390),
    .B(_06135_),
    .Y(_06201_));
 sky130_fd_sc_hd__o22a_1 _11180_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_srl_sra[20] ),
    .A2(net412),
    .B1(_06196_),
    .B2(_06201_),
    .X(_01597_));
 sky130_fd_sc_hd__nor2_1 _11181_ (.A(net390),
    .B(_06143_),
    .Y(_06202_));
 sky130_fd_sc_hd__o22a_1 _11182_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_srl_sra[21] ),
    .A2(net413),
    .B1(_06196_),
    .B2(_06202_),
    .X(_01598_));
 sky130_fd_sc_hd__a21o_1 _11183_ (.A1(net392),
    .A2(_06150_),
    .B1(_06196_),
    .X(_06203_));
 sky130_fd_sc_hd__o21a_1 _11184_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_srl_sra[22] ),
    .A2(net412),
    .B1(_06203_),
    .X(_01599_));
 sky130_fd_sc_hd__nor2_1 _11185_ (.A(net391),
    .B(_06158_),
    .Y(_06204_));
 sky130_fd_sc_hd__o22a_1 _11186_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_srl_sra[23] ),
    .A2(net412),
    .B1(_06196_),
    .B2(_06204_),
    .X(_01600_));
 sky130_fd_sc_hd__nor2_1 _11187_ (.A(net390),
    .B(_06164_),
    .Y(_06205_));
 sky130_fd_sc_hd__o22a_1 _11188_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_srl_sra[24] ),
    .A2(net413),
    .B1(_06196_),
    .B2(_06205_),
    .X(_01601_));
 sky130_fd_sc_hd__nor2_1 _11189_ (.A(net390),
    .B(_06168_),
    .Y(_06206_));
 sky130_fd_sc_hd__o22a_1 _11190_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_srl_sra[25] ),
    .A2(net413),
    .B1(_06196_),
    .B2(_06206_),
    .X(_01602_));
 sky130_fd_sc_hd__nor2_1 _11191_ (.A(net390),
    .B(_06172_),
    .Y(_06207_));
 sky130_fd_sc_hd__o22a_1 _11192_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_srl_sra[26] ),
    .A2(net413),
    .B1(_06196_),
    .B2(_06207_),
    .X(_01603_));
 sky130_fd_sc_hd__nor2_1 _11193_ (.A(net390),
    .B(_06176_),
    .Y(_06208_));
 sky130_fd_sc_hd__o22a_1 _11194_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_srl_sra[27] ),
    .A2(net413),
    .B1(_06196_),
    .B2(_06208_),
    .X(_01604_));
 sky130_fd_sc_hd__nor2_1 _11195_ (.A(net390),
    .B(_06180_),
    .Y(_06209_));
 sky130_fd_sc_hd__o22a_1 _11196_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_srl_sra[28] ),
    .A2(net413),
    .B1(_06196_),
    .B2(_06209_),
    .X(_01605_));
 sky130_fd_sc_hd__nor2_1 _11197_ (.A(net390),
    .B(_06184_),
    .Y(_06210_));
 sky130_fd_sc_hd__o22a_1 _11198_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_srl_sra[29] ),
    .A2(net412),
    .B1(_06196_),
    .B2(_06210_),
    .X(_01606_));
 sky130_fd_sc_hd__nor2_1 _11199_ (.A(net390),
    .B(_06188_),
    .Y(_06211_));
 sky130_fd_sc_hd__o22a_1 _11200_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_srl_sra[30] ),
    .A2(net412),
    .B1(_06196_),
    .B2(_06211_),
    .X(_01607_));
 sky130_fd_sc_hd__nand2_1 _11201_ (.A(net459),
    .B(net391),
    .Y(_06212_));
 sky130_fd_sc_hd__and3_1 _11202_ (.A(net412),
    .B(_06193_),
    .C(_06212_),
    .X(_06213_));
 sky130_fd_sc_hd__a22o_1 _11203_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_srl_sra[31] ),
    .A2(_06026_),
    .B1(_06213_),
    .B2(_05614_),
    .X(_01608_));
 sky130_fd_sc_hd__or3b_2 _11204_ (.A(\core_pipeline.decode_to_execute_alu_function[1] ),
    .B(\core_pipeline.decode_to_execute_alu_function[0] ),
    .C_N(\core_pipeline.decode_to_execute_alu_function[2] ),
    .X(_06214_));
 sky130_fd_sc_hd__mux2_1 _11205_ (.A0(_05816_),
    .A1(\core_pipeline.pipeline_execute.ex_alu.result_xor[0] ),
    .S(net411),
    .X(_01609_));
 sky130_fd_sc_hd__mux2_1 _11206_ (.A0(_05819_),
    .A1(\core_pipeline.pipeline_execute.ex_alu.result_xor[1] ),
    .S(net411),
    .X(_01610_));
 sky130_fd_sc_hd__mux2_1 _11207_ (.A0(_05815_),
    .A1(\core_pipeline.pipeline_execute.ex_alu.result_xor[2] ),
    .S(net411),
    .X(_01611_));
 sky130_fd_sc_hd__mux2_1 _11208_ (.A0(_05814_),
    .A1(\core_pipeline.pipeline_execute.ex_alu.result_xor[3] ),
    .S(net411),
    .X(_01612_));
 sky130_fd_sc_hd__mux2_1 _11209_ (.A0(_05674_),
    .A1(\core_pipeline.pipeline_execute.ex_alu.result_xor[4] ),
    .S(net411),
    .X(_01613_));
 sky130_fd_sc_hd__mux2_1 _11210_ (.A0(_05675_),
    .A1(\core_pipeline.pipeline_execute.ex_alu.result_xor[5] ),
    .S(net411),
    .X(_01614_));
 sky130_fd_sc_hd__mux2_1 _11211_ (.A0(_05663_),
    .A1(\core_pipeline.pipeline_execute.ex_alu.result_xor[6] ),
    .S(net411),
    .X(_01615_));
 sky130_fd_sc_hd__mux2_1 _11212_ (.A0(_05660_),
    .A1(\core_pipeline.pipeline_execute.ex_alu.result_xor[7] ),
    .S(net411),
    .X(_01616_));
 sky130_fd_sc_hd__mux2_1 _11213_ (.A0(_05634_),
    .A1(\core_pipeline.pipeline_execute.ex_alu.result_xor[8] ),
    .S(net410),
    .X(_01617_));
 sky130_fd_sc_hd__mux2_1 _11214_ (.A0(_05637_),
    .A1(\core_pipeline.pipeline_execute.ex_alu.result_xor[9] ),
    .S(net410),
    .X(_01618_));
 sky130_fd_sc_hd__mux2_1 _11215_ (.A0(_05654_),
    .A1(\core_pipeline.pipeline_execute.ex_alu.result_xor[10] ),
    .S(net410),
    .X(_01619_));
 sky130_fd_sc_hd__mux2_1 _11216_ (.A0(_05640_),
    .A1(\core_pipeline.pipeline_execute.ex_alu.result_xor[11] ),
    .S(net410),
    .X(_01620_));
 sky130_fd_sc_hd__mux2_1 _11217_ (.A0(_05646_),
    .A1(\core_pipeline.pipeline_execute.ex_alu.result_xor[12] ),
    .S(net410),
    .X(_01621_));
 sky130_fd_sc_hd__nand2b_1 _11218_ (.A_N(\core_pipeline.pipeline_execute.ex_alu.result_xor[13] ),
    .B(net410),
    .Y(_06215_));
 sky130_fd_sc_hd__o31a_1 _11219_ (.A1(_05624_),
    .A2(_05649_),
    .A3(net410),
    .B1(_06215_),
    .X(_01622_));
 sky130_fd_sc_hd__mux2_1 _11220_ (.A0(_05621_),
    .A1(\core_pipeline.pipeline_execute.ex_alu.result_xor[14] ),
    .S(net410),
    .X(_01623_));
 sky130_fd_sc_hd__mux2_1 _11221_ (.A0(_05630_),
    .A1(\core_pipeline.pipeline_execute.ex_alu.result_xor[15] ),
    .S(net410),
    .X(_01624_));
 sky130_fd_sc_hd__mux2_1 _11222_ (.A0(_05761_),
    .A1(\core_pipeline.pipeline_execute.ex_alu.result_xor[16] ),
    .S(net410),
    .X(_01625_));
 sky130_fd_sc_hd__mux2_1 _11223_ (.A0(_05749_),
    .A1(\core_pipeline.pipeline_execute.ex_alu.result_xor[17] ),
    .S(net410),
    .X(_01626_));
 sky130_fd_sc_hd__mux2_1 _11224_ (.A0(_05784_),
    .A1(\core_pipeline.pipeline_execute.ex_alu.result_xor[18] ),
    .S(net410),
    .X(_01627_));
 sky130_fd_sc_hd__mux2_1 _11225_ (.A0(_05791_),
    .A1(\core_pipeline.pipeline_execute.ex_alu.result_xor[19] ),
    .S(net410),
    .X(_01628_));
 sky130_fd_sc_hd__mux2_1 _11226_ (.A0(_05777_),
    .A1(\core_pipeline.pipeline_execute.ex_alu.result_xor[20] ),
    .S(net410),
    .X(_01629_));
 sky130_fd_sc_hd__mux2_1 _11227_ (.A0(_05769_),
    .A1(\core_pipeline.pipeline_execute.ex_alu.result_xor[21] ),
    .S(net411),
    .X(_01630_));
 sky130_fd_sc_hd__mux2_1 _11228_ (.A0(_05756_),
    .A1(\core_pipeline.pipeline_execute.ex_alu.result_xor[22] ),
    .S(net411),
    .X(_01631_));
 sky130_fd_sc_hd__mux2_1 _11229_ (.A0(_05743_),
    .A1(\core_pipeline.pipeline_execute.ex_alu.result_xor[23] ),
    .S(net411),
    .X(_01632_));
 sky130_fd_sc_hd__mux2_1 _11230_ (.A0(_05720_),
    .A1(\core_pipeline.pipeline_execute.ex_alu.result_xor[24] ),
    .S(net410),
    .X(_01633_));
 sky130_fd_sc_hd__mux2_1 _11231_ (.A0(_05734_),
    .A1(\core_pipeline.pipeline_execute.ex_alu.result_xor[25] ),
    .S(net410),
    .X(_01634_));
 sky130_fd_sc_hd__mux2_1 _11232_ (.A0(_05713_),
    .A1(\core_pipeline.pipeline_execute.ex_alu.result_xor[26] ),
    .S(net410),
    .X(_01635_));
 sky130_fd_sc_hd__mux2_1 _11233_ (.A0(_05727_),
    .A1(\core_pipeline.pipeline_execute.ex_alu.result_xor[27] ),
    .S(net411),
    .X(_01636_));
 sky130_fd_sc_hd__mux2_1 _11234_ (.A0(_05700_),
    .A1(\core_pipeline.pipeline_execute.ex_alu.result_xor[28] ),
    .S(net411),
    .X(_01637_));
 sky130_fd_sc_hd__mux2_1 _11235_ (.A0(_05708_),
    .A1(\core_pipeline.pipeline_execute.ex_alu.result_xor[29] ),
    .S(net411),
    .X(_01638_));
 sky130_fd_sc_hd__mux2_1 _11236_ (.A0(_05694_),
    .A1(\core_pipeline.pipeline_execute.ex_alu.result_xor[30] ),
    .S(net411),
    .X(_01639_));
 sky130_fd_sc_hd__mux2_1 _11237_ (.A0(_05685_),
    .A1(\core_pipeline.pipeline_execute.ex_alu.result_xor[31] ),
    .S(net411),
    .X(_01640_));
 sky130_fd_sc_hd__or3b_1 _11238_ (.A(\core_pipeline.decode_to_execute_alu_function[2] ),
    .B(\core_pipeline.decode_to_execute_alu_function[0] ),
    .C_N(\core_pipeline.decode_to_execute_alu_function[1] ),
    .X(_06216_));
 sky130_fd_sc_hd__nand2b_1 _11239_ (.A_N(_05685_),
    .B(_05813_),
    .Y(_06217_));
 sky130_fd_sc_hd__nor2_1 _11240_ (.A(_05823_),
    .B(_06216_),
    .Y(_06218_));
 sky130_fd_sc_hd__a32o_1 _11241_ (.A1(_05616_),
    .A2(_06217_),
    .A3(_06218_),
    .B1(_06216_),
    .B2(\core_pipeline.pipeline_execute.ex_alu.result_slt[0] ),
    .X(_01641_));
 sky130_fd_sc_hd__nor2_1 _11242_ (.A(_06012_),
    .B(_06031_),
    .Y(_06219_));
 sky130_fd_sc_hd__mux2_1 _11243_ (.A0(_04610_),
    .A1(_06219_),
    .S(net381),
    .X(_06220_));
 sky130_fd_sc_hd__mux2_1 _11244_ (.A0(_04593_),
    .A1(_06220_),
    .S(net386),
    .X(_06221_));
 sky130_fd_sc_hd__nand2_1 _11245_ (.A(net396),
    .B(_06221_),
    .Y(_06222_));
 sky130_fd_sc_hd__o211a_1 _11246_ (.A1(net396),
    .A2(_04560_),
    .B1(_06222_),
    .C1(net392),
    .X(_06223_));
 sky130_fd_sc_hd__a31o_1 _11247_ (.A1(net391),
    .A2(_04495_),
    .A3(_04500_),
    .B1(net435),
    .X(_06224_));
 sky130_fd_sc_hd__o22a_1 _11248_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_sll[16] ),
    .A2(_04471_),
    .B1(_06223_),
    .B2(_06224_),
    .X(_01642_));
 sky130_fd_sc_hd__nor2_1 _11249_ (.A(_06060_),
    .B(_06078_),
    .Y(_06225_));
 sky130_fd_sc_hd__mux2_1 _11250_ (.A0(_04619_),
    .A1(_06225_),
    .S(net381),
    .X(_06226_));
 sky130_fd_sc_hd__inv_2 _11251_ (.A(_06226_),
    .Y(_06227_));
 sky130_fd_sc_hd__nor2_1 _11252_ (.A(net385),
    .B(_06226_),
    .Y(_06228_));
 sky130_fd_sc_hd__a21oi_1 _11253_ (.A1(net385),
    .A2(_04603_),
    .B1(_06228_),
    .Y(_06229_));
 sky130_fd_sc_hd__nand2_1 _11254_ (.A(net396),
    .B(_06229_),
    .Y(_06230_));
 sky130_fd_sc_hd__o211a_1 _11255_ (.A1(net396),
    .A2(_04570_),
    .B1(_06230_),
    .C1(net392),
    .X(_06231_));
 sky130_fd_sc_hd__a31o_1 _11256_ (.A1(net389),
    .A2(_04498_),
    .A3(_04507_),
    .B1(net436),
    .X(_06232_));
 sky130_fd_sc_hd__o22a_1 _11257_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_sll[17] ),
    .A2(net437),
    .B1(_06231_),
    .B2(_06232_),
    .X(_01643_));
 sky130_fd_sc_hd__nor2_1 _11258_ (.A(_06009_),
    .B(_06011_),
    .Y(_06233_));
 sky130_fd_sc_hd__mux2_1 _11259_ (.A0(_06219_),
    .A1(_06233_),
    .S(net382),
    .X(_06234_));
 sky130_fd_sc_hd__mux2_1 _11260_ (.A0(_04611_),
    .A1(_06234_),
    .S(net386),
    .X(_06235_));
 sky130_fd_sc_hd__mux2_1 _11261_ (.A0(_04577_),
    .A1(_06235_),
    .S(net397),
    .X(_06236_));
 sky130_fd_sc_hd__nor2_1 _11262_ (.A(net389),
    .B(_06236_),
    .Y(_06237_));
 sky130_fd_sc_hd__a31o_1 _11263_ (.A1(net389),
    .A2(_04498_),
    .A3(_04514_),
    .B1(net436),
    .X(_06238_));
 sky130_fd_sc_hd__o22a_1 _11264_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_sll[18] ),
    .A2(net437),
    .B1(_06237_),
    .B2(_06238_),
    .X(_01644_));
 sky130_fd_sc_hd__o21ba_1 _11265_ (.A1(net372),
    .A2(_05788_),
    .B1_N(_06059_),
    .X(_06239_));
 sky130_fd_sc_hd__mux2_1 _11266_ (.A0(_06225_),
    .A1(_06239_),
    .S(net381),
    .X(_06240_));
 sky130_fd_sc_hd__mux2_1 _11267_ (.A0(_04620_),
    .A1(_06240_),
    .S(net386),
    .X(_06241_));
 sky130_fd_sc_hd__nand2_1 _11268_ (.A(net396),
    .B(_06241_),
    .Y(_06242_));
 sky130_fd_sc_hd__o211a_1 _11269_ (.A1(net396),
    .A2(_04586_),
    .B1(_06242_),
    .C1(net392),
    .X(_06243_));
 sky130_fd_sc_hd__a31o_1 _11270_ (.A1(net389),
    .A2(_04498_),
    .A3(_04520_),
    .B1(net435),
    .X(_06244_));
 sky130_fd_sc_hd__o22a_1 _11271_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_sll[19] ),
    .A2(net438),
    .B1(_06243_),
    .B2(_06244_),
    .X(_01645_));
 sky130_fd_sc_hd__nor2_1 _11272_ (.A(_06008_),
    .B(_06019_),
    .Y(_06245_));
 sky130_fd_sc_hd__mux2_1 _11273_ (.A0(_06233_),
    .A1(_06245_),
    .S(net381),
    .X(_06246_));
 sky130_fd_sc_hd__mux2_1 _11274_ (.A0(_06220_),
    .A1(_06246_),
    .S(net386),
    .X(_06247_));
 sky130_fd_sc_hd__nand2_1 _11275_ (.A(net397),
    .B(_06247_),
    .Y(_06248_));
 sky130_fd_sc_hd__o211a_1 _11276_ (.A1(net397),
    .A2(_04595_),
    .B1(_06248_),
    .C1(net392),
    .X(_06249_));
 sky130_fd_sc_hd__a31o_1 _11277_ (.A1(net396),
    .A2(net389),
    .A3(_04527_),
    .B1(net436),
    .X(_06250_));
 sky130_fd_sc_hd__o22a_1 _11278_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_sll[20] ),
    .A2(net438),
    .B1(_06249_),
    .B2(_06250_),
    .X(_01646_));
 sky130_fd_sc_hd__o21ai_1 _11279_ (.A1(net375),
    .A2(_05773_),
    .B1(_06066_),
    .Y(_06251_));
 sky130_fd_sc_hd__nor2_1 _11280_ (.A(net378),
    .B(_06251_),
    .Y(_06252_));
 sky130_fd_sc_hd__a21oi_1 _11281_ (.A1(net378),
    .A2(_06239_),
    .B1(_06252_),
    .Y(_06253_));
 sky130_fd_sc_hd__mux2_1 _11282_ (.A0(_06227_),
    .A1(_06253_),
    .S(net386),
    .X(_06254_));
 sky130_fd_sc_hd__or2_1 _11283_ (.A(net396),
    .B(_04604_),
    .X(_06255_));
 sky130_fd_sc_hd__o211a_1 _11284_ (.A1(net394),
    .A2(_06254_),
    .B1(_06255_),
    .C1(net392),
    .X(_06256_));
 sky130_fd_sc_hd__a31o_1 _11285_ (.A1(net396),
    .A2(net391),
    .A3(_04534_),
    .B1(net435),
    .X(_06257_));
 sky130_fd_sc_hd__o22a_1 _11286_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_sll[21] ),
    .A2(net438),
    .B1(_06256_),
    .B2(_06257_),
    .X(_01647_));
 sky130_fd_sc_hd__and3_1 _11287_ (.A(net381),
    .B(_06016_),
    .C(_06018_),
    .X(_06258_));
 sky130_fd_sc_hd__a21o_1 _11288_ (.A1(net378),
    .A2(_06245_),
    .B1(_06258_),
    .X(_06259_));
 sky130_fd_sc_hd__mux2_1 _11289_ (.A0(_06234_),
    .A1(_06259_),
    .S(net386),
    .X(_06260_));
 sky130_fd_sc_hd__nor2_1 _11290_ (.A(net397),
    .B(_04612_),
    .Y(_06261_));
 sky130_fd_sc_hd__o21ai_1 _11291_ (.A1(net394),
    .A2(_06260_),
    .B1(net392),
    .Y(_06262_));
 sky130_fd_sc_hd__o221a_1 _11292_ (.A1(net392),
    .A2(_04542_),
    .B1(_06261_),
    .B2(_06262_),
    .C1(net438),
    .X(_06263_));
 sky130_fd_sc_hd__a21o_1 _11293_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_sll[22] ),
    .A2(net435),
    .B1(_06263_),
    .X(_01648_));
 sky130_fd_sc_hd__nand2_1 _11294_ (.A(_06064_),
    .B(_06067_),
    .Y(_06264_));
 sky130_fd_sc_hd__mux2_1 _11295_ (.A0(_06251_),
    .A1(_06264_),
    .S(net381),
    .X(_06265_));
 sky130_fd_sc_hd__inv_2 _11296_ (.A(_06265_),
    .Y(_06266_));
 sky130_fd_sc_hd__mux2_1 _11297_ (.A0(_06240_),
    .A1(_06266_),
    .S(net386),
    .X(_06267_));
 sky130_fd_sc_hd__nor2_1 _11298_ (.A(net399),
    .B(_04621_),
    .Y(_06268_));
 sky130_fd_sc_hd__o21ai_1 _11299_ (.A1(net395),
    .A2(_06267_),
    .B1(net393),
    .Y(_06269_));
 sky130_fd_sc_hd__o221a_1 _11300_ (.A1(net393),
    .A2(_04551_),
    .B1(_06268_),
    .B2(_06269_),
    .C1(net438),
    .X(_06270_));
 sky130_fd_sc_hd__a21o_1 _11301_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_sll[23] ),
    .A2(net435),
    .B1(_06270_),
    .X(_01649_));
 sky130_fd_sc_hd__nand2_4 _11302_ (.A(net437),
    .B(net389),
    .Y(_06271_));
 sky130_fd_sc_hd__inv_2 _11303_ (.A(_06271_),
    .Y(_06272_));
 sky130_fd_sc_hd__a21oi_2 _11304_ (.A1(net372),
    .A2(_05740_),
    .B1(_05999_),
    .Y(_06273_));
 sky130_fd_sc_hd__and3_1 _11305_ (.A(net378),
    .B(_06016_),
    .C(_06018_),
    .X(_06274_));
 sky130_fd_sc_hd__a21oi_1 _11306_ (.A1(net381),
    .A2(_06273_),
    .B1(_06274_),
    .Y(_06275_));
 sky130_fd_sc_hd__nor2_1 _11307_ (.A(_04499_),
    .B(_06275_),
    .Y(_06276_));
 sky130_fd_sc_hd__a221o_1 _11308_ (.A1(net394),
    .A2(_06221_),
    .B1(_06246_),
    .B2(_06088_),
    .C1(_06276_),
    .X(_06277_));
 sky130_fd_sc_hd__nand2_1 _11309_ (.A(_04481_),
    .B(_06277_),
    .Y(_06278_));
 sky130_fd_sc_hd__o221a_1 _11310_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_sll[24] ),
    .A2(net437),
    .B1(_04562_),
    .B2(_06271_),
    .C1(_06278_),
    .X(_01650_));
 sky130_fd_sc_hd__nand2_1 _11311_ (.A(net394),
    .B(_06229_),
    .Y(_06279_));
 sky130_fd_sc_hd__nand2_1 _11312_ (.A(_06049_),
    .B(_06063_),
    .Y(_06280_));
 sky130_fd_sc_hd__mux2_1 _11313_ (.A0(_06264_),
    .A1(_06280_),
    .S(net383),
    .X(_06281_));
 sky130_fd_sc_hd__o221a_1 _11314_ (.A1(_06089_),
    .A2(_06253_),
    .B1(_06281_),
    .B2(_04499_),
    .C1(_06279_),
    .X(_06282_));
 sky130_fd_sc_hd__or2_1 _11315_ (.A(_04482_),
    .B(_06282_),
    .X(_06283_));
 sky130_fd_sc_hd__o221a_1 _11316_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_sll[25] ),
    .A2(net437),
    .B1(_04571_),
    .B2(_06271_),
    .C1(_06283_),
    .X(_01651_));
 sky130_fd_sc_hd__nor2_1 _11317_ (.A(_05995_),
    .B(_05998_),
    .Y(_06284_));
 sky130_fd_sc_hd__mux2_1 _11318_ (.A0(_06273_),
    .A1(_06284_),
    .S(net381),
    .X(_06285_));
 sky130_fd_sc_hd__a221o_1 _11319_ (.A1(_06088_),
    .A2(_06259_),
    .B1(_06285_),
    .B2(_04498_),
    .C1(net389),
    .X(_06286_));
 sky130_fd_sc_hd__a21oi_1 _11320_ (.A1(net394),
    .A2(_06235_),
    .B1(_06286_),
    .Y(_06287_));
 sky130_fd_sc_hd__a211o_1 _11321_ (.A1(net389),
    .A2(_04578_),
    .B1(_06287_),
    .C1(net436),
    .X(_06288_));
 sky130_fd_sc_hd__o21a_1 _11322_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_sll[26] ),
    .A2(net437),
    .B1(_06288_),
    .X(_01652_));
 sky130_fd_sc_hd__nand2_1 _11323_ (.A(net394),
    .B(_06241_),
    .Y(_06289_));
 sky130_fd_sc_hd__nand2_1 _11324_ (.A(_06047_),
    .B(_06050_),
    .Y(_06290_));
 sky130_fd_sc_hd__mux2_2 _11325_ (.A0(_06280_),
    .A1(_06290_),
    .S(net383),
    .X(_06291_));
 sky130_fd_sc_hd__o221a_1 _11326_ (.A1(_06089_),
    .A2(_06265_),
    .B1(_06291_),
    .B2(_04499_),
    .C1(_06289_),
    .X(_06292_));
 sky130_fd_sc_hd__or2_1 _11327_ (.A(_04482_),
    .B(_06292_),
    .X(_06293_));
 sky130_fd_sc_hd__o221a_1 _11328_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_sll[27] ),
    .A2(net437),
    .B1(_04587_),
    .B2(_06271_),
    .C1(_06293_),
    .X(_01653_));
 sky130_fd_sc_hd__nor2_1 _11329_ (.A(net397),
    .B(_06247_),
    .Y(_06294_));
 sky130_fd_sc_hd__nand2_1 _11330_ (.A(net378),
    .B(_06284_),
    .Y(_06295_));
 sky130_fd_sc_hd__o21ai_2 _11331_ (.A1(net376),
    .A2(net360),
    .B1(_06004_),
    .Y(_06296_));
 sky130_fd_sc_hd__o211a_1 _11332_ (.A1(net378),
    .A2(_06296_),
    .B1(_06295_),
    .C1(_04498_),
    .X(_06297_));
 sky130_fd_sc_hd__a211o_1 _11333_ (.A1(_06088_),
    .A2(_06275_),
    .B1(_06297_),
    .C1(net389),
    .X(_06298_));
 sky130_fd_sc_hd__o221a_1 _11334_ (.A1(net392),
    .A2(_04596_),
    .B1(_06294_),
    .B2(_06298_),
    .C1(net438),
    .X(_06299_));
 sky130_fd_sc_hd__a21o_1 _11335_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_sll[28] ),
    .A2(net436),
    .B1(_06299_),
    .X(_01654_));
 sky130_fd_sc_hd__a21oi_1 _11336_ (.A1(_06046_),
    .A2(_06054_),
    .B1(_04488_),
    .Y(_06300_));
 sky130_fd_sc_hd__a211o_1 _11337_ (.A1(_04488_),
    .A2(_06290_),
    .B1(_06300_),
    .C1(_04499_),
    .X(_06301_));
 sky130_fd_sc_hd__o211a_1 _11338_ (.A1(_06089_),
    .A2(_06281_),
    .B1(_06301_),
    .C1(net280),
    .X(_06302_));
 sky130_fd_sc_hd__o21a_1 _11339_ (.A1(net396),
    .A2(_06254_),
    .B1(_06302_),
    .X(_06303_));
 sky130_fd_sc_hd__a221o_1 _11340_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_sll[29] ),
    .A2(net435),
    .B1(_04605_),
    .B2(_06272_),
    .C1(_06303_),
    .X(_01655_));
 sky130_fd_sc_hd__o211ai_4 _11341_ (.A1(net373),
    .A2(_05688_),
    .B1(_06003_),
    .C1(net382),
    .Y(_06304_));
 sky130_fd_sc_hd__o211a_1 _11342_ (.A1(net382),
    .A2(_06296_),
    .B1(_06304_),
    .C1(_04498_),
    .X(_06305_));
 sky130_fd_sc_hd__o22a_1 _11343_ (.A1(net397),
    .A2(_06260_),
    .B1(_06285_),
    .B2(_06089_),
    .X(_06306_));
 sky130_fd_sc_hd__or3b_1 _11344_ (.A(net389),
    .B(_06305_),
    .C_N(_06306_),
    .X(_06307_));
 sky130_fd_sc_hd__o211a_1 _11345_ (.A1(net392),
    .A2(_04614_),
    .B1(_06307_),
    .C1(net438),
    .X(_06308_));
 sky130_fd_sc_hd__a21o_1 _11346_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_sll[30] ),
    .A2(net436),
    .B1(_06308_),
    .X(_01656_));
 sky130_fd_sc_hd__nand2_1 _11347_ (.A(net394),
    .B(_06267_),
    .Y(_06309_));
 sky130_fd_sc_hd__a21oi_1 _11348_ (.A1(_06046_),
    .A2(_06054_),
    .B1(net382),
    .Y(_06310_));
 sky130_fd_sc_hd__and3_1 _11349_ (.A(net383),
    .B(net374),
    .C(_05687_),
    .X(_06311_));
 sky130_fd_sc_hd__a211o_1 _11350_ (.A1(_04492_),
    .A2(_05614_),
    .B1(_06311_),
    .C1(_04499_),
    .X(_06312_));
 sky130_fd_sc_hd__o221a_1 _11351_ (.A1(_06089_),
    .A2(_06291_),
    .B1(_06310_),
    .B2(_06312_),
    .C1(net280),
    .X(_06313_));
 sky130_fd_sc_hd__a22oi_1 _11352_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_sll[31] ),
    .A2(net435),
    .B1(_06309_),
    .B2(_06313_),
    .Y(_06314_));
 sky130_fd_sc_hd__o21ai_1 _11353_ (.A1(_04622_),
    .A2(_06271_),
    .B1(_06314_),
    .Y(_01657_));
 sky130_fd_sc_hd__or3_2 _11354_ (.A(\core_pipeline.decode_to_execute_alu_function[2] ),
    .B(\core_pipeline.decode_to_execute_alu_function[1] ),
    .C(\core_pipeline.decode_to_execute_alu_function[0] ),
    .X(_06315_));
 sky130_fd_sc_hd__mux2_1 _11355_ (.A0(_05816_),
    .A1(net493),
    .S(net409),
    .X(_01658_));
 sky130_fd_sc_hd__or3_1 _11356_ (.A(net631),
    .B(net379),
    .C(net377),
    .X(_06316_));
 sky130_fd_sc_hd__and3_1 _11357_ (.A(_04502_),
    .B(_06053_),
    .C(_06316_),
    .X(_06317_));
 sky130_fd_sc_hd__a21oi_1 _11358_ (.A1(_06053_),
    .A2(_06316_),
    .B1(_04502_),
    .Y(_06318_));
 sky130_fd_sc_hd__nor2_1 _11359_ (.A(_06317_),
    .B(_06318_),
    .Y(_06319_));
 sky130_fd_sc_hd__xnor2_1 _11360_ (.A(_04503_),
    .B(_06319_),
    .Y(_06320_));
 sky130_fd_sc_hd__mux2_1 _11361_ (.A0(_06320_),
    .A1(net492),
    .S(net409),
    .X(_01659_));
 sky130_fd_sc_hd__or3_1 _11362_ (.A(net631),
    .B(net384),
    .C(_04492_),
    .X(_06321_));
 sky130_fd_sc_hd__and3b_1 _11363_ (.A_N(_04511_),
    .B(_06117_),
    .C(_06321_),
    .X(_06322_));
 sky130_fd_sc_hd__a21bo_1 _11364_ (.A1(_06117_),
    .A2(_06321_),
    .B1_N(_04511_),
    .X(_06323_));
 sky130_fd_sc_hd__and2b_1 _11365_ (.A_N(_06322_),
    .B(_06323_),
    .X(_06324_));
 sky130_fd_sc_hd__a21o_1 _11366_ (.A1(_04504_),
    .A2(_06319_),
    .B1(_06317_),
    .X(_06325_));
 sky130_fd_sc_hd__nor2_1 _11367_ (.A(_06324_),
    .B(_06325_),
    .Y(_06326_));
 sky130_fd_sc_hd__and2_1 _11368_ (.A(_06324_),
    .B(_06325_),
    .X(_06327_));
 sky130_fd_sc_hd__or3_1 _11369_ (.A(net409),
    .B(_06326_),
    .C(_06327_),
    .X(_06328_));
 sky130_fd_sc_hd__a21bo_1 _11370_ (.A1(\core_busio.mem_address[2] ),
    .A2(net409),
    .B1_N(_06328_),
    .X(_01660_));
 sky130_fd_sc_hd__or2_1 _11371_ (.A(net395),
    .B(_06155_),
    .X(_06329_));
 sky130_fd_sc_hd__a21bo_2 _11372_ (.A1(_06156_),
    .A2(_06329_),
    .B1_N(_04517_),
    .X(_06330_));
 sky130_fd_sc_hd__inv_2 _11373_ (.A(_06330_),
    .Y(_06331_));
 sky130_fd_sc_hd__a21oi_1 _11374_ (.A1(_06323_),
    .A2(_06325_),
    .B1(_06322_),
    .Y(_06332_));
 sky130_fd_sc_hd__and3b_1 _11375_ (.A_N(_04517_),
    .B(_06156_),
    .C(_06329_),
    .X(_06333_));
 sky130_fd_sc_hd__a211o_1 _11376_ (.A1(_06324_),
    .A2(_06325_),
    .B1(_06333_),
    .C1(_06322_),
    .X(_06334_));
 sky130_fd_sc_hd__nor2_1 _11377_ (.A(_06331_),
    .B(_06333_),
    .Y(_06335_));
 sky130_fd_sc_hd__xnor2_1 _11378_ (.A(_06332_),
    .B(_06335_),
    .Y(_06336_));
 sky130_fd_sc_hd__mux2_1 _11379_ (.A0(_06336_),
    .A1(\core_busio.mem_address[3] ),
    .S(net409),
    .X(_01661_));
 sky130_fd_sc_hd__xnor2_2 _11380_ (.A(net391),
    .B(_06193_),
    .Y(_06337_));
 sky130_fd_sc_hd__nor2_2 _11381_ (.A(_04523_),
    .B(_06337_),
    .Y(_06338_));
 sky130_fd_sc_hd__inv_2 _11382_ (.A(_06338_),
    .Y(_06339_));
 sky130_fd_sc_hd__and2_1 _11383_ (.A(_04523_),
    .B(_06337_),
    .X(_06340_));
 sky130_fd_sc_hd__nor2_1 _11384_ (.A(_06338_),
    .B(_06340_),
    .Y(_06341_));
 sky130_fd_sc_hd__and2_1 _11385_ (.A(_06330_),
    .B(_06334_),
    .X(_06342_));
 sky130_fd_sc_hd__xor2_1 _11386_ (.A(_06341_),
    .B(_06342_),
    .X(_06343_));
 sky130_fd_sc_hd__mux2_1 _11387_ (.A0(_06343_),
    .A1(\core_busio.mem_address[4] ),
    .S(net409),
    .X(_01662_));
 sky130_fd_sc_hd__a21bo_1 _11388_ (.A1(_06193_),
    .A2(_06212_),
    .B1_N(_05666_),
    .X(_06344_));
 sky130_fd_sc_hd__nand3b_2 _11389_ (.A_N(_05666_),
    .B(_06193_),
    .C(_06212_),
    .Y(_06345_));
 sky130_fd_sc_hd__nand3_2 _11390_ (.A(_04530_),
    .B(_06344_),
    .C(_06345_),
    .Y(_06346_));
 sky130_fd_sc_hd__a21o_1 _11391_ (.A1(_06344_),
    .A2(_06345_),
    .B1(_04530_),
    .X(_06347_));
 sky130_fd_sc_hd__nand2_1 _11392_ (.A(_06346_),
    .B(_06347_),
    .Y(_06348_));
 sky130_fd_sc_hd__a31o_1 _11393_ (.A1(_06330_),
    .A2(_06334_),
    .A3(_06341_),
    .B1(_06338_),
    .X(_06349_));
 sky130_fd_sc_hd__xnor2_1 _11394_ (.A(_06348_),
    .B(_06349_),
    .Y(_06350_));
 sky130_fd_sc_hd__mux2_1 _11395_ (.A0(_06350_),
    .A1(\core_busio.mem_address[5] ),
    .S(net409),
    .X(_01663_));
 sky130_fd_sc_hd__a31o_1 _11396_ (.A1(net393),
    .A2(_04500_),
    .A3(_05666_),
    .B1(net632),
    .X(_06351_));
 sky130_fd_sc_hd__xnor2_1 _11397_ (.A(_05662_),
    .B(_06351_),
    .Y(_06352_));
 sky130_fd_sc_hd__and2_1 _11398_ (.A(_04538_),
    .B(_06352_),
    .X(_06353_));
 sky130_fd_sc_hd__nor2_1 _11399_ (.A(_04538_),
    .B(_06352_),
    .Y(_06354_));
 sky130_fd_sc_hd__nor2_2 _11400_ (.A(_06353_),
    .B(_06354_),
    .Y(_06355_));
 sky130_fd_sc_hd__and3_1 _11401_ (.A(_06341_),
    .B(_06346_),
    .C(_06347_),
    .X(_06356_));
 sky130_fd_sc_hd__a21boi_2 _11402_ (.A1(_06339_),
    .A2(_06346_),
    .B1_N(_06347_),
    .Y(_06357_));
 sky130_fd_sc_hd__a21oi_2 _11403_ (.A1(_06342_),
    .A2(_06356_),
    .B1(_06357_),
    .Y(_06358_));
 sky130_fd_sc_hd__xnor2_1 _11404_ (.A(_06355_),
    .B(_06358_),
    .Y(_06359_));
 sky130_fd_sc_hd__mux2_1 _11405_ (.A0(_06359_),
    .A1(\core_busio.mem_address[6] ),
    .S(net409),
    .X(_01664_));
 sky130_fd_sc_hd__a41o_1 _11406_ (.A1(net393),
    .A2(_04500_),
    .A3(_05662_),
    .A4(_05666_),
    .B1(net631),
    .X(_06360_));
 sky130_fd_sc_hd__xor2_1 _11407_ (.A(_05657_),
    .B(_06360_),
    .X(_06361_));
 sky130_fd_sc_hd__nor2_1 _11408_ (.A(_04545_),
    .B(_06361_),
    .Y(_06362_));
 sky130_fd_sc_hd__nand2_1 _11409_ (.A(_04545_),
    .B(_06361_),
    .Y(_06363_));
 sky130_fd_sc_hd__and2b_1 _11410_ (.A_N(_06362_),
    .B(_06363_),
    .X(_06364_));
 sky130_fd_sc_hd__o21ba_1 _11411_ (.A1(_06354_),
    .A2(_06358_),
    .B1_N(_06353_),
    .X(_06365_));
 sky130_fd_sc_hd__xnor2_1 _11412_ (.A(_06364_),
    .B(_06365_),
    .Y(_06366_));
 sky130_fd_sc_hd__mux2_1 _11413_ (.A0(_06366_),
    .A1(\core_busio.mem_address[7] ),
    .S(net409),
    .X(_01665_));
 sky130_fd_sc_hd__and4_4 _11414_ (.A(net393),
    .B(_05657_),
    .C(_05662_),
    .D(_05666_),
    .X(_06367_));
 sky130_fd_sc_hd__a21oi_1 _11415_ (.A1(_04500_),
    .A2(_06367_),
    .B1(net635),
    .Y(_06368_));
 sky130_fd_sc_hd__xnor2_1 _11416_ (.A(_05633_),
    .B(_06368_),
    .Y(_06369_));
 sky130_fd_sc_hd__or2_1 _11417_ (.A(_04553_),
    .B(_06369_),
    .X(_06370_));
 sky130_fd_sc_hd__and2_1 _11418_ (.A(_04553_),
    .B(_06369_),
    .X(_06371_));
 sky130_fd_sc_hd__nand2_1 _11419_ (.A(_04553_),
    .B(_06369_),
    .Y(_06372_));
 sky130_fd_sc_hd__and2_1 _11420_ (.A(_06370_),
    .B(_06372_),
    .X(_06373_));
 sky130_fd_sc_hd__or2_1 _11421_ (.A(_06353_),
    .B(_06362_),
    .X(_06374_));
 sky130_fd_sc_hd__a32o_2 _11422_ (.A1(_06355_),
    .A2(_06357_),
    .A3(_06364_),
    .B1(_06374_),
    .B2(_06363_),
    .X(_06375_));
 sky130_fd_sc_hd__and4_2 _11423_ (.A(_06330_),
    .B(_06334_),
    .C(_06356_),
    .D(_06364_),
    .X(_06376_));
 sky130_fd_sc_hd__a21oi_4 _11424_ (.A1(_06355_),
    .A2(_06376_),
    .B1(_06375_),
    .Y(_06377_));
 sky130_fd_sc_hd__xnor2_1 _11425_ (.A(_06373_),
    .B(_06377_),
    .Y(_06378_));
 sky130_fd_sc_hd__mux2_1 _11426_ (.A0(_06378_),
    .A1(\core_busio.mem_address[8] ),
    .S(net408),
    .X(_01666_));
 sky130_fd_sc_hd__a31o_1 _11427_ (.A1(_04500_),
    .A2(_05633_),
    .A3(_06367_),
    .B1(net635),
    .X(_06379_));
 sky130_fd_sc_hd__xor2_2 _11428_ (.A(_05636_),
    .B(_06379_),
    .X(_06380_));
 sky130_fd_sc_hd__nor2_1 _11429_ (.A(_04565_),
    .B(_06380_),
    .Y(_06381_));
 sky130_fd_sc_hd__or2_1 _11430_ (.A(_04565_),
    .B(_06380_),
    .X(_06382_));
 sky130_fd_sc_hd__and2_1 _11431_ (.A(_04565_),
    .B(_06380_),
    .X(_06383_));
 sky130_fd_sc_hd__nor2_1 _11432_ (.A(_06381_),
    .B(_06383_),
    .Y(_06384_));
 sky130_fd_sc_hd__o21a_1 _11433_ (.A1(_06371_),
    .A2(_06377_),
    .B1(_06370_),
    .X(_06385_));
 sky130_fd_sc_hd__xnor2_1 _11434_ (.A(_06384_),
    .B(_06385_),
    .Y(_06386_));
 sky130_fd_sc_hd__mux2_1 _11435_ (.A0(_06386_),
    .A1(\core_busio.mem_address[9] ),
    .S(net408),
    .X(_01667_));
 sky130_fd_sc_hd__and2_1 _11436_ (.A(_05633_),
    .B(_05636_),
    .X(_06387_));
 sky130_fd_sc_hd__and3_2 _11437_ (.A(_04500_),
    .B(_06367_),
    .C(_06387_),
    .X(_06388_));
 sky130_fd_sc_hd__or2_4 _11438_ (.A(net635),
    .B(_06388_),
    .X(_06389_));
 sky130_fd_sc_hd__xnor2_4 _11439_ (.A(_05651_),
    .B(_06389_),
    .Y(_06390_));
 sky130_fd_sc_hd__xnor2_2 _11440_ (.A(_04574_),
    .B(_06390_),
    .Y(_06391_));
 sky130_fd_sc_hd__or2_1 _11441_ (.A(_06383_),
    .B(_06385_),
    .X(_06392_));
 sky130_fd_sc_hd__a21oi_1 _11442_ (.A1(_06370_),
    .A2(_06382_),
    .B1(_06383_),
    .Y(_06393_));
 sky130_fd_sc_hd__a21oi_1 _11443_ (.A1(_06382_),
    .A2(_06392_),
    .B1(_06391_),
    .Y(_06394_));
 sky130_fd_sc_hd__a31o_1 _11444_ (.A1(_06382_),
    .A2(_06391_),
    .A3(_06392_),
    .B1(net408),
    .X(_06395_));
 sky130_fd_sc_hd__a2bb2o_1 _11445_ (.A1_N(_06394_),
    .A2_N(_06395_),
    .B1(\core_busio.mem_address[10] ),
    .B2(net408),
    .X(_01668_));
 sky130_fd_sc_hd__a21oi_1 _11446_ (.A1(_05651_),
    .A2(_06388_),
    .B1(net635),
    .Y(_06396_));
 sky130_fd_sc_hd__xnor2_1 _11447_ (.A(_05639_),
    .B(_06396_),
    .Y(_06397_));
 sky130_fd_sc_hd__nand2_1 _11448_ (.A(_04581_),
    .B(_06397_),
    .Y(_06398_));
 sky130_fd_sc_hd__or2_1 _11449_ (.A(_04581_),
    .B(_06397_),
    .X(_06399_));
 sky130_fd_sc_hd__and2_1 _11450_ (.A(_06398_),
    .B(_06399_),
    .X(_06400_));
 sky130_fd_sc_hd__a21oi_1 _11451_ (.A1(_04574_),
    .A2(_06390_),
    .B1(_06394_),
    .Y(_06401_));
 sky130_fd_sc_hd__xnor2_1 _11452_ (.A(_06400_),
    .B(_06401_),
    .Y(_06402_));
 sky130_fd_sc_hd__mux2_1 _11453_ (.A0(_06402_),
    .A1(\core_busio.mem_address[11] ),
    .S(net408),
    .X(_01669_));
 sky130_fd_sc_hd__a31o_1 _11454_ (.A1(_05639_),
    .A2(_05651_),
    .A3(_06388_),
    .B1(net635),
    .X(_06403_));
 sky130_fd_sc_hd__xnor2_1 _11455_ (.A(_05642_),
    .B(_06403_),
    .Y(_06404_));
 sky130_fd_sc_hd__nor2_1 _11456_ (.A(net371),
    .B(_06404_),
    .Y(_06405_));
 sky130_fd_sc_hd__and2_1 _11457_ (.A(net371),
    .B(_06404_),
    .X(_06406_));
 sky130_fd_sc_hd__nor2_1 _11458_ (.A(_06405_),
    .B(_06406_),
    .Y(_06407_));
 sky130_fd_sc_hd__and2b_1 _11459_ (.A_N(_06391_),
    .B(_06400_),
    .X(_06408_));
 sky130_fd_sc_hd__and4b_2 _11460_ (.A_N(_06377_),
    .B(_06384_),
    .C(_06408_),
    .D(_06373_),
    .X(_06409_));
 sky130_fd_sc_hd__a21bo_1 _11461_ (.A1(_04574_),
    .A2(_06390_),
    .B1_N(_06399_),
    .X(_06410_));
 sky130_fd_sc_hd__a22o_1 _11462_ (.A1(_06393_),
    .A2(_06408_),
    .B1(_06410_),
    .B2(_06398_),
    .X(_06411_));
 sky130_fd_sc_hd__o21a_1 _11463_ (.A1(_06409_),
    .A2(_06411_),
    .B1(_06407_),
    .X(_06412_));
 sky130_fd_sc_hd__nor3_1 _11464_ (.A(_06407_),
    .B(_06409_),
    .C(_06411_),
    .Y(_06413_));
 sky130_fd_sc_hd__or3_1 _11465_ (.A(net408),
    .B(_06412_),
    .C(_06413_),
    .X(_06414_));
 sky130_fd_sc_hd__a21bo_1 _11466_ (.A1(\core_busio.mem_address[12] ),
    .A2(net408),
    .B1_N(_06414_),
    .X(_01670_));
 sky130_fd_sc_hd__a21boi_1 _11467_ (.A1(_03423_),
    .A2(_05642_),
    .B1_N(_06403_),
    .Y(_06415_));
 sky130_fd_sc_hd__xnor2_1 _11468_ (.A(_05623_),
    .B(_06415_),
    .Y(_06416_));
 sky130_fd_sc_hd__nor2_1 _11469_ (.A(_04599_),
    .B(_06416_),
    .Y(_06417_));
 sky130_fd_sc_hd__and2_1 _11470_ (.A(_04599_),
    .B(_06416_),
    .X(_06418_));
 sky130_fd_sc_hd__nor2_1 _11471_ (.A(_06417_),
    .B(_06418_),
    .Y(_06419_));
 sky130_fd_sc_hd__nor2_1 _11472_ (.A(_06405_),
    .B(_06412_),
    .Y(_06420_));
 sky130_fd_sc_hd__xnor2_1 _11473_ (.A(_06419_),
    .B(_06420_),
    .Y(_06421_));
 sky130_fd_sc_hd__mux2_1 _11474_ (.A0(_06421_),
    .A1(\core_busio.mem_address[13] ),
    .S(net408),
    .X(_01671_));
 sky130_fd_sc_hd__nor2_1 _11475_ (.A(_05623_),
    .B(_05642_),
    .Y(_06422_));
 sky130_fd_sc_hd__and4_1 _11476_ (.A(_05639_),
    .B(_05651_),
    .C(_06388_),
    .D(_06422_),
    .X(_06423_));
 sky130_fd_sc_hd__or2_2 _11477_ (.A(net634),
    .B(_06423_),
    .X(_06424_));
 sky130_fd_sc_hd__xor2_2 _11478_ (.A(_05618_),
    .B(_06424_),
    .X(_06425_));
 sky130_fd_sc_hd__nor2_2 _11479_ (.A(_04608_),
    .B(_06425_),
    .Y(_06426_));
 sky130_fd_sc_hd__and2_1 _11480_ (.A(_04608_),
    .B(_06425_),
    .X(_06427_));
 sky130_fd_sc_hd__nor2_2 _11481_ (.A(_06426_),
    .B(_06427_),
    .Y(_06428_));
 sky130_fd_sc_hd__o21ba_1 _11482_ (.A1(_06405_),
    .A2(_06417_),
    .B1_N(_06418_),
    .X(_06429_));
 sky130_fd_sc_hd__a21o_1 _11483_ (.A1(_06412_),
    .A2(_06419_),
    .B1(_06429_),
    .X(_06430_));
 sky130_fd_sc_hd__nand2_1 _11484_ (.A(_06428_),
    .B(_06430_),
    .Y(_06431_));
 sky130_fd_sc_hd__o21ba_1 _11485_ (.A1(_06428_),
    .A2(_06430_),
    .B1_N(net408),
    .X(_06432_));
 sky130_fd_sc_hd__a22o_1 _11486_ (.A1(\core_busio.mem_address[14] ),
    .A2(net407),
    .B1(_06431_),
    .B2(_06432_),
    .X(_01672_));
 sky130_fd_sc_hd__a211o_1 _11487_ (.A1(_05618_),
    .A2(_06423_),
    .B1(_05627_),
    .C1(net634),
    .X(_06433_));
 sky130_fd_sc_hd__o211ai_2 _11488_ (.A1(net634),
    .A2(_05618_),
    .B1(_05627_),
    .C1(_06424_),
    .Y(_06434_));
 sky130_fd_sc_hd__a21oi_1 _11489_ (.A1(_06433_),
    .A2(_06434_),
    .B1(_04618_),
    .Y(_06435_));
 sky130_fd_sc_hd__a21o_1 _11490_ (.A1(_06428_),
    .A2(_06430_),
    .B1(_06426_),
    .X(_06436_));
 sky130_fd_sc_hd__and3_1 _11491_ (.A(_04618_),
    .B(_06433_),
    .C(_06434_),
    .X(_06437_));
 sky130_fd_sc_hd__nor2_1 _11492_ (.A(_06435_),
    .B(_06437_),
    .Y(_06438_));
 sky130_fd_sc_hd__nand2_1 _11493_ (.A(_06436_),
    .B(_06438_),
    .Y(_06439_));
 sky130_fd_sc_hd__o21ba_1 _11494_ (.A1(_06436_),
    .A2(_06438_),
    .B1_N(net408),
    .X(_06440_));
 sky130_fd_sc_hd__a22o_1 _11495_ (.A1(\core_busio.mem_address[15] ),
    .A2(net408),
    .B1(_06439_),
    .B2(_06440_),
    .X(_01673_));
 sky130_fd_sc_hd__and3_2 _11496_ (.A(_05618_),
    .B(_05626_),
    .C(_06423_),
    .X(_06441_));
 sky130_fd_sc_hd__or2_1 _11497_ (.A(net633),
    .B(_06441_),
    .X(_06442_));
 sky130_fd_sc_hd__xnor2_1 _11498_ (.A(_05758_),
    .B(_06442_),
    .Y(_06443_));
 sky130_fd_sc_hd__nand2_1 _11499_ (.A(_05760_),
    .B(_06443_),
    .Y(_06444_));
 sky130_fd_sc_hd__or2_1 _11500_ (.A(_05760_),
    .B(_06443_),
    .X(_06445_));
 sky130_fd_sc_hd__and2_2 _11501_ (.A(_06444_),
    .B(_06445_),
    .X(_06446_));
 sky130_fd_sc_hd__nor2_1 _11502_ (.A(_06426_),
    .B(_06437_),
    .Y(_06447_));
 sky130_fd_sc_hd__and2_1 _11503_ (.A(_06428_),
    .B(_06438_),
    .X(_06448_));
 sky130_fd_sc_hd__a2bb2o_1 _11504_ (.A1_N(_06435_),
    .A2_N(_06447_),
    .B1(_06448_),
    .B2(_06429_),
    .X(_06449_));
 sky130_fd_sc_hd__and4_1 _11505_ (.A(_06407_),
    .B(_06419_),
    .C(_06428_),
    .D(_06438_),
    .X(_06450_));
 sky130_fd_sc_hd__o21a_1 _11506_ (.A1(_06409_),
    .A2(_06411_),
    .B1(_06450_),
    .X(_06451_));
 sky130_fd_sc_hd__or2_4 _11507_ (.A(_06449_),
    .B(_06451_),
    .X(_06452_));
 sky130_fd_sc_hd__xor2_1 _11508_ (.A(_06446_),
    .B(_06452_),
    .X(_06453_));
 sky130_fd_sc_hd__mux2_1 _11509_ (.A0(_06453_),
    .A1(\core_busio.mem_address[16] ),
    .S(net407),
    .X(_01674_));
 sky130_fd_sc_hd__a21o_1 _11510_ (.A1(_05758_),
    .A2(_06441_),
    .B1(net634),
    .X(_06454_));
 sky130_fd_sc_hd__xor2_1 _11511_ (.A(_05745_),
    .B(_06454_),
    .X(_06455_));
 sky130_fd_sc_hd__and2b_1 _11512_ (.A_N(_05748_),
    .B(_06455_),
    .X(_06456_));
 sky130_fd_sc_hd__a21bo_1 _11513_ (.A1(_06446_),
    .A2(_06452_),
    .B1_N(_06444_),
    .X(_06457_));
 sky130_fd_sc_hd__o21bai_1 _11514_ (.A1(_05746_),
    .A2(_05747_),
    .B1_N(_06455_),
    .Y(_06458_));
 sky130_fd_sc_hd__and2b_1 _11515_ (.A_N(_06456_),
    .B(_06458_),
    .X(_06459_));
 sky130_fd_sc_hd__xor2_1 _11516_ (.A(_06457_),
    .B(_06459_),
    .X(_06460_));
 sky130_fd_sc_hd__mux2_1 _11517_ (.A0(_06460_),
    .A1(\core_busio.mem_address[17] ),
    .S(net407),
    .X(_01675_));
 sky130_fd_sc_hd__a31o_1 _11518_ (.A1(_05745_),
    .A2(_05758_),
    .A3(_06441_),
    .B1(net633),
    .X(_06461_));
 sky130_fd_sc_hd__xnor2_1 _11519_ (.A(_05779_),
    .B(_06461_),
    .Y(_06462_));
 sky130_fd_sc_hd__nand2_1 _11520_ (.A(_05781_),
    .B(_06462_),
    .Y(_06463_));
 sky130_fd_sc_hd__or2_1 _11521_ (.A(_05781_),
    .B(_06462_),
    .X(_06464_));
 sky130_fd_sc_hd__nand2_1 _11522_ (.A(_06463_),
    .B(_06464_),
    .Y(_06465_));
 sky130_fd_sc_hd__a21oi_1 _11523_ (.A1(_06444_),
    .A2(_06458_),
    .B1(_06456_),
    .Y(_06466_));
 sky130_fd_sc_hd__a31o_1 _11524_ (.A1(_06446_),
    .A2(_06452_),
    .A3(_06459_),
    .B1(_06466_),
    .X(_06467_));
 sky130_fd_sc_hd__nand2b_1 _11525_ (.A_N(_06465_),
    .B(_06467_),
    .Y(_06468_));
 sky130_fd_sc_hd__xnor2_1 _11526_ (.A(_06465_),
    .B(_06467_),
    .Y(_06469_));
 sky130_fd_sc_hd__mux2_1 _11527_ (.A0(_06469_),
    .A1(\core_busio.mem_address[18] ),
    .S(net407),
    .X(_01676_));
 sky130_fd_sc_hd__a41o_1 _11528_ (.A1(_05745_),
    .A2(_05758_),
    .A3(_05779_),
    .A4(_06441_),
    .B1(net633),
    .X(_06470_));
 sky130_fd_sc_hd__xor2_1 _11529_ (.A(_05786_),
    .B(_06470_),
    .X(_06471_));
 sky130_fd_sc_hd__and2_1 _11530_ (.A(_05788_),
    .B(_06471_),
    .X(_06472_));
 sky130_fd_sc_hd__nand2_1 _11531_ (.A(_06463_),
    .B(_06468_),
    .Y(_06473_));
 sky130_fd_sc_hd__or2_1 _11532_ (.A(_05788_),
    .B(_06471_),
    .X(_06474_));
 sky130_fd_sc_hd__nand2b_1 _11533_ (.A_N(_06472_),
    .B(_06474_),
    .Y(_06475_));
 sky130_fd_sc_hd__xnor2_1 _11534_ (.A(_06473_),
    .B(_06475_),
    .Y(_06476_));
 sky130_fd_sc_hd__mux2_1 _11535_ (.A0(_06476_),
    .A1(\core_busio.mem_address[19] ),
    .S(net407),
    .X(_01677_));
 sky130_fd_sc_hd__and4_1 _11536_ (.A(_05745_),
    .B(_05758_),
    .C(_05779_),
    .D(_05786_),
    .X(_06477_));
 sky130_fd_sc_hd__and2_1 _11537_ (.A(_06441_),
    .B(_06477_),
    .X(_06478_));
 sky130_fd_sc_hd__nor2_1 _11538_ (.A(net633),
    .B(_06478_),
    .Y(_06479_));
 sky130_fd_sc_hd__xnor2_1 _11539_ (.A(_05771_),
    .B(_06479_),
    .Y(_06480_));
 sky130_fd_sc_hd__or2_2 _11540_ (.A(_05773_),
    .B(_06480_),
    .X(_06481_));
 sky130_fd_sc_hd__nand2_1 _11541_ (.A(_05773_),
    .B(_06480_),
    .Y(_06482_));
 sky130_fd_sc_hd__nand2_1 _11542_ (.A(_06481_),
    .B(_06482_),
    .Y(_06483_));
 sky130_fd_sc_hd__a21oi_1 _11543_ (.A1(_06463_),
    .A2(_06474_),
    .B1(_06472_),
    .Y(_06484_));
 sky130_fd_sc_hd__nor2_1 _11544_ (.A(_06465_),
    .B(_06475_),
    .Y(_06485_));
 sky130_fd_sc_hd__a21o_1 _11545_ (.A1(_06466_),
    .A2(_06485_),
    .B1(_06484_),
    .X(_06486_));
 sky130_fd_sc_hd__and3_1 _11546_ (.A(_06446_),
    .B(_06459_),
    .C(_06485_),
    .X(_06487_));
 sky130_fd_sc_hd__a21o_2 _11547_ (.A1(_06452_),
    .A2(_06487_),
    .B1(_06486_),
    .X(_06488_));
 sky130_fd_sc_hd__nand2b_1 _11548_ (.A_N(_06483_),
    .B(_06488_),
    .Y(_06489_));
 sky130_fd_sc_hd__xnor2_1 _11549_ (.A(_06483_),
    .B(_06488_),
    .Y(_06490_));
 sky130_fd_sc_hd__mux2_1 _11550_ (.A0(_06490_),
    .A1(\core_busio.mem_address[20] ),
    .S(net407),
    .X(_01678_));
 sky130_fd_sc_hd__a31o_1 _11551_ (.A1(_05771_),
    .A2(_06441_),
    .A3(_06477_),
    .B1(net633),
    .X(_06491_));
 sky130_fd_sc_hd__xor2_2 _11552_ (.A(_05763_),
    .B(_06491_),
    .X(_06492_));
 sky130_fd_sc_hd__or2_1 _11553_ (.A(_05766_),
    .B(_06492_),
    .X(_06493_));
 sky130_fd_sc_hd__and2_1 _11554_ (.A(_05766_),
    .B(_06492_),
    .X(_06494_));
 sky130_fd_sc_hd__nand2_1 _11555_ (.A(_05766_),
    .B(_06492_),
    .Y(_06495_));
 sky130_fd_sc_hd__nand2_1 _11556_ (.A(_06493_),
    .B(_06495_),
    .Y(_06496_));
 sky130_fd_sc_hd__a21oi_1 _11557_ (.A1(_06481_),
    .A2(_06489_),
    .B1(_06496_),
    .Y(_06497_));
 sky130_fd_sc_hd__a31o_1 _11558_ (.A1(_06481_),
    .A2(_06489_),
    .A3(_06496_),
    .B1(net407),
    .X(_06498_));
 sky130_fd_sc_hd__a2bb2o_1 _11559_ (.A1_N(_06497_),
    .A2_N(_06498_),
    .B1(\core_busio.mem_address[21] ),
    .B2(net407),
    .X(_01679_));
 sky130_fd_sc_hd__a31o_1 _11560_ (.A1(_05763_),
    .A2(_05771_),
    .A3(_06478_),
    .B1(net633),
    .X(_06499_));
 sky130_fd_sc_hd__xor2_2 _11561_ (.A(_05751_),
    .B(_06499_),
    .X(_06500_));
 sky130_fd_sc_hd__nand2_2 _11562_ (.A(_05753_),
    .B(_06500_),
    .Y(_06501_));
 sky130_fd_sc_hd__or2_1 _11563_ (.A(_05753_),
    .B(_06500_),
    .X(_06502_));
 sky130_fd_sc_hd__nand2_2 _11564_ (.A(_06501_),
    .B(_06502_),
    .Y(_06503_));
 sky130_fd_sc_hd__a31o_1 _11565_ (.A1(_06481_),
    .A2(_06489_),
    .A3(_06493_),
    .B1(_06494_),
    .X(_06504_));
 sky130_fd_sc_hd__or2_1 _11566_ (.A(_06503_),
    .B(_06504_),
    .X(_06505_));
 sky130_fd_sc_hd__xor2_1 _11567_ (.A(_06503_),
    .B(_06504_),
    .X(_06506_));
 sky130_fd_sc_hd__mux2_1 _11568_ (.A0(_06506_),
    .A1(\core_busio.mem_address[22] ),
    .S(net407),
    .X(_01680_));
 sky130_fd_sc_hd__and4b_1 _11569_ (.A_N(_05751_),
    .B(_05763_),
    .C(_05771_),
    .D(_06478_),
    .X(_06507_));
 sky130_fd_sc_hd__or2_4 _11570_ (.A(net633),
    .B(_06507_),
    .X(_06508_));
 sky130_fd_sc_hd__xnor2_4 _11571_ (.A(_05738_),
    .B(_06508_),
    .Y(_06509_));
 sky130_fd_sc_hd__xnor2_4 _11572_ (.A(_05740_),
    .B(_06509_),
    .Y(_06510_));
 sky130_fd_sc_hd__a21oi_1 _11573_ (.A1(_06501_),
    .A2(_06505_),
    .B1(_06510_),
    .Y(_06511_));
 sky130_fd_sc_hd__a31o_1 _11574_ (.A1(_06501_),
    .A2(_06505_),
    .A3(_06510_),
    .B1(net407),
    .X(_06512_));
 sky130_fd_sc_hd__a2bb2o_1 _11575_ (.A1_N(_06511_),
    .A2_N(_06512_),
    .B1(\core_busio.mem_address[23] ),
    .B2(net407),
    .X(_01681_));
 sky130_fd_sc_hd__nor4_1 _11576_ (.A(_06483_),
    .B(_06496_),
    .C(_06503_),
    .D(_06510_),
    .Y(_06513_));
 sky130_fd_sc_hd__a21bo_1 _11577_ (.A1(_05740_),
    .A2(_06509_),
    .B1_N(_06501_),
    .X(_06514_));
 sky130_fd_sc_hd__o21a_1 _11578_ (.A1(_05740_),
    .A2(_06509_),
    .B1(_06514_),
    .X(_06515_));
 sky130_fd_sc_hd__a2111oi_1 _11579_ (.A1(_06481_),
    .A2(_06493_),
    .B1(_06494_),
    .C1(_06503_),
    .D1(_06510_),
    .Y(_06516_));
 sky130_fd_sc_hd__a211o_2 _11580_ (.A1(_06488_),
    .A2(_06513_),
    .B1(_06515_),
    .C1(_06516_),
    .X(_06517_));
 sky130_fd_sc_hd__a21o_1 _11581_ (.A1(_05738_),
    .A2(_06507_),
    .B1(net633),
    .X(_06518_));
 sky130_fd_sc_hd__xor2_1 _11582_ (.A(_05715_),
    .B(_06518_),
    .X(_06519_));
 sky130_fd_sc_hd__and2_1 _11583_ (.A(_05717_),
    .B(_06519_),
    .X(_06520_));
 sky130_fd_sc_hd__nor2_1 _11584_ (.A(_05717_),
    .B(_06519_),
    .Y(_06521_));
 sky130_fd_sc_hd__nor2_2 _11585_ (.A(_06520_),
    .B(_06521_),
    .Y(_06522_));
 sky130_fd_sc_hd__nand2_1 _11586_ (.A(_06517_),
    .B(_06522_),
    .Y(_06523_));
 sky130_fd_sc_hd__o21ba_1 _11587_ (.A1(_06517_),
    .A2(_06522_),
    .B1_N(net407),
    .X(_06524_));
 sky130_fd_sc_hd__a22o_1 _11588_ (.A1(\core_busio.mem_address[24] ),
    .A2(net407),
    .B1(_06523_),
    .B2(_06524_),
    .X(_01682_));
 sky130_fd_sc_hd__nand3b_1 _11589_ (.A_N(_05715_),
    .B(_05738_),
    .C(_06507_),
    .Y(_06525_));
 sky130_fd_sc_hd__and2_1 _11590_ (.A(net459),
    .B(_06525_),
    .X(_06526_));
 sky130_fd_sc_hd__xnor2_1 _11591_ (.A(_05729_),
    .B(_06526_),
    .Y(_06527_));
 sky130_fd_sc_hd__and2_1 _11592_ (.A(_05731_),
    .B(_06527_),
    .X(_06528_));
 sky130_fd_sc_hd__nor2_1 _11593_ (.A(_05731_),
    .B(_06527_),
    .Y(_06529_));
 sky130_fd_sc_hd__nor2_1 _11594_ (.A(_06528_),
    .B(_06529_),
    .Y(_06530_));
 sky130_fd_sc_hd__a21oi_2 _11595_ (.A1(_06517_),
    .A2(_06522_),
    .B1(_06520_),
    .Y(_06531_));
 sky130_fd_sc_hd__xnor2_1 _11596_ (.A(_06530_),
    .B(_06531_),
    .Y(_06532_));
 sky130_fd_sc_hd__mux2_1 _11597_ (.A0(_06532_),
    .A1(\core_busio.mem_address[25] ),
    .S(net407),
    .X(_01683_));
 sky130_fd_sc_hd__nor2_1 _11598_ (.A(_05729_),
    .B(_06525_),
    .Y(_06533_));
 sky130_fd_sc_hd__or2_1 _11599_ (.A(net633),
    .B(_06533_),
    .X(_06534_));
 sky130_fd_sc_hd__xnor2_1 _11600_ (.A(_05710_),
    .B(_06534_),
    .Y(_06535_));
 sky130_fd_sc_hd__and2_1 _11601_ (.A(_05712_),
    .B(_06535_),
    .X(_06536_));
 sky130_fd_sc_hd__nor2_1 _11602_ (.A(_05712_),
    .B(_06535_),
    .Y(_06537_));
 sky130_fd_sc_hd__nor2_1 _11603_ (.A(_06536_),
    .B(_06537_),
    .Y(_06538_));
 sky130_fd_sc_hd__nor2_1 _11604_ (.A(_06529_),
    .B(_06531_),
    .Y(_06539_));
 sky130_fd_sc_hd__o21a_1 _11605_ (.A1(_06528_),
    .A2(_06539_),
    .B1(_06538_),
    .X(_06540_));
 sky130_fd_sc_hd__or3_1 _11606_ (.A(_06528_),
    .B(_06538_),
    .C(_06539_),
    .X(_06541_));
 sky130_fd_sc_hd__or3b_1 _11607_ (.A(net407),
    .B(_06540_),
    .C_N(_06541_),
    .X(_06542_));
 sky130_fd_sc_hd__a21bo_1 _11608_ (.A1(\core_busio.mem_address[26] ),
    .A2(net407),
    .B1_N(_06542_),
    .X(_01684_));
 sky130_fd_sc_hd__a21o_2 _11609_ (.A1(_05710_),
    .A2(_06533_),
    .B1(net633),
    .X(_06543_));
 sky130_fd_sc_hd__xnor2_2 _11610_ (.A(_05722_),
    .B(_06543_),
    .Y(_06544_));
 sky130_fd_sc_hd__nor2_1 _11611_ (.A(_06536_),
    .B(_06540_),
    .Y(_06545_));
 sky130_fd_sc_hd__xor2_1 _11612_ (.A(net360),
    .B(_06544_),
    .X(_06546_));
 sky130_fd_sc_hd__xnor2_1 _11613_ (.A(_06545_),
    .B(_06546_),
    .Y(_06547_));
 sky130_fd_sc_hd__mux2_1 _11614_ (.A0(_06547_),
    .A1(\core_busio.mem_address[27] ),
    .S(net407),
    .X(_01685_));
 sky130_fd_sc_hd__a21boi_4 _11615_ (.A1(net459),
    .A2(_05722_),
    .B1_N(_06543_),
    .Y(_06548_));
 sky130_fd_sc_hd__xor2_4 _11616_ (.A(_05697_),
    .B(_06548_),
    .X(_06549_));
 sky130_fd_sc_hd__inv_2 _11617_ (.A(_06549_),
    .Y(_06550_));
 sky130_fd_sc_hd__xor2_2 _11618_ (.A(_05699_),
    .B(_06549_),
    .X(_06551_));
 sky130_fd_sc_hd__a2bb2o_1 _11619_ (.A1_N(_06536_),
    .A2_N(_06540_),
    .B1(_06544_),
    .B2(net360),
    .X(_06552_));
 sky130_fd_sc_hd__o21a_1 _11620_ (.A1(net360),
    .A2(_06544_),
    .B1(_06552_),
    .X(_06553_));
 sky130_fd_sc_hd__xor2_1 _11621_ (.A(_06551_),
    .B(_06553_),
    .X(_06554_));
 sky130_fd_sc_hd__mux2_1 _11622_ (.A0(_06554_),
    .A1(\core_busio.mem_address[28] ),
    .S(net409),
    .X(_01686_));
 sky130_fd_sc_hd__o21a_1 _11623_ (.A1(net633),
    .A2(_05697_),
    .B1(_06548_),
    .X(_06555_));
 sky130_fd_sc_hd__xnor2_1 _11624_ (.A(_05702_),
    .B(_06555_),
    .Y(_06556_));
 sky130_fd_sc_hd__nor2_1 _11625_ (.A(_05704_),
    .B(_06556_),
    .Y(_06557_));
 sky130_fd_sc_hd__nand2_1 _11626_ (.A(_05704_),
    .B(_06556_),
    .Y(_06558_));
 sky130_fd_sc_hd__nand2b_1 _11627_ (.A_N(_06557_),
    .B(_06558_),
    .Y(_06559_));
 sky130_fd_sc_hd__a2bb2o_2 _11628_ (.A1_N(_06551_),
    .A2_N(_06553_),
    .B1(_05699_),
    .B2(_06550_),
    .X(_06560_));
 sky130_fd_sc_hd__xnor2_1 _11629_ (.A(_06559_),
    .B(_06560_),
    .Y(_06561_));
 sky130_fd_sc_hd__mux2_1 _11630_ (.A0(_06561_),
    .A1(\core_busio.mem_address[29] ),
    .S(net409),
    .X(_01687_));
 sky130_fd_sc_hd__a21boi_4 _11631_ (.A1(net459),
    .A2(_05702_),
    .B1_N(_06555_),
    .Y(_06562_));
 sky130_fd_sc_hd__xnor2_2 _11632_ (.A(_05690_),
    .B(_06562_),
    .Y(_06563_));
 sky130_fd_sc_hd__xnor2_2 _11633_ (.A(_05688_),
    .B(_06563_),
    .Y(_06564_));
 sky130_fd_sc_hd__o21ai_2 _11634_ (.A1(_06557_),
    .A2(_06560_),
    .B1(_06558_),
    .Y(_06565_));
 sky130_fd_sc_hd__xor2_1 _11635_ (.A(_06564_),
    .B(_06565_),
    .X(_06566_));
 sky130_fd_sc_hd__mux2_1 _11636_ (.A0(_06566_),
    .A1(\core_busio.mem_address[30] ),
    .S(net409),
    .X(_01688_));
 sky130_fd_sc_hd__o22a_1 _11637_ (.A1(_05688_),
    .A2(_06563_),
    .B1(_06564_),
    .B2(_06565_),
    .X(_06567_));
 sky130_fd_sc_hd__o21ai_1 _11638_ (.A1(net632),
    .A2(_05691_),
    .B1(_06562_),
    .Y(_06568_));
 sky130_fd_sc_hd__xnor2_1 _11639_ (.A(_05685_),
    .B(_06568_),
    .Y(_06569_));
 sky130_fd_sc_hd__xnor2_1 _11640_ (.A(_06567_),
    .B(_06569_),
    .Y(_06570_));
 sky130_fd_sc_hd__mux2_1 _11641_ (.A0(_06570_),
    .A1(\core_busio.mem_address[31] ),
    .S(net409),
    .X(_01689_));
 sky130_fd_sc_hd__mux2_1 _11642_ (.A0(\core_pipeline.execute_to_memory_wfi ),
    .A1(\core_pipeline.decode_to_execute_wfi ),
    .S(net147),
    .X(_01690_));
 sky130_fd_sc_hd__or4_4 _11643_ (.A(\core_pipeline.memory_to_writeback_rd_address[2] ),
    .B(\core_pipeline.memory_to_writeback_rd_address[3] ),
    .C(_03912_),
    .D(_05589_),
    .X(_06571_));
 sky130_fd_sc_hd__mux2_1 _11644_ (.A0(net349),
    .A1(\core_pipeline.pipeline_registers.registers[17][0] ),
    .S(net179),
    .X(_01691_));
 sky130_fd_sc_hd__mux2_1 _11645_ (.A0(net346),
    .A1(\core_pipeline.pipeline_registers.registers[17][1] ),
    .S(net180),
    .X(_01692_));
 sky130_fd_sc_hd__mux2_1 _11646_ (.A0(net345),
    .A1(\core_pipeline.pipeline_registers.registers[17][2] ),
    .S(net180),
    .X(_01693_));
 sky130_fd_sc_hd__mux2_1 _11647_ (.A0(net343),
    .A1(\core_pipeline.pipeline_registers.registers[17][3] ),
    .S(net179),
    .X(_01694_));
 sky130_fd_sc_hd__mux2_1 _11648_ (.A0(net341),
    .A1(\core_pipeline.pipeline_registers.registers[17][4] ),
    .S(net179),
    .X(_01695_));
 sky130_fd_sc_hd__mux2_1 _11649_ (.A0(net338),
    .A1(\core_pipeline.pipeline_registers.registers[17][5] ),
    .S(net180),
    .X(_01696_));
 sky130_fd_sc_hd__mux2_1 _11650_ (.A0(net336),
    .A1(\core_pipeline.pipeline_registers.registers[17][6] ),
    .S(net180),
    .X(_01697_));
 sky130_fd_sc_hd__mux2_1 _11651_ (.A0(net333),
    .A1(\core_pipeline.pipeline_registers.registers[17][7] ),
    .S(net179),
    .X(_01698_));
 sky130_fd_sc_hd__mux2_1 _11652_ (.A0(net331),
    .A1(\core_pipeline.pipeline_registers.registers[17][8] ),
    .S(net179),
    .X(_01699_));
 sky130_fd_sc_hd__mux2_1 _11653_ (.A0(net330),
    .A1(\core_pipeline.pipeline_registers.registers[17][9] ),
    .S(net179),
    .X(_01700_));
 sky130_fd_sc_hd__mux2_1 _11654_ (.A0(net327),
    .A1(\core_pipeline.pipeline_registers.registers[17][10] ),
    .S(net179),
    .X(_01701_));
 sky130_fd_sc_hd__mux2_1 _11655_ (.A0(net326),
    .A1(\core_pipeline.pipeline_registers.registers[17][11] ),
    .S(net179),
    .X(_01702_));
 sky130_fd_sc_hd__mux2_1 _11656_ (.A0(net323),
    .A1(\core_pipeline.pipeline_registers.registers[17][12] ),
    .S(net179),
    .X(_01703_));
 sky130_fd_sc_hd__mux2_1 _11657_ (.A0(net321),
    .A1(\core_pipeline.pipeline_registers.registers[17][13] ),
    .S(net179),
    .X(_01704_));
 sky130_fd_sc_hd__mux2_1 _11658_ (.A0(net319),
    .A1(\core_pipeline.pipeline_registers.registers[17][14] ),
    .S(net179),
    .X(_01705_));
 sky130_fd_sc_hd__mux2_1 _11659_ (.A0(net318),
    .A1(\core_pipeline.pipeline_registers.registers[17][15] ),
    .S(net179),
    .X(_01706_));
 sky130_fd_sc_hd__mux2_1 _11660_ (.A0(net316),
    .A1(\core_pipeline.pipeline_registers.registers[17][16] ),
    .S(net179),
    .X(_01707_));
 sky130_fd_sc_hd__mux2_1 _11661_ (.A0(net313),
    .A1(\core_pipeline.pipeline_registers.registers[17][17] ),
    .S(net180),
    .X(_01708_));
 sky130_fd_sc_hd__mux2_1 _11662_ (.A0(net310),
    .A1(\core_pipeline.pipeline_registers.registers[17][18] ),
    .S(net180),
    .X(_01709_));
 sky130_fd_sc_hd__mux2_1 _11663_ (.A0(net309),
    .A1(\core_pipeline.pipeline_registers.registers[17][19] ),
    .S(net180),
    .X(_01710_));
 sky130_fd_sc_hd__mux2_1 _11664_ (.A0(net305),
    .A1(\core_pipeline.pipeline_registers.registers[17][20] ),
    .S(net180),
    .X(_01711_));
 sky130_fd_sc_hd__mux2_1 _11665_ (.A0(net303),
    .A1(\core_pipeline.pipeline_registers.registers[17][21] ),
    .S(net180),
    .X(_01712_));
 sky130_fd_sc_hd__mux2_1 _11666_ (.A0(net302),
    .A1(\core_pipeline.pipeline_registers.registers[17][22] ),
    .S(net179),
    .X(_01713_));
 sky130_fd_sc_hd__mux2_1 _11667_ (.A0(net299),
    .A1(\core_pipeline.pipeline_registers.registers[17][23] ),
    .S(net180),
    .X(_01714_));
 sky130_fd_sc_hd__mux2_1 _11668_ (.A0(net298),
    .A1(\core_pipeline.pipeline_registers.registers[17][24] ),
    .S(net179),
    .X(_01715_));
 sky130_fd_sc_hd__mux2_1 _11669_ (.A0(net296),
    .A1(\core_pipeline.pipeline_registers.registers[17][25] ),
    .S(net179),
    .X(_01716_));
 sky130_fd_sc_hd__mux2_1 _11670_ (.A0(net293),
    .A1(\core_pipeline.pipeline_registers.registers[17][26] ),
    .S(net179),
    .X(_01717_));
 sky130_fd_sc_hd__mux2_1 _11671_ (.A0(net291),
    .A1(\core_pipeline.pipeline_registers.registers[17][27] ),
    .S(net180),
    .X(_01718_));
 sky130_fd_sc_hd__mux2_1 _11672_ (.A0(net289),
    .A1(\core_pipeline.pipeline_registers.registers[17][28] ),
    .S(net180),
    .X(_01719_));
 sky130_fd_sc_hd__mux2_1 _11673_ (.A0(net286),
    .A1(\core_pipeline.pipeline_registers.registers[17][29] ),
    .S(net180),
    .X(_01720_));
 sky130_fd_sc_hd__mux2_1 _11674_ (.A0(net285),
    .A1(\core_pipeline.pipeline_registers.registers[17][30] ),
    .S(net180),
    .X(_01721_));
 sky130_fd_sc_hd__mux2_1 _11675_ (.A0(net282),
    .A1(\core_pipeline.pipeline_registers.registers[17][31] ),
    .S(net180),
    .X(_01722_));
 sky130_fd_sc_hd__or4_4 _11676_ (.A(\core_pipeline.memory_to_writeback_rd_address[2] ),
    .B(\core_pipeline.memory_to_writeback_rd_address[3] ),
    .C(_03912_),
    .D(_04939_),
    .X(_06572_));
 sky130_fd_sc_hd__mux2_1 _11677_ (.A0(net349),
    .A1(\core_pipeline.pipeline_registers.registers[16][0] ),
    .S(net177),
    .X(_01723_));
 sky130_fd_sc_hd__mux2_1 _11678_ (.A0(net346),
    .A1(\core_pipeline.pipeline_registers.registers[16][1] ),
    .S(net178),
    .X(_01724_));
 sky130_fd_sc_hd__mux2_1 _11679_ (.A0(net345),
    .A1(\core_pipeline.pipeline_registers.registers[16][2] ),
    .S(net178),
    .X(_01725_));
 sky130_fd_sc_hd__mux2_1 _11680_ (.A0(net342),
    .A1(\core_pipeline.pipeline_registers.registers[16][3] ),
    .S(net177),
    .X(_01726_));
 sky130_fd_sc_hd__mux2_1 _11681_ (.A0(net341),
    .A1(\core_pipeline.pipeline_registers.registers[16][4] ),
    .S(net177),
    .X(_01727_));
 sky130_fd_sc_hd__mux2_1 _11682_ (.A0(net339),
    .A1(\core_pipeline.pipeline_registers.registers[16][5] ),
    .S(net178),
    .X(_01728_));
 sky130_fd_sc_hd__mux2_1 _11683_ (.A0(net336),
    .A1(\core_pipeline.pipeline_registers.registers[16][6] ),
    .S(net178),
    .X(_01729_));
 sky130_fd_sc_hd__mux2_1 _11684_ (.A0(net333),
    .A1(\core_pipeline.pipeline_registers.registers[16][7] ),
    .S(net177),
    .X(_01730_));
 sky130_fd_sc_hd__mux2_1 _11685_ (.A0(net331),
    .A1(\core_pipeline.pipeline_registers.registers[16][8] ),
    .S(net177),
    .X(_01731_));
 sky130_fd_sc_hd__mux2_1 _11686_ (.A0(net330),
    .A1(\core_pipeline.pipeline_registers.registers[16][9] ),
    .S(net177),
    .X(_01732_));
 sky130_fd_sc_hd__mux2_1 _11687_ (.A0(net327),
    .A1(\core_pipeline.pipeline_registers.registers[16][10] ),
    .S(net177),
    .X(_01733_));
 sky130_fd_sc_hd__mux2_1 _11688_ (.A0(net326),
    .A1(\core_pipeline.pipeline_registers.registers[16][11] ),
    .S(net177),
    .X(_01734_));
 sky130_fd_sc_hd__mux2_1 _11689_ (.A0(net324),
    .A1(\core_pipeline.pipeline_registers.registers[16][12] ),
    .S(net177),
    .X(_01735_));
 sky130_fd_sc_hd__mux2_1 _11690_ (.A0(net321),
    .A1(\core_pipeline.pipeline_registers.registers[16][13] ),
    .S(net177),
    .X(_01736_));
 sky130_fd_sc_hd__mux2_1 _11691_ (.A0(net319),
    .A1(\core_pipeline.pipeline_registers.registers[16][14] ),
    .S(net177),
    .X(_01737_));
 sky130_fd_sc_hd__mux2_1 _11692_ (.A0(net318),
    .A1(\core_pipeline.pipeline_registers.registers[16][15] ),
    .S(net177),
    .X(_01738_));
 sky130_fd_sc_hd__mux2_1 _11693_ (.A0(net316),
    .A1(\core_pipeline.pipeline_registers.registers[16][16] ),
    .S(net177),
    .X(_01739_));
 sky130_fd_sc_hd__mux2_1 _11694_ (.A0(net313),
    .A1(\core_pipeline.pipeline_registers.registers[16][17] ),
    .S(net178),
    .X(_01740_));
 sky130_fd_sc_hd__mux2_1 _11695_ (.A0(net310),
    .A1(\core_pipeline.pipeline_registers.registers[16][18] ),
    .S(net178),
    .X(_01741_));
 sky130_fd_sc_hd__mux2_1 _11696_ (.A0(net309),
    .A1(\core_pipeline.pipeline_registers.registers[16][19] ),
    .S(net178),
    .X(_01742_));
 sky130_fd_sc_hd__mux2_1 _11697_ (.A0(net305),
    .A1(\core_pipeline.pipeline_registers.registers[16][20] ),
    .S(net178),
    .X(_01743_));
 sky130_fd_sc_hd__mux2_1 _11698_ (.A0(net303),
    .A1(\core_pipeline.pipeline_registers.registers[16][21] ),
    .S(net178),
    .X(_01744_));
 sky130_fd_sc_hd__mux2_1 _11699_ (.A0(net302),
    .A1(\core_pipeline.pipeline_registers.registers[16][22] ),
    .S(net177),
    .X(_01745_));
 sky130_fd_sc_hd__mux2_1 _11700_ (.A0(net299),
    .A1(\core_pipeline.pipeline_registers.registers[16][23] ),
    .S(net178),
    .X(_01746_));
 sky130_fd_sc_hd__mux2_1 _11701_ (.A0(net298),
    .A1(\core_pipeline.pipeline_registers.registers[16][24] ),
    .S(net177),
    .X(_01747_));
 sky130_fd_sc_hd__mux2_1 _11702_ (.A0(net296),
    .A1(\core_pipeline.pipeline_registers.registers[16][25] ),
    .S(net177),
    .X(_01748_));
 sky130_fd_sc_hd__mux2_1 _11703_ (.A0(net293),
    .A1(\core_pipeline.pipeline_registers.registers[16][26] ),
    .S(net177),
    .X(_01749_));
 sky130_fd_sc_hd__mux2_1 _11704_ (.A0(net291),
    .A1(\core_pipeline.pipeline_registers.registers[16][27] ),
    .S(net178),
    .X(_01750_));
 sky130_fd_sc_hd__mux2_1 _11705_ (.A0(net289),
    .A1(\core_pipeline.pipeline_registers.registers[16][28] ),
    .S(net178),
    .X(_01751_));
 sky130_fd_sc_hd__mux2_1 _11706_ (.A0(net286),
    .A1(\core_pipeline.pipeline_registers.registers[16][29] ),
    .S(net178),
    .X(_01752_));
 sky130_fd_sc_hd__mux2_1 _11707_ (.A0(net284),
    .A1(\core_pipeline.pipeline_registers.registers[16][30] ),
    .S(net178),
    .X(_01753_));
 sky130_fd_sc_hd__mux2_1 _11708_ (.A0(net282),
    .A1(\core_pipeline.pipeline_registers.registers[16][31] ),
    .S(net178),
    .X(_01754_));
 sky130_fd_sc_hd__or3b_4 _11709_ (.A(\core_pipeline.memory_to_writeback_rd_address[4] ),
    .B(_04468_),
    .C_N(\core_pipeline.memory_to_writeback_rd_address[2] ),
    .X(_06573_));
 sky130_fd_sc_hd__nor2_8 _11710_ (.A(_03915_),
    .B(_06573_),
    .Y(_06574_));
 sky130_fd_sc_hd__mux2_1 _11711_ (.A0(\core_pipeline.pipeline_registers.registers[15][0] ),
    .A1(net348),
    .S(net175),
    .X(_01755_));
 sky130_fd_sc_hd__mux2_1 _11712_ (.A0(\core_pipeline.pipeline_registers.registers[15][1] ),
    .A1(net347),
    .S(net176),
    .X(_01756_));
 sky130_fd_sc_hd__mux2_1 _11713_ (.A0(\core_pipeline.pipeline_registers.registers[15][2] ),
    .A1(net344),
    .S(net176),
    .X(_01757_));
 sky130_fd_sc_hd__mux2_1 _11714_ (.A0(\core_pipeline.pipeline_registers.registers[15][3] ),
    .A1(net343),
    .S(net175),
    .X(_01758_));
 sky130_fd_sc_hd__mux2_1 _11715_ (.A0(\core_pipeline.pipeline_registers.registers[15][4] ),
    .A1(net340),
    .S(net175),
    .X(_01759_));
 sky130_fd_sc_hd__mux2_1 _11716_ (.A0(\core_pipeline.pipeline_registers.registers[15][5] ),
    .A1(net337),
    .S(net176),
    .X(_01760_));
 sky130_fd_sc_hd__mux2_1 _11717_ (.A0(\core_pipeline.pipeline_registers.registers[15][6] ),
    .A1(net335),
    .S(net176),
    .X(_01761_));
 sky130_fd_sc_hd__mux2_1 _11718_ (.A0(\core_pipeline.pipeline_registers.registers[15][7] ),
    .A1(net334),
    .S(net175),
    .X(_01762_));
 sky130_fd_sc_hd__mux2_1 _11719_ (.A0(\core_pipeline.pipeline_registers.registers[15][8] ),
    .A1(net331),
    .S(net175),
    .X(_01763_));
 sky130_fd_sc_hd__mux2_1 _11720_ (.A0(\core_pipeline.pipeline_registers.registers[15][9] ),
    .A1(net329),
    .S(net175),
    .X(_01764_));
 sky130_fd_sc_hd__mux2_1 _11721_ (.A0(\core_pipeline.pipeline_registers.registers[15][10] ),
    .A1(net327),
    .S(net175),
    .X(_01765_));
 sky130_fd_sc_hd__mux2_1 _11722_ (.A0(\core_pipeline.pipeline_registers.registers[15][11] ),
    .A1(net325),
    .S(net175),
    .X(_01766_));
 sky130_fd_sc_hd__mux2_1 _11723_ (.A0(\core_pipeline.pipeline_registers.registers[15][12] ),
    .A1(net323),
    .S(net175),
    .X(_01767_));
 sky130_fd_sc_hd__mux2_1 _11724_ (.A0(\core_pipeline.pipeline_registers.registers[15][13] ),
    .A1(net321),
    .S(net175),
    .X(_01768_));
 sky130_fd_sc_hd__mux2_1 _11725_ (.A0(\core_pipeline.pipeline_registers.registers[15][14] ),
    .A1(net320),
    .S(net175),
    .X(_01769_));
 sky130_fd_sc_hd__mux2_1 _11726_ (.A0(\core_pipeline.pipeline_registers.registers[15][15] ),
    .A1(net317),
    .S(net175),
    .X(_01770_));
 sky130_fd_sc_hd__mux2_1 _11727_ (.A0(\core_pipeline.pipeline_registers.registers[15][16] ),
    .A1(net315),
    .S(net175),
    .X(_01771_));
 sky130_fd_sc_hd__mux2_1 _11728_ (.A0(\core_pipeline.pipeline_registers.registers[15][17] ),
    .A1(net313),
    .S(net176),
    .X(_01772_));
 sky130_fd_sc_hd__mux2_1 _11729_ (.A0(\core_pipeline.pipeline_registers.registers[15][18] ),
    .A1(net311),
    .S(net176),
    .X(_01773_));
 sky130_fd_sc_hd__mux2_1 _11730_ (.A0(\core_pipeline.pipeline_registers.registers[15][19] ),
    .A1(net308),
    .S(net176),
    .X(_01774_));
 sky130_fd_sc_hd__mux2_1 _11731_ (.A0(\core_pipeline.pipeline_registers.registers[15][20] ),
    .A1(net305),
    .S(net176),
    .X(_01775_));
 sky130_fd_sc_hd__mux2_1 _11732_ (.A0(\core_pipeline.pipeline_registers.registers[15][21] ),
    .A1(net304),
    .S(net176),
    .X(_01776_));
 sky130_fd_sc_hd__mux2_1 _11733_ (.A0(\core_pipeline.pipeline_registers.registers[15][22] ),
    .A1(net301),
    .S(net176),
    .X(_01777_));
 sky130_fd_sc_hd__mux2_1 _11734_ (.A0(\core_pipeline.pipeline_registers.registers[15][23] ),
    .A1(net299),
    .S(net176),
    .X(_01778_));
 sky130_fd_sc_hd__mux2_1 _11735_ (.A0(\core_pipeline.pipeline_registers.registers[15][24] ),
    .A1(net297),
    .S(net175),
    .X(_01779_));
 sky130_fd_sc_hd__mux2_1 _11736_ (.A0(\core_pipeline.pipeline_registers.registers[15][25] ),
    .A1(net295),
    .S(net175),
    .X(_01780_));
 sky130_fd_sc_hd__mux2_1 _11737_ (.A0(\core_pipeline.pipeline_registers.registers[15][26] ),
    .A1(net294),
    .S(net175),
    .X(_01781_));
 sky130_fd_sc_hd__mux2_1 _11738_ (.A0(\core_pipeline.pipeline_registers.registers[15][27] ),
    .A1(net292),
    .S(net176),
    .X(_01782_));
 sky130_fd_sc_hd__mux2_1 _11739_ (.A0(\core_pipeline.pipeline_registers.registers[15][28] ),
    .A1(net289),
    .S(net176),
    .X(_01783_));
 sky130_fd_sc_hd__mux2_1 _11740_ (.A0(\core_pipeline.pipeline_registers.registers[15][29] ),
    .A1(net286),
    .S(net176),
    .X(_01784_));
 sky130_fd_sc_hd__mux2_1 _11741_ (.A0(\core_pipeline.pipeline_registers.registers[15][30] ),
    .A1(net285),
    .S(net175),
    .X(_01785_));
 sky130_fd_sc_hd__mux2_1 _11742_ (.A0(\core_pipeline.pipeline_registers.registers[15][31] ),
    .A1(net282),
    .S(net176),
    .X(_01786_));
 sky130_fd_sc_hd__or4_4 _11743_ (.A(\core_pipeline.memory_to_writeback_rd_address[2] ),
    .B(\core_pipeline.memory_to_writeback_rd_address[4] ),
    .C(_04468_),
    .D(_05589_),
    .X(_06575_));
 sky130_fd_sc_hd__mux2_1 _11744_ (.A0(net348),
    .A1(\core_pipeline.pipeline_registers.registers[9][0] ),
    .S(net173),
    .X(_01787_));
 sky130_fd_sc_hd__mux2_1 _11745_ (.A0(net346),
    .A1(\core_pipeline.pipeline_registers.registers[9][1] ),
    .S(net174),
    .X(_01788_));
 sky130_fd_sc_hd__mux2_1 _11746_ (.A0(net344),
    .A1(\core_pipeline.pipeline_registers.registers[9][2] ),
    .S(net174),
    .X(_01789_));
 sky130_fd_sc_hd__mux2_1 _11747_ (.A0(net343),
    .A1(\core_pipeline.pipeline_registers.registers[9][3] ),
    .S(net173),
    .X(_01790_));
 sky130_fd_sc_hd__mux2_1 _11748_ (.A0(net340),
    .A1(\core_pipeline.pipeline_registers.registers[9][4] ),
    .S(net173),
    .X(_01791_));
 sky130_fd_sc_hd__mux2_1 _11749_ (.A0(net337),
    .A1(\core_pipeline.pipeline_registers.registers[9][5] ),
    .S(net174),
    .X(_01792_));
 sky130_fd_sc_hd__mux2_1 _11750_ (.A0(net335),
    .A1(\core_pipeline.pipeline_registers.registers[9][6] ),
    .S(net174),
    .X(_01793_));
 sky130_fd_sc_hd__mux2_1 _11751_ (.A0(net334),
    .A1(\core_pipeline.pipeline_registers.registers[9][7] ),
    .S(net173),
    .X(_01794_));
 sky130_fd_sc_hd__mux2_1 _11752_ (.A0(net332),
    .A1(\core_pipeline.pipeline_registers.registers[9][8] ),
    .S(net173),
    .X(_01795_));
 sky130_fd_sc_hd__mux2_1 _11753_ (.A0(net329),
    .A1(\core_pipeline.pipeline_registers.registers[9][9] ),
    .S(net173),
    .X(_01796_));
 sky130_fd_sc_hd__mux2_1 _11754_ (.A0(net327),
    .A1(\core_pipeline.pipeline_registers.registers[9][10] ),
    .S(net173),
    .X(_01797_));
 sky130_fd_sc_hd__mux2_1 _11755_ (.A0(net325),
    .A1(\core_pipeline.pipeline_registers.registers[9][11] ),
    .S(net173),
    .X(_01798_));
 sky130_fd_sc_hd__mux2_1 _11756_ (.A0(net323),
    .A1(\core_pipeline.pipeline_registers.registers[9][12] ),
    .S(net173),
    .X(_01799_));
 sky130_fd_sc_hd__mux2_1 _11757_ (.A0(net321),
    .A1(\core_pipeline.pipeline_registers.registers[9][13] ),
    .S(net173),
    .X(_01800_));
 sky130_fd_sc_hd__mux2_1 _11758_ (.A0(net320),
    .A1(\core_pipeline.pipeline_registers.registers[9][14] ),
    .S(net173),
    .X(_01801_));
 sky130_fd_sc_hd__mux2_1 _11759_ (.A0(net318),
    .A1(\core_pipeline.pipeline_registers.registers[9][15] ),
    .S(net173),
    .X(_01802_));
 sky130_fd_sc_hd__mux2_1 _11760_ (.A0(net315),
    .A1(\core_pipeline.pipeline_registers.registers[9][16] ),
    .S(net173),
    .X(_01803_));
 sky130_fd_sc_hd__mux2_1 _11761_ (.A0(net312),
    .A1(\core_pipeline.pipeline_registers.registers[9][17] ),
    .S(net174),
    .X(_01804_));
 sky130_fd_sc_hd__mux2_1 _11762_ (.A0(net311),
    .A1(\core_pipeline.pipeline_registers.registers[9][18] ),
    .S(net174),
    .X(_01805_));
 sky130_fd_sc_hd__mux2_1 _11763_ (.A0(net308),
    .A1(\core_pipeline.pipeline_registers.registers[9][19] ),
    .S(net174),
    .X(_01806_));
 sky130_fd_sc_hd__mux2_1 _11764_ (.A0(net306),
    .A1(\core_pipeline.pipeline_registers.registers[9][20] ),
    .S(net174),
    .X(_01807_));
 sky130_fd_sc_hd__mux2_1 _11765_ (.A0(net303),
    .A1(\core_pipeline.pipeline_registers.registers[9][21] ),
    .S(net174),
    .X(_01808_));
 sky130_fd_sc_hd__mux2_1 _11766_ (.A0(net301),
    .A1(\core_pipeline.pipeline_registers.registers[9][22] ),
    .S(net174),
    .X(_01809_));
 sky130_fd_sc_hd__mux2_1 _11767_ (.A0(net300),
    .A1(\core_pipeline.pipeline_registers.registers[9][23] ),
    .S(net174),
    .X(_01810_));
 sky130_fd_sc_hd__mux2_1 _11768_ (.A0(net298),
    .A1(\core_pipeline.pipeline_registers.registers[9][24] ),
    .S(net173),
    .X(_01811_));
 sky130_fd_sc_hd__mux2_1 _11769_ (.A0(net295),
    .A1(\core_pipeline.pipeline_registers.registers[9][25] ),
    .S(net173),
    .X(_01812_));
 sky130_fd_sc_hd__mux2_1 _11770_ (.A0(net293),
    .A1(\core_pipeline.pipeline_registers.registers[9][26] ),
    .S(net173),
    .X(_01813_));
 sky130_fd_sc_hd__mux2_1 _11771_ (.A0(net292),
    .A1(\core_pipeline.pipeline_registers.registers[9][27] ),
    .S(net174),
    .X(_01814_));
 sky130_fd_sc_hd__mux2_1 _11772_ (.A0(net289),
    .A1(\core_pipeline.pipeline_registers.registers[9][28] ),
    .S(net174),
    .X(_01815_));
 sky130_fd_sc_hd__mux2_1 _11773_ (.A0(net287),
    .A1(\core_pipeline.pipeline_registers.registers[9][29] ),
    .S(net174),
    .X(_01816_));
 sky130_fd_sc_hd__mux2_1 _11774_ (.A0(net284),
    .A1(\core_pipeline.pipeline_registers.registers[9][30] ),
    .S(net173),
    .X(_01817_));
 sky130_fd_sc_hd__mux2_1 _11775_ (.A0(net282),
    .A1(\core_pipeline.pipeline_registers.registers[9][31] ),
    .S(net174),
    .X(_01818_));
 sky130_fd_sc_hd__or2_1 _11776_ (.A(\core_pipeline.execute_to_memory_ecause[1] ),
    .B(_05825_),
    .X(_06576_));
 sky130_fd_sc_hd__nand2_1 _11777_ (.A(\core_pipeline.execute_to_memory_load ),
    .B(_05825_),
    .Y(_06577_));
 sky130_fd_sc_hd__a32o_1 _11778_ (.A1(_05826_),
    .A2(_06576_),
    .A3(_06577_),
    .B1(net458),
    .B2(\core_pipeline.memory_to_writeback_ecause[1] ),
    .X(_01819_));
 sky130_fd_sc_hd__a22o_1 _11779_ (.A1(\core_pipeline.memory_to_writeback_ecause[2] ),
    .A2(net458),
    .B1(_05825_),
    .B2(_05826_),
    .X(_01820_));
 sky130_fd_sc_hd__o21a_1 _11780_ (.A1(\core_pipeline.decode_to_execute_exception ),
    .A2(_05966_),
    .B1(net147),
    .X(_06578_));
 sky130_fd_sc_hd__inv_2 _11781_ (.A(_06578_),
    .Y(_06579_));
 sky130_fd_sc_hd__a22o_1 _11782_ (.A1(\core_pipeline.execute_to_memory_ecause[0] ),
    .A2(net133),
    .B1(_06578_),
    .B2(\core_pipeline.decode_to_execute_ecause[0] ),
    .X(_01821_));
 sky130_fd_sc_hd__o22a_1 _11783_ (.A1(\core_pipeline.execute_to_memory_ecause[1] ),
    .A2(net147),
    .B1(_06579_),
    .B2(\core_pipeline.decode_to_execute_ecause[1] ),
    .X(_01822_));
 sky130_fd_sc_hd__a22o_1 _11784_ (.A1(\core_pipeline.execute_to_memory_ecause[3] ),
    .A2(net133),
    .B1(_06578_),
    .B2(\core_pipeline.decode_to_execute_ecause[3] ),
    .X(_01823_));
 sky130_fd_sc_hd__nor2_8 _11785_ (.A(_04934_),
    .B(_06573_),
    .Y(_06580_));
 sky130_fd_sc_hd__mux2_1 _11786_ (.A0(\core_pipeline.pipeline_registers.registers[14][0] ),
    .A1(net348),
    .S(net171),
    .X(_01824_));
 sky130_fd_sc_hd__mux2_1 _11787_ (.A0(\core_pipeline.pipeline_registers.registers[14][1] ),
    .A1(net347),
    .S(net172),
    .X(_01825_));
 sky130_fd_sc_hd__mux2_1 _11788_ (.A0(\core_pipeline.pipeline_registers.registers[14][2] ),
    .A1(net344),
    .S(net172),
    .X(_01826_));
 sky130_fd_sc_hd__mux2_1 _11789_ (.A0(\core_pipeline.pipeline_registers.registers[14][3] ),
    .A1(net343),
    .S(net171),
    .X(_01827_));
 sky130_fd_sc_hd__mux2_1 _11790_ (.A0(\core_pipeline.pipeline_registers.registers[14][4] ),
    .A1(net340),
    .S(net171),
    .X(_01828_));
 sky130_fd_sc_hd__mux2_1 _11791_ (.A0(\core_pipeline.pipeline_registers.registers[14][5] ),
    .A1(net337),
    .S(net172),
    .X(_01829_));
 sky130_fd_sc_hd__mux2_1 _11792_ (.A0(\core_pipeline.pipeline_registers.registers[14][6] ),
    .A1(net335),
    .S(net172),
    .X(_01830_));
 sky130_fd_sc_hd__mux2_1 _11793_ (.A0(\core_pipeline.pipeline_registers.registers[14][7] ),
    .A1(net334),
    .S(net171),
    .X(_01831_));
 sky130_fd_sc_hd__mux2_1 _11794_ (.A0(\core_pipeline.pipeline_registers.registers[14][8] ),
    .A1(net331),
    .S(net171),
    .X(_01832_));
 sky130_fd_sc_hd__mux2_1 _11795_ (.A0(\core_pipeline.pipeline_registers.registers[14][9] ),
    .A1(net329),
    .S(net171),
    .X(_01833_));
 sky130_fd_sc_hd__mux2_1 _11796_ (.A0(\core_pipeline.pipeline_registers.registers[14][10] ),
    .A1(net327),
    .S(net171),
    .X(_01834_));
 sky130_fd_sc_hd__mux2_1 _11797_ (.A0(\core_pipeline.pipeline_registers.registers[14][11] ),
    .A1(net325),
    .S(net171),
    .X(_01835_));
 sky130_fd_sc_hd__mux2_1 _11798_ (.A0(\core_pipeline.pipeline_registers.registers[14][12] ),
    .A1(net323),
    .S(net171),
    .X(_01836_));
 sky130_fd_sc_hd__mux2_1 _11799_ (.A0(\core_pipeline.pipeline_registers.registers[14][13] ),
    .A1(net321),
    .S(net171),
    .X(_01837_));
 sky130_fd_sc_hd__mux2_1 _11800_ (.A0(\core_pipeline.pipeline_registers.registers[14][14] ),
    .A1(net320),
    .S(net171),
    .X(_01838_));
 sky130_fd_sc_hd__mux2_1 _11801_ (.A0(\core_pipeline.pipeline_registers.registers[14][15] ),
    .A1(net318),
    .S(net171),
    .X(_01839_));
 sky130_fd_sc_hd__mux2_1 _11802_ (.A0(\core_pipeline.pipeline_registers.registers[14][16] ),
    .A1(net315),
    .S(net171),
    .X(_01840_));
 sky130_fd_sc_hd__mux2_1 _11803_ (.A0(\core_pipeline.pipeline_registers.registers[14][17] ),
    .A1(net314),
    .S(net172),
    .X(_01841_));
 sky130_fd_sc_hd__mux2_1 _11804_ (.A0(\core_pipeline.pipeline_registers.registers[14][18] ),
    .A1(net311),
    .S(net172),
    .X(_01842_));
 sky130_fd_sc_hd__mux2_1 _11805_ (.A0(\core_pipeline.pipeline_registers.registers[14][19] ),
    .A1(net308),
    .S(net172),
    .X(_01843_));
 sky130_fd_sc_hd__mux2_1 _11806_ (.A0(\core_pipeline.pipeline_registers.registers[14][20] ),
    .A1(net305),
    .S(net172),
    .X(_01844_));
 sky130_fd_sc_hd__mux2_1 _11807_ (.A0(\core_pipeline.pipeline_registers.registers[14][21] ),
    .A1(net304),
    .S(net172),
    .X(_01845_));
 sky130_fd_sc_hd__mux2_1 _11808_ (.A0(\core_pipeline.pipeline_registers.registers[14][22] ),
    .A1(net301),
    .S(net172),
    .X(_01846_));
 sky130_fd_sc_hd__mux2_1 _11809_ (.A0(\core_pipeline.pipeline_registers.registers[14][23] ),
    .A1(net299),
    .S(net172),
    .X(_01847_));
 sky130_fd_sc_hd__mux2_1 _11810_ (.A0(\core_pipeline.pipeline_registers.registers[14][24] ),
    .A1(net297),
    .S(net171),
    .X(_01848_));
 sky130_fd_sc_hd__mux2_1 _11811_ (.A0(\core_pipeline.pipeline_registers.registers[14][25] ),
    .A1(net295),
    .S(net171),
    .X(_01849_));
 sky130_fd_sc_hd__mux2_1 _11812_ (.A0(\core_pipeline.pipeline_registers.registers[14][26] ),
    .A1(net294),
    .S(net171),
    .X(_01850_));
 sky130_fd_sc_hd__mux2_1 _11813_ (.A0(\core_pipeline.pipeline_registers.registers[14][27] ),
    .A1(net292),
    .S(net172),
    .X(_01851_));
 sky130_fd_sc_hd__mux2_1 _11814_ (.A0(\core_pipeline.pipeline_registers.registers[14][28] ),
    .A1(net289),
    .S(net172),
    .X(_01852_));
 sky130_fd_sc_hd__mux2_1 _11815_ (.A0(\core_pipeline.pipeline_registers.registers[14][29] ),
    .A1(net286),
    .S(net172),
    .X(_01853_));
 sky130_fd_sc_hd__mux2_1 _11816_ (.A0(\core_pipeline.pipeline_registers.registers[14][30] ),
    .A1(net284),
    .S(net171),
    .X(_01854_));
 sky130_fd_sc_hd__mux2_1 _11817_ (.A0(\core_pipeline.pipeline_registers.registers[14][31] ),
    .A1(net282),
    .S(net172),
    .X(_01855_));
 sky130_fd_sc_hd__nor2_8 _11818_ (.A(_05589_),
    .B(_06573_),
    .Y(_06581_));
 sky130_fd_sc_hd__mux2_1 _11819_ (.A0(\core_pipeline.pipeline_registers.registers[13][0] ),
    .A1(net348),
    .S(net169),
    .X(_01856_));
 sky130_fd_sc_hd__mux2_1 _11820_ (.A0(\core_pipeline.pipeline_registers.registers[13][1] ),
    .A1(net347),
    .S(net170),
    .X(_01857_));
 sky130_fd_sc_hd__mux2_1 _11821_ (.A0(\core_pipeline.pipeline_registers.registers[13][2] ),
    .A1(net344),
    .S(net170),
    .X(_01858_));
 sky130_fd_sc_hd__mux2_1 _11822_ (.A0(\core_pipeline.pipeline_registers.registers[13][3] ),
    .A1(net343),
    .S(net169),
    .X(_01859_));
 sky130_fd_sc_hd__mux2_1 _11823_ (.A0(\core_pipeline.pipeline_registers.registers[13][4] ),
    .A1(net340),
    .S(net169),
    .X(_01860_));
 sky130_fd_sc_hd__mux2_1 _11824_ (.A0(\core_pipeline.pipeline_registers.registers[13][5] ),
    .A1(net337),
    .S(net170),
    .X(_01861_));
 sky130_fd_sc_hd__mux2_1 _11825_ (.A0(\core_pipeline.pipeline_registers.registers[13][6] ),
    .A1(net335),
    .S(net170),
    .X(_01862_));
 sky130_fd_sc_hd__mux2_1 _11826_ (.A0(\core_pipeline.pipeline_registers.registers[13][7] ),
    .A1(net334),
    .S(net169),
    .X(_01863_));
 sky130_fd_sc_hd__mux2_1 _11827_ (.A0(\core_pipeline.pipeline_registers.registers[13][8] ),
    .A1(net332),
    .S(net169),
    .X(_01864_));
 sky130_fd_sc_hd__mux2_1 _11828_ (.A0(\core_pipeline.pipeline_registers.registers[13][9] ),
    .A1(net329),
    .S(net169),
    .X(_01865_));
 sky130_fd_sc_hd__mux2_1 _11829_ (.A0(\core_pipeline.pipeline_registers.registers[13][10] ),
    .A1(net328),
    .S(net169),
    .X(_01866_));
 sky130_fd_sc_hd__mux2_1 _11830_ (.A0(\core_pipeline.pipeline_registers.registers[13][11] ),
    .A1(net325),
    .S(net169),
    .X(_01867_));
 sky130_fd_sc_hd__mux2_1 _11831_ (.A0(\core_pipeline.pipeline_registers.registers[13][12] ),
    .A1(net323),
    .S(net169),
    .X(_01868_));
 sky130_fd_sc_hd__mux2_1 _11832_ (.A0(\core_pipeline.pipeline_registers.registers[13][13] ),
    .A1(net321),
    .S(net169),
    .X(_01869_));
 sky130_fd_sc_hd__mux2_1 _11833_ (.A0(\core_pipeline.pipeline_registers.registers[13][14] ),
    .A1(net320),
    .S(net169),
    .X(_01870_));
 sky130_fd_sc_hd__mux2_1 _11834_ (.A0(\core_pipeline.pipeline_registers.registers[13][15] ),
    .A1(net317),
    .S(net169),
    .X(_01871_));
 sky130_fd_sc_hd__mux2_1 _11835_ (.A0(\core_pipeline.pipeline_registers.registers[13][16] ),
    .A1(net315),
    .S(net169),
    .X(_01872_));
 sky130_fd_sc_hd__mux2_1 _11836_ (.A0(\core_pipeline.pipeline_registers.registers[13][17] ),
    .A1(net313),
    .S(net170),
    .X(_01873_));
 sky130_fd_sc_hd__mux2_1 _11837_ (.A0(\core_pipeline.pipeline_registers.registers[13][18] ),
    .A1(net311),
    .S(net170),
    .X(_01874_));
 sky130_fd_sc_hd__mux2_1 _11838_ (.A0(\core_pipeline.pipeline_registers.registers[13][19] ),
    .A1(net308),
    .S(net170),
    .X(_01875_));
 sky130_fd_sc_hd__mux2_1 _11839_ (.A0(\core_pipeline.pipeline_registers.registers[13][20] ),
    .A1(net305),
    .S(net170),
    .X(_01876_));
 sky130_fd_sc_hd__mux2_1 _11840_ (.A0(\core_pipeline.pipeline_registers.registers[13][21] ),
    .A1(net303),
    .S(net170),
    .X(_01877_));
 sky130_fd_sc_hd__mux2_1 _11841_ (.A0(\core_pipeline.pipeline_registers.registers[13][22] ),
    .A1(net301),
    .S(net170),
    .X(_01878_));
 sky130_fd_sc_hd__mux2_1 _11842_ (.A0(\core_pipeline.pipeline_registers.registers[13][23] ),
    .A1(net299),
    .S(net170),
    .X(_01879_));
 sky130_fd_sc_hd__mux2_1 _11843_ (.A0(\core_pipeline.pipeline_registers.registers[13][24] ),
    .A1(net297),
    .S(net169),
    .X(_01880_));
 sky130_fd_sc_hd__mux2_1 _11844_ (.A0(\core_pipeline.pipeline_registers.registers[13][25] ),
    .A1(net295),
    .S(net169),
    .X(_01881_));
 sky130_fd_sc_hd__mux2_1 _11845_ (.A0(\core_pipeline.pipeline_registers.registers[13][26] ),
    .A1(net294),
    .S(net169),
    .X(_01882_));
 sky130_fd_sc_hd__mux2_1 _11846_ (.A0(\core_pipeline.pipeline_registers.registers[13][27] ),
    .A1(net292),
    .S(net170),
    .X(_01883_));
 sky130_fd_sc_hd__mux2_1 _11847_ (.A0(\core_pipeline.pipeline_registers.registers[13][28] ),
    .A1(net289),
    .S(net170),
    .X(_01884_));
 sky130_fd_sc_hd__mux2_1 _11848_ (.A0(\core_pipeline.pipeline_registers.registers[13][29] ),
    .A1(net286),
    .S(net170),
    .X(_01885_));
 sky130_fd_sc_hd__mux2_1 _11849_ (.A0(\core_pipeline.pipeline_registers.registers[13][30] ),
    .A1(net285),
    .S(net169),
    .X(_01886_));
 sky130_fd_sc_hd__mux2_1 _11850_ (.A0(\core_pipeline.pipeline_registers.registers[13][31] ),
    .A1(net283),
    .S(net170),
    .X(_01887_));
 sky130_fd_sc_hd__nor2_8 _11851_ (.A(_04939_),
    .B(_06573_),
    .Y(_06582_));
 sky130_fd_sc_hd__mux2_1 _11852_ (.A0(\core_pipeline.pipeline_registers.registers[12][0] ),
    .A1(net348),
    .S(net167),
    .X(_01888_));
 sky130_fd_sc_hd__mux2_1 _11853_ (.A0(\core_pipeline.pipeline_registers.registers[12][1] ),
    .A1(net346),
    .S(net168),
    .X(_01889_));
 sky130_fd_sc_hd__mux2_1 _11854_ (.A0(\core_pipeline.pipeline_registers.registers[12][2] ),
    .A1(net344),
    .S(net168),
    .X(_01890_));
 sky130_fd_sc_hd__mux2_1 _11855_ (.A0(\core_pipeline.pipeline_registers.registers[12][3] ),
    .A1(net343),
    .S(net167),
    .X(_01891_));
 sky130_fd_sc_hd__mux2_1 _11856_ (.A0(\core_pipeline.pipeline_registers.registers[12][4] ),
    .A1(net340),
    .S(net167),
    .X(_01892_));
 sky130_fd_sc_hd__mux2_1 _11857_ (.A0(\core_pipeline.pipeline_registers.registers[12][5] ),
    .A1(net337),
    .S(net168),
    .X(_01893_));
 sky130_fd_sc_hd__mux2_1 _11858_ (.A0(\core_pipeline.pipeline_registers.registers[12][6] ),
    .A1(net335),
    .S(net167),
    .X(_01894_));
 sky130_fd_sc_hd__mux2_1 _11859_ (.A0(\core_pipeline.pipeline_registers.registers[12][7] ),
    .A1(net334),
    .S(net167),
    .X(_01895_));
 sky130_fd_sc_hd__mux2_1 _11860_ (.A0(\core_pipeline.pipeline_registers.registers[12][8] ),
    .A1(net332),
    .S(net167),
    .X(_01896_));
 sky130_fd_sc_hd__mux2_1 _11861_ (.A0(\core_pipeline.pipeline_registers.registers[12][9] ),
    .A1(net329),
    .S(net167),
    .X(_01897_));
 sky130_fd_sc_hd__mux2_1 _11862_ (.A0(\core_pipeline.pipeline_registers.registers[12][10] ),
    .A1(net327),
    .S(net167),
    .X(_01898_));
 sky130_fd_sc_hd__mux2_1 _11863_ (.A0(\core_pipeline.pipeline_registers.registers[12][11] ),
    .A1(net325),
    .S(net167),
    .X(_01899_));
 sky130_fd_sc_hd__mux2_1 _11864_ (.A0(\core_pipeline.pipeline_registers.registers[12][12] ),
    .A1(net323),
    .S(net167),
    .X(_01900_));
 sky130_fd_sc_hd__mux2_1 _11865_ (.A0(\core_pipeline.pipeline_registers.registers[12][13] ),
    .A1(net321),
    .S(net167),
    .X(_01901_));
 sky130_fd_sc_hd__mux2_1 _11866_ (.A0(\core_pipeline.pipeline_registers.registers[12][14] ),
    .A1(net320),
    .S(net167),
    .X(_01902_));
 sky130_fd_sc_hd__mux2_1 _11867_ (.A0(\core_pipeline.pipeline_registers.registers[12][15] ),
    .A1(net317),
    .S(net167),
    .X(_01903_));
 sky130_fd_sc_hd__mux2_1 _11868_ (.A0(\core_pipeline.pipeline_registers.registers[12][16] ),
    .A1(net315),
    .S(net167),
    .X(_01904_));
 sky130_fd_sc_hd__mux2_1 _11869_ (.A0(\core_pipeline.pipeline_registers.registers[12][17] ),
    .A1(net313),
    .S(net168),
    .X(_01905_));
 sky130_fd_sc_hd__mux2_1 _11870_ (.A0(\core_pipeline.pipeline_registers.registers[12][18] ),
    .A1(net311),
    .S(net168),
    .X(_01906_));
 sky130_fd_sc_hd__mux2_1 _11871_ (.A0(\core_pipeline.pipeline_registers.registers[12][19] ),
    .A1(net309),
    .S(net168),
    .X(_01907_));
 sky130_fd_sc_hd__mux2_1 _11872_ (.A0(\core_pipeline.pipeline_registers.registers[12][20] ),
    .A1(net305),
    .S(net168),
    .X(_01908_));
 sky130_fd_sc_hd__mux2_1 _11873_ (.A0(\core_pipeline.pipeline_registers.registers[12][21] ),
    .A1(net303),
    .S(net168),
    .X(_01909_));
 sky130_fd_sc_hd__mux2_1 _11874_ (.A0(\core_pipeline.pipeline_registers.registers[12][22] ),
    .A1(net301),
    .S(net168),
    .X(_01910_));
 sky130_fd_sc_hd__mux2_1 _11875_ (.A0(\core_pipeline.pipeline_registers.registers[12][23] ),
    .A1(net299),
    .S(net168),
    .X(_01911_));
 sky130_fd_sc_hd__mux2_1 _11876_ (.A0(\core_pipeline.pipeline_registers.registers[12][24] ),
    .A1(net297),
    .S(net167),
    .X(_01912_));
 sky130_fd_sc_hd__mux2_1 _11877_ (.A0(\core_pipeline.pipeline_registers.registers[12][25] ),
    .A1(net295),
    .S(net167),
    .X(_01913_));
 sky130_fd_sc_hd__mux2_1 _11878_ (.A0(\core_pipeline.pipeline_registers.registers[12][26] ),
    .A1(net293),
    .S(net167),
    .X(_01914_));
 sky130_fd_sc_hd__mux2_1 _11879_ (.A0(\core_pipeline.pipeline_registers.registers[12][27] ),
    .A1(net292),
    .S(net168),
    .X(_01915_));
 sky130_fd_sc_hd__mux2_1 _11880_ (.A0(\core_pipeline.pipeline_registers.registers[12][28] ),
    .A1(net290),
    .S(net168),
    .X(_01916_));
 sky130_fd_sc_hd__mux2_1 _11881_ (.A0(\core_pipeline.pipeline_registers.registers[12][29] ),
    .A1(net286),
    .S(net168),
    .X(_01917_));
 sky130_fd_sc_hd__mux2_1 _11882_ (.A0(\core_pipeline.pipeline_registers.registers[12][30] ),
    .A1(net285),
    .S(net168),
    .X(_01918_));
 sky130_fd_sc_hd__mux2_1 _11883_ (.A0(\core_pipeline.pipeline_registers.registers[12][31] ),
    .A1(net283),
    .S(net168),
    .X(_01919_));
 sky130_fd_sc_hd__a22o_1 _11884_ (.A1(\core_pipeline.memory_to_writeback_ecause[3] ),
    .A2(net458),
    .B1(_05827_),
    .B2(\core_pipeline.execute_to_memory_ecause[3] ),
    .X(_01920_));
 sky130_fd_sc_hd__mux4_1 _11885_ (.A0(\core_pipeline.pipeline_registers.registers[4][0] ),
    .A1(\core_pipeline.pipeline_registers.registers[5][0] ),
    .A2(\core_pipeline.pipeline_registers.registers[6][0] ),
    .A3(\core_pipeline.pipeline_registers.registers[7][0] ),
    .S0(net604),
    .S1(net582),
    .X(_06583_));
 sky130_fd_sc_hd__mux4_1 _11886_ (.A0(\core_pipeline.pipeline_registers.registers[0][0] ),
    .A1(\core_pipeline.pipeline_registers.registers[1][0] ),
    .A2(\core_pipeline.pipeline_registers.registers[2][0] ),
    .A3(\core_pipeline.pipeline_registers.registers[3][0] ),
    .S0(net603),
    .S1(net582),
    .X(_06584_));
 sky130_fd_sc_hd__mux4_1 _11887_ (.A0(\core_pipeline.pipeline_registers.registers[20][0] ),
    .A1(\core_pipeline.pipeline_registers.registers[21][0] ),
    .A2(\core_pipeline.pipeline_registers.registers[22][0] ),
    .A3(\core_pipeline.pipeline_registers.registers[23][0] ),
    .S0(net604),
    .S1(net582),
    .X(_06585_));
 sky130_fd_sc_hd__mux4_1 _11888_ (.A0(\core_pipeline.pipeline_registers.registers[16][0] ),
    .A1(\core_pipeline.pipeline_registers.registers[17][0] ),
    .A2(\core_pipeline.pipeline_registers.registers[18][0] ),
    .A3(\core_pipeline.pipeline_registers.registers[19][0] ),
    .S0(net603),
    .S1(net583),
    .X(_06586_));
 sky130_fd_sc_hd__mux2_1 _11889_ (.A0(_06583_),
    .A1(_06584_),
    .S(net472),
    .X(_06587_));
 sky130_fd_sc_hd__mux4_1 _11890_ (.A0(\core_pipeline.pipeline_registers.registers[8][0] ),
    .A1(\core_pipeline.pipeline_registers.registers[9][0] ),
    .A2(\core_pipeline.pipeline_registers.registers[10][0] ),
    .A3(\core_pipeline.pipeline_registers.registers[11][0] ),
    .S0(net603),
    .S1(net582),
    .X(_06588_));
 sky130_fd_sc_hd__mux4_1 _11891_ (.A0(\core_pipeline.pipeline_registers.registers[12][0] ),
    .A1(\core_pipeline.pipeline_registers.registers[13][0] ),
    .A2(\core_pipeline.pipeline_registers.registers[14][0] ),
    .A3(\core_pipeline.pipeline_registers.registers[15][0] ),
    .S0(net603),
    .S1(net582),
    .X(_06589_));
 sky130_fd_sc_hd__or2_1 _11892_ (.A(net472),
    .B(_06589_),
    .X(_06590_));
 sky130_fd_sc_hd__o21a_1 _11893_ (.A1(net576),
    .A2(_06588_),
    .B1(net570),
    .X(_06591_));
 sky130_fd_sc_hd__a221o_1 _11894_ (.A1(net468),
    .A2(_06587_),
    .B1(_06590_),
    .B2(_06591_),
    .C1(net567),
    .X(_06592_));
 sky130_fd_sc_hd__mux2_1 _11895_ (.A0(\core_pipeline.pipeline_registers.registers[30][0] ),
    .A1(\core_pipeline.pipeline_registers.registers[31][0] ),
    .S(net607),
    .X(_06593_));
 sky130_fd_sc_hd__and2_1 _11896_ (.A(net586),
    .B(_06593_),
    .X(_06594_));
 sky130_fd_sc_hd__mux2_1 _11897_ (.A0(\core_pipeline.pipeline_registers.registers[28][0] ),
    .A1(\core_pipeline.pipeline_registers.registers[29][0] ),
    .S(net607),
    .X(_06595_));
 sky130_fd_sc_hd__a21o_1 _11898_ (.A1(net482),
    .A2(_06595_),
    .B1(net472),
    .X(_06596_));
 sky130_fd_sc_hd__mux2_1 _11899_ (.A0(\core_pipeline.pipeline_registers.registers[26][0] ),
    .A1(\core_pipeline.pipeline_registers.registers[27][0] ),
    .S(net607),
    .X(_06597_));
 sky130_fd_sc_hd__and2_1 _11900_ (.A(net586),
    .B(_06597_),
    .X(_06598_));
 sky130_fd_sc_hd__mux2_1 _11901_ (.A0(\core_pipeline.pipeline_registers.registers[24][0] ),
    .A1(\core_pipeline.pipeline_registers.registers[25][0] ),
    .S(net607),
    .X(_06599_));
 sky130_fd_sc_hd__a21o_1 _11902_ (.A1(net482),
    .A2(_06599_),
    .B1(net576),
    .X(_06600_));
 sky130_fd_sc_hd__o221a_1 _11903_ (.A1(_06594_),
    .A2(_06596_),
    .B1(_06598_),
    .B2(_06600_),
    .C1(net570),
    .X(_06601_));
 sky130_fd_sc_hd__mux2_1 _11904_ (.A0(_06585_),
    .A1(_06586_),
    .S(net472),
    .X(_06602_));
 sky130_fd_sc_hd__a211o_1 _11905_ (.A1(net468),
    .A2(_06602_),
    .B1(_06601_),
    .C1(net467),
    .X(_06603_));
 sky130_fd_sc_hd__and3_4 _11906_ (.A(net144),
    .B(_06592_),
    .C(_06603_),
    .X(_06604_));
 sky130_fd_sc_hd__a21o_1 _11907_ (.A1(\core_pipeline.decode_to_execute_rs1_data[0] ),
    .A2(net122),
    .B1(_06604_),
    .X(_01921_));
 sky130_fd_sc_hd__mux4_1 _11908_ (.A0(\core_pipeline.pipeline_registers.registers[4][1] ),
    .A1(\core_pipeline.pipeline_registers.registers[5][1] ),
    .A2(\core_pipeline.pipeline_registers.registers[6][1] ),
    .A3(\core_pipeline.pipeline_registers.registers[7][1] ),
    .S0(net624),
    .S1(net601),
    .X(_06605_));
 sky130_fd_sc_hd__mux4_1 _11909_ (.A0(\core_pipeline.pipeline_registers.registers[0][1] ),
    .A1(\core_pipeline.pipeline_registers.registers[1][1] ),
    .A2(\core_pipeline.pipeline_registers.registers[2][1] ),
    .A3(\core_pipeline.pipeline_registers.registers[3][1] ),
    .S0(net626),
    .S1(net602),
    .X(_06606_));
 sky130_fd_sc_hd__mux4_1 _11910_ (.A0(\core_pipeline.pipeline_registers.registers[20][1] ),
    .A1(\core_pipeline.pipeline_registers.registers[21][1] ),
    .A2(\core_pipeline.pipeline_registers.registers[22][1] ),
    .A3(\core_pipeline.pipeline_registers.registers[23][1] ),
    .S0(net626),
    .S1(net594),
    .X(_06607_));
 sky130_fd_sc_hd__mux4_1 _11911_ (.A0(\core_pipeline.pipeline_registers.registers[16][1] ),
    .A1(\core_pipeline.pipeline_registers.registers[17][1] ),
    .A2(\core_pipeline.pipeline_registers.registers[18][1] ),
    .A3(\core_pipeline.pipeline_registers.registers[19][1] ),
    .S0(net621),
    .S1(net598),
    .X(_06608_));
 sky130_fd_sc_hd__mux2_1 _11912_ (.A0(_06605_),
    .A1(_06606_),
    .S(net479),
    .X(_06609_));
 sky130_fd_sc_hd__mux4_1 _11913_ (.A0(\core_pipeline.pipeline_registers.registers[8][1] ),
    .A1(\core_pipeline.pipeline_registers.registers[9][1] ),
    .A2(\core_pipeline.pipeline_registers.registers[10][1] ),
    .A3(\core_pipeline.pipeline_registers.registers[11][1] ),
    .S0(net624),
    .S1(net601),
    .X(_06610_));
 sky130_fd_sc_hd__mux4_1 _11914_ (.A0(\core_pipeline.pipeline_registers.registers[12][1] ),
    .A1(\core_pipeline.pipeline_registers.registers[13][1] ),
    .A2(\core_pipeline.pipeline_registers.registers[14][1] ),
    .A3(\core_pipeline.pipeline_registers.registers[15][1] ),
    .S0(net624),
    .S1(net601),
    .X(_06611_));
 sky130_fd_sc_hd__or2_1 _11915_ (.A(net480),
    .B(_06611_),
    .X(_06612_));
 sky130_fd_sc_hd__o21a_1 _11916_ (.A1(net581),
    .A2(_06610_),
    .B1(net575),
    .X(_06613_));
 sky130_fd_sc_hd__a221o_1 _11917_ (.A1(net471),
    .A2(_06609_),
    .B1(_06612_),
    .B2(_06613_),
    .C1(net568),
    .X(_06614_));
 sky130_fd_sc_hd__mux2_1 _11918_ (.A0(\core_pipeline.pipeline_registers.registers[30][1] ),
    .A1(\core_pipeline.pipeline_registers.registers[31][1] ),
    .S(net621),
    .X(_06615_));
 sky130_fd_sc_hd__and2_1 _11919_ (.A(net598),
    .B(_06615_),
    .X(_06616_));
 sky130_fd_sc_hd__mux2_1 _11920_ (.A0(\core_pipeline.pipeline_registers.registers[28][1] ),
    .A1(\core_pipeline.pipeline_registers.registers[29][1] ),
    .S(net624),
    .X(_06617_));
 sky130_fd_sc_hd__a21o_1 _11921_ (.A1(net485),
    .A2(_06617_),
    .B1(net479),
    .X(_06618_));
 sky130_fd_sc_hd__mux2_1 _11922_ (.A0(\core_pipeline.pipeline_registers.registers[26][1] ),
    .A1(\core_pipeline.pipeline_registers.registers[27][1] ),
    .S(net621),
    .X(_06619_));
 sky130_fd_sc_hd__and2_1 _11923_ (.A(net598),
    .B(_06619_),
    .X(_06620_));
 sky130_fd_sc_hd__mux2_1 _11924_ (.A0(\core_pipeline.pipeline_registers.registers[24][1] ),
    .A1(\core_pipeline.pipeline_registers.registers[25][1] ),
    .S(net621),
    .X(_06621_));
 sky130_fd_sc_hd__a21o_1 _11925_ (.A1(net485),
    .A2(_06621_),
    .B1(net580),
    .X(_06622_));
 sky130_fd_sc_hd__o221a_1 _11926_ (.A1(_06616_),
    .A2(_06618_),
    .B1(_06620_),
    .B2(_06622_),
    .C1(net574),
    .X(_06623_));
 sky130_fd_sc_hd__mux2_1 _11927_ (.A0(_06607_),
    .A1(_06608_),
    .S(net479),
    .X(_06624_));
 sky130_fd_sc_hd__a211o_1 _11928_ (.A1(net471),
    .A2(_06624_),
    .B1(_06623_),
    .C1(net466),
    .X(_06625_));
 sky130_fd_sc_hd__and3_2 _11929_ (.A(net146),
    .B(_06614_),
    .C(_06625_),
    .X(_06626_));
 sky130_fd_sc_hd__a21o_1 _11930_ (.A1(\core_pipeline.decode_to_execute_rs1_data[1] ),
    .A2(net125),
    .B1(_06626_),
    .X(_01922_));
 sky130_fd_sc_hd__mux4_1 _11931_ (.A0(\core_pipeline.pipeline_registers.registers[4][2] ),
    .A1(\core_pipeline.pipeline_registers.registers[5][2] ),
    .A2(\core_pipeline.pipeline_registers.registers[6][2] ),
    .A3(\core_pipeline.pipeline_registers.registers[7][2] ),
    .S0(net619),
    .S1(net596),
    .X(_06627_));
 sky130_fd_sc_hd__mux4_1 _11932_ (.A0(\core_pipeline.pipeline_registers.registers[0][2] ),
    .A1(\core_pipeline.pipeline_registers.registers[1][2] ),
    .A2(\core_pipeline.pipeline_registers.registers[2][2] ),
    .A3(\core_pipeline.pipeline_registers.registers[3][2] ),
    .S0(net619),
    .S1(net596),
    .X(_06628_));
 sky130_fd_sc_hd__mux4_1 _11933_ (.A0(\core_pipeline.pipeline_registers.registers[20][2] ),
    .A1(\core_pipeline.pipeline_registers.registers[21][2] ),
    .A2(\core_pipeline.pipeline_registers.registers[22][2] ),
    .A3(\core_pipeline.pipeline_registers.registers[23][2] ),
    .S0(net616),
    .S1(net593),
    .X(_06629_));
 sky130_fd_sc_hd__mux4_1 _11934_ (.A0(\core_pipeline.pipeline_registers.registers[16][2] ),
    .A1(\core_pipeline.pipeline_registers.registers[17][2] ),
    .A2(\core_pipeline.pipeline_registers.registers[18][2] ),
    .A3(\core_pipeline.pipeline_registers.registers[19][2] ),
    .S0(net616),
    .S1(net593),
    .X(_06630_));
 sky130_fd_sc_hd__mux2_1 _11935_ (.A0(_06627_),
    .A1(_06628_),
    .S(net478),
    .X(_06631_));
 sky130_fd_sc_hd__mux4_2 _11936_ (.A0(\core_pipeline.pipeline_registers.registers[8][2] ),
    .A1(\core_pipeline.pipeline_registers.registers[9][2] ),
    .A2(\core_pipeline.pipeline_registers.registers[10][2] ),
    .A3(\core_pipeline.pipeline_registers.registers[11][2] ),
    .S0(net619),
    .S1(net596),
    .X(_06632_));
 sky130_fd_sc_hd__mux4_1 _11937_ (.A0(\core_pipeline.pipeline_registers.registers[12][2] ),
    .A1(\core_pipeline.pipeline_registers.registers[13][2] ),
    .A2(\core_pipeline.pipeline_registers.registers[14][2] ),
    .A3(\core_pipeline.pipeline_registers.registers[15][2] ),
    .S0(net619),
    .S1(net596),
    .X(_06633_));
 sky130_fd_sc_hd__or2_1 _11938_ (.A(net478),
    .B(_06633_),
    .X(_06634_));
 sky130_fd_sc_hd__o21a_1 _11939_ (.A1(net580),
    .A2(_06632_),
    .B1(net574),
    .X(_06635_));
 sky130_fd_sc_hd__a221o_1 _11940_ (.A1(net471),
    .A2(_06631_),
    .B1(_06634_),
    .B2(_06635_),
    .C1(net568),
    .X(_06636_));
 sky130_fd_sc_hd__mux2_1 _11941_ (.A0(\core_pipeline.pipeline_registers.registers[30][2] ),
    .A1(\core_pipeline.pipeline_registers.registers[31][2] ),
    .S(net619),
    .X(_06637_));
 sky130_fd_sc_hd__and2_1 _11942_ (.A(net596),
    .B(_06637_),
    .X(_06638_));
 sky130_fd_sc_hd__mux2_1 _11943_ (.A0(\core_pipeline.pipeline_registers.registers[28][2] ),
    .A1(\core_pipeline.pipeline_registers.registers[29][2] ),
    .S(net616),
    .X(_06639_));
 sky130_fd_sc_hd__a21o_1 _11944_ (.A1(net485),
    .A2(_06639_),
    .B1(net477),
    .X(_06640_));
 sky130_fd_sc_hd__mux2_1 _11945_ (.A0(\core_pipeline.pipeline_registers.registers[26][2] ),
    .A1(\core_pipeline.pipeline_registers.registers[27][2] ),
    .S(net619),
    .X(_06641_));
 sky130_fd_sc_hd__and2_1 _11946_ (.A(net593),
    .B(_06641_),
    .X(_06642_));
 sky130_fd_sc_hd__mux2_1 _11947_ (.A0(\core_pipeline.pipeline_registers.registers[24][2] ),
    .A1(\core_pipeline.pipeline_registers.registers[25][2] ),
    .S(net616),
    .X(_06643_));
 sky130_fd_sc_hd__a21o_1 _11948_ (.A1(net485),
    .A2(_06643_),
    .B1(net580),
    .X(_06644_));
 sky130_fd_sc_hd__o221a_1 _11949_ (.A1(_06638_),
    .A2(_06640_),
    .B1(_06642_),
    .B2(_06644_),
    .C1(net573),
    .X(_06645_));
 sky130_fd_sc_hd__mux2_1 _11950_ (.A0(_06629_),
    .A1(_06630_),
    .S(net477),
    .X(_06646_));
 sky130_fd_sc_hd__a211o_1 _11951_ (.A1(net470),
    .A2(_06646_),
    .B1(_06645_),
    .C1(net466),
    .X(_06647_));
 sky130_fd_sc_hd__and3_2 _11952_ (.A(net145),
    .B(_06636_),
    .C(_06647_),
    .X(_06648_));
 sky130_fd_sc_hd__a21o_1 _11953_ (.A1(\core_pipeline.decode_to_execute_rs1_data[2] ),
    .A2(net130),
    .B1(_06648_),
    .X(_01923_));
 sky130_fd_sc_hd__mux4_1 _11954_ (.A0(\core_pipeline.pipeline_registers.registers[4][3] ),
    .A1(\core_pipeline.pipeline_registers.registers[5][3] ),
    .A2(\core_pipeline.pipeline_registers.registers[6][3] ),
    .A3(\core_pipeline.pipeline_registers.registers[7][3] ),
    .S0(net608),
    .S1(net586),
    .X(_06649_));
 sky130_fd_sc_hd__mux4_1 _11955_ (.A0(\core_pipeline.pipeline_registers.registers[0][3] ),
    .A1(\core_pipeline.pipeline_registers.registers[1][3] ),
    .A2(\core_pipeline.pipeline_registers.registers[2][3] ),
    .A3(\core_pipeline.pipeline_registers.registers[3][3] ),
    .S0(net608),
    .S1(net586),
    .X(_06650_));
 sky130_fd_sc_hd__mux4_1 _11956_ (.A0(\core_pipeline.pipeline_registers.registers[20][3] ),
    .A1(\core_pipeline.pipeline_registers.registers[21][3] ),
    .A2(\core_pipeline.pipeline_registers.registers[22][3] ),
    .A3(\core_pipeline.pipeline_registers.registers[23][3] ),
    .S0(net608),
    .S1(net587),
    .X(_06651_));
 sky130_fd_sc_hd__mux4_1 _11957_ (.A0(\core_pipeline.pipeline_registers.registers[16][3] ),
    .A1(\core_pipeline.pipeline_registers.registers[17][3] ),
    .A2(\core_pipeline.pipeline_registers.registers[18][3] ),
    .A3(\core_pipeline.pipeline_registers.registers[19][3] ),
    .S0(net610),
    .S1(net589),
    .X(_06652_));
 sky130_fd_sc_hd__mux2_1 _11958_ (.A0(_06649_),
    .A1(_06650_),
    .S(net473),
    .X(_06653_));
 sky130_fd_sc_hd__mux4_1 _11959_ (.A0(\core_pipeline.pipeline_registers.registers[8][3] ),
    .A1(\core_pipeline.pipeline_registers.registers[9][3] ),
    .A2(\core_pipeline.pipeline_registers.registers[10][3] ),
    .A3(\core_pipeline.pipeline_registers.registers[11][3] ),
    .S0(net607),
    .S1(net586),
    .X(_06654_));
 sky130_fd_sc_hd__mux4_1 _11960_ (.A0(\core_pipeline.pipeline_registers.registers[12][3] ),
    .A1(\core_pipeline.pipeline_registers.registers[13][3] ),
    .A2(\core_pipeline.pipeline_registers.registers[14][3] ),
    .A3(\core_pipeline.pipeline_registers.registers[15][3] ),
    .S0(net608),
    .S1(net586),
    .X(_06655_));
 sky130_fd_sc_hd__or2_1 _11961_ (.A(net473),
    .B(_06655_),
    .X(_06656_));
 sky130_fd_sc_hd__o21a_1 _11962_ (.A1(net577),
    .A2(_06654_),
    .B1(net571),
    .X(_06657_));
 sky130_fd_sc_hd__a221o_1 _11963_ (.A1(net468),
    .A2(_06653_),
    .B1(_06656_),
    .B2(_06657_),
    .C1(net567),
    .X(_02294_));
 sky130_fd_sc_hd__mux2_1 _11964_ (.A0(\core_pipeline.pipeline_registers.registers[30][3] ),
    .A1(\core_pipeline.pipeline_registers.registers[31][3] ),
    .S(net608),
    .X(_02295_));
 sky130_fd_sc_hd__and2_1 _11965_ (.A(net587),
    .B(_02295_),
    .X(_02296_));
 sky130_fd_sc_hd__mux2_1 _11966_ (.A0(\core_pipeline.pipeline_registers.registers[28][3] ),
    .A1(\core_pipeline.pipeline_registers.registers[29][3] ),
    .S(net608),
    .X(_02297_));
 sky130_fd_sc_hd__a21o_1 _11967_ (.A1(net482),
    .A2(_02297_),
    .B1(net473),
    .X(_02298_));
 sky130_fd_sc_hd__mux2_1 _11968_ (.A0(\core_pipeline.pipeline_registers.registers[26][3] ),
    .A1(\core_pipeline.pipeline_registers.registers[27][3] ),
    .S(net608),
    .X(_02299_));
 sky130_fd_sc_hd__and2_1 _11969_ (.A(net587),
    .B(_02299_),
    .X(_02300_));
 sky130_fd_sc_hd__mux2_1 _11970_ (.A0(\core_pipeline.pipeline_registers.registers[24][3] ),
    .A1(\core_pipeline.pipeline_registers.registers[25][3] ),
    .S(net608),
    .X(_02301_));
 sky130_fd_sc_hd__a21o_1 _11971_ (.A1(net482),
    .A2(_02301_),
    .B1(net577),
    .X(_02302_));
 sky130_fd_sc_hd__o221a_1 _11972_ (.A1(_02296_),
    .A2(_02298_),
    .B1(_02300_),
    .B2(_02302_),
    .C1(net571),
    .X(_02303_));
 sky130_fd_sc_hd__mux2_1 _11973_ (.A0(_06651_),
    .A1(_06652_),
    .S(net473),
    .X(_02304_));
 sky130_fd_sc_hd__a211o_1 _11974_ (.A1(net468),
    .A2(_02304_),
    .B1(_02303_),
    .C1(net467),
    .X(_02305_));
 sky130_fd_sc_hd__and3_2 _11975_ (.A(net144),
    .B(_02294_),
    .C(_02305_),
    .X(_02306_));
 sky130_fd_sc_hd__a21o_1 _11976_ (.A1(\core_pipeline.decode_to_execute_rs1_data[3] ),
    .A2(net121),
    .B1(_02306_),
    .X(_01924_));
 sky130_fd_sc_hd__mux4_1 _11977_ (.A0(\core_pipeline.pipeline_registers.registers[4][4] ),
    .A1(\core_pipeline.pipeline_registers.registers[5][4] ),
    .A2(\core_pipeline.pipeline_registers.registers[6][4] ),
    .A3(\core_pipeline.pipeline_registers.registers[7][4] ),
    .S0(net603),
    .S1(net582),
    .X(_02307_));
 sky130_fd_sc_hd__mux4_1 _11978_ (.A0(\core_pipeline.pipeline_registers.registers[0][4] ),
    .A1(\core_pipeline.pipeline_registers.registers[1][4] ),
    .A2(\core_pipeline.pipeline_registers.registers[2][4] ),
    .A3(\core_pipeline.pipeline_registers.registers[3][4] ),
    .S0(net603),
    .S1(net582),
    .X(_02308_));
 sky130_fd_sc_hd__mux4_1 _11979_ (.A0(\core_pipeline.pipeline_registers.registers[20][4] ),
    .A1(\core_pipeline.pipeline_registers.registers[21][4] ),
    .A2(\core_pipeline.pipeline_registers.registers[22][4] ),
    .A3(\core_pipeline.pipeline_registers.registers[23][4] ),
    .S0(net604),
    .S1(net583),
    .X(_02309_));
 sky130_fd_sc_hd__mux4_1 _11980_ (.A0(\core_pipeline.pipeline_registers.registers[16][4] ),
    .A1(\core_pipeline.pipeline_registers.registers[17][4] ),
    .A2(\core_pipeline.pipeline_registers.registers[18][4] ),
    .A3(\core_pipeline.pipeline_registers.registers[19][4] ),
    .S0(net604),
    .S1(net583),
    .X(_02310_));
 sky130_fd_sc_hd__mux2_1 _11981_ (.A0(_02307_),
    .A1(_02308_),
    .S(net472),
    .X(_02311_));
 sky130_fd_sc_hd__mux4_1 _11982_ (.A0(\core_pipeline.pipeline_registers.registers[8][4] ),
    .A1(\core_pipeline.pipeline_registers.registers[9][4] ),
    .A2(\core_pipeline.pipeline_registers.registers[10][4] ),
    .A3(\core_pipeline.pipeline_registers.registers[11][4] ),
    .S0(net603),
    .S1(net582),
    .X(_02312_));
 sky130_fd_sc_hd__mux4_1 _11983_ (.A0(\core_pipeline.pipeline_registers.registers[12][4] ),
    .A1(\core_pipeline.pipeline_registers.registers[13][4] ),
    .A2(\core_pipeline.pipeline_registers.registers[14][4] ),
    .A3(\core_pipeline.pipeline_registers.registers[15][4] ),
    .S0(net603),
    .S1(net582),
    .X(_02313_));
 sky130_fd_sc_hd__or2_1 _11984_ (.A(net472),
    .B(_02313_),
    .X(_02314_));
 sky130_fd_sc_hd__o21a_1 _11985_ (.A1(net576),
    .A2(_02312_),
    .B1(net570),
    .X(_02315_));
 sky130_fd_sc_hd__a221o_1 _11986_ (.A1(net468),
    .A2(_02311_),
    .B1(_02314_),
    .B2(_02315_),
    .C1(net567),
    .X(_02316_));
 sky130_fd_sc_hd__mux2_1 _11987_ (.A0(\core_pipeline.pipeline_registers.registers[30][4] ),
    .A1(\core_pipeline.pipeline_registers.registers[31][4] ),
    .S(net608),
    .X(_02317_));
 sky130_fd_sc_hd__and2_1 _11988_ (.A(net583),
    .B(_02317_),
    .X(_02318_));
 sky130_fd_sc_hd__mux2_1 _11989_ (.A0(\core_pipeline.pipeline_registers.registers[28][4] ),
    .A1(\core_pipeline.pipeline_registers.registers[29][4] ),
    .S(net604),
    .X(_02319_));
 sky130_fd_sc_hd__a21o_1 _11990_ (.A1(net482),
    .A2(_02319_),
    .B1(net472),
    .X(_02320_));
 sky130_fd_sc_hd__mux2_1 _11991_ (.A0(\core_pipeline.pipeline_registers.registers[26][4] ),
    .A1(\core_pipeline.pipeline_registers.registers[27][4] ),
    .S(net604),
    .X(_02321_));
 sky130_fd_sc_hd__and2_1 _11992_ (.A(net583),
    .B(_02321_),
    .X(_02322_));
 sky130_fd_sc_hd__mux2_1 _11993_ (.A0(\core_pipeline.pipeline_registers.registers[24][4] ),
    .A1(\core_pipeline.pipeline_registers.registers[25][4] ),
    .S(net604),
    .X(_02323_));
 sky130_fd_sc_hd__a21o_1 _11994_ (.A1(net482),
    .A2(_02323_),
    .B1(net576),
    .X(_02324_));
 sky130_fd_sc_hd__o221a_1 _11995_ (.A1(_02318_),
    .A2(_02320_),
    .B1(_02322_),
    .B2(_02324_),
    .C1(net570),
    .X(_02325_));
 sky130_fd_sc_hd__mux2_1 _11996_ (.A0(_02309_),
    .A1(_02310_),
    .S(net472),
    .X(_02326_));
 sky130_fd_sc_hd__a211o_1 _11997_ (.A1(net468),
    .A2(_02326_),
    .B1(_02325_),
    .C1(net467),
    .X(_02327_));
 sky130_fd_sc_hd__and3_2 _11998_ (.A(net144),
    .B(_02316_),
    .C(_02327_),
    .X(_02328_));
 sky130_fd_sc_hd__a21o_1 _11999_ (.A1(\core_pipeline.decode_to_execute_rs1_data[4] ),
    .A2(net123),
    .B1(_02328_),
    .X(_01925_));
 sky130_fd_sc_hd__mux4_1 _12000_ (.A0(\core_pipeline.pipeline_registers.registers[4][5] ),
    .A1(\core_pipeline.pipeline_registers.registers[5][5] ),
    .A2(\core_pipeline.pipeline_registers.registers[6][5] ),
    .A3(\core_pipeline.pipeline_registers.registers[7][5] ),
    .S0(net616),
    .S1(net593),
    .X(_02329_));
 sky130_fd_sc_hd__mux4_1 _12001_ (.A0(\core_pipeline.pipeline_registers.registers[0][5] ),
    .A1(\core_pipeline.pipeline_registers.registers[1][5] ),
    .A2(\core_pipeline.pipeline_registers.registers[2][5] ),
    .A3(\core_pipeline.pipeline_registers.registers[3][5] ),
    .S0(net616),
    .S1(net593),
    .X(_02330_));
 sky130_fd_sc_hd__mux4_1 _12002_ (.A0(\core_pipeline.pipeline_registers.registers[20][5] ),
    .A1(\core_pipeline.pipeline_registers.registers[21][5] ),
    .A2(\core_pipeline.pipeline_registers.registers[22][5] ),
    .A3(\core_pipeline.pipeline_registers.registers[23][5] ),
    .S0(net623),
    .S1(net593),
    .X(_02331_));
 sky130_fd_sc_hd__mux4_1 _12003_ (.A0(\core_pipeline.pipeline_registers.registers[16][5] ),
    .A1(\core_pipeline.pipeline_registers.registers[17][5] ),
    .A2(\core_pipeline.pipeline_registers.registers[18][5] ),
    .A3(\core_pipeline.pipeline_registers.registers[19][5] ),
    .S0(net616),
    .S1(net592),
    .X(_02332_));
 sky130_fd_sc_hd__mux2_1 _12004_ (.A0(_02329_),
    .A1(_02330_),
    .S(net477),
    .X(_02333_));
 sky130_fd_sc_hd__mux4_1 _12005_ (.A0(\core_pipeline.pipeline_registers.registers[8][5] ),
    .A1(\core_pipeline.pipeline_registers.registers[9][5] ),
    .A2(\core_pipeline.pipeline_registers.registers[10][5] ),
    .A3(\core_pipeline.pipeline_registers.registers[11][5] ),
    .S0(net616),
    .S1(net593),
    .X(_02334_));
 sky130_fd_sc_hd__mux4_1 _12006_ (.A0(\core_pipeline.pipeline_registers.registers[12][5] ),
    .A1(\core_pipeline.pipeline_registers.registers[13][5] ),
    .A2(\core_pipeline.pipeline_registers.registers[14][5] ),
    .A3(\core_pipeline.pipeline_registers.registers[15][5] ),
    .S0(net616),
    .S1(net593),
    .X(_02335_));
 sky130_fd_sc_hd__or2_1 _12007_ (.A(net477),
    .B(_02335_),
    .X(_02336_));
 sky130_fd_sc_hd__o21a_1 _12008_ (.A1(net579),
    .A2(_02334_),
    .B1(net573),
    .X(_02337_));
 sky130_fd_sc_hd__a221o_1 _12009_ (.A1(net470),
    .A2(_02333_),
    .B1(_02336_),
    .B2(_02337_),
    .C1(net568),
    .X(_02338_));
 sky130_fd_sc_hd__mux2_1 _12010_ (.A0(\core_pipeline.pipeline_registers.registers[30][5] ),
    .A1(\core_pipeline.pipeline_registers.registers[31][5] ),
    .S(net616),
    .X(_02339_));
 sky130_fd_sc_hd__and2_1 _12011_ (.A(net592),
    .B(_02339_),
    .X(_02340_));
 sky130_fd_sc_hd__mux2_1 _12012_ (.A0(\core_pipeline.pipeline_registers.registers[28][5] ),
    .A1(\core_pipeline.pipeline_registers.registers[29][5] ),
    .S(net616),
    .X(_02341_));
 sky130_fd_sc_hd__a21o_1 _12013_ (.A1(net484),
    .A2(_02341_),
    .B1(net477),
    .X(_02342_));
 sky130_fd_sc_hd__mux2_1 _12014_ (.A0(\core_pipeline.pipeline_registers.registers[26][5] ),
    .A1(\core_pipeline.pipeline_registers.registers[27][5] ),
    .S(net616),
    .X(_02343_));
 sky130_fd_sc_hd__and2_1 _12015_ (.A(net592),
    .B(_02343_),
    .X(_02344_));
 sky130_fd_sc_hd__mux2_1 _12016_ (.A0(\core_pipeline.pipeline_registers.registers[24][5] ),
    .A1(\core_pipeline.pipeline_registers.registers[25][5] ),
    .S(net616),
    .X(_02345_));
 sky130_fd_sc_hd__a21o_1 _12017_ (.A1(net484),
    .A2(_02345_),
    .B1(net579),
    .X(_02346_));
 sky130_fd_sc_hd__o221a_1 _12018_ (.A1(_02340_),
    .A2(_02342_),
    .B1(_02344_),
    .B2(_02346_),
    .C1(net573),
    .X(_02347_));
 sky130_fd_sc_hd__mux2_1 _12019_ (.A0(_02331_),
    .A1(_02332_),
    .S(net477),
    .X(_02348_));
 sky130_fd_sc_hd__a211o_1 _12020_ (.A1(net470),
    .A2(_02348_),
    .B1(_02347_),
    .C1(net466),
    .X(_02349_));
 sky130_fd_sc_hd__and3_2 _12021_ (.A(net145),
    .B(_02338_),
    .C(_02349_),
    .X(_02350_));
 sky130_fd_sc_hd__a21o_1 _12022_ (.A1(\core_pipeline.decode_to_execute_rs1_data[5] ),
    .A2(net130),
    .B1(_02350_),
    .X(_01926_));
 sky130_fd_sc_hd__mux4_1 _12023_ (.A0(\core_pipeline.pipeline_registers.registers[4][6] ),
    .A1(\core_pipeline.pipeline_registers.registers[5][6] ),
    .A2(\core_pipeline.pipeline_registers.registers[6][6] ),
    .A3(\core_pipeline.pipeline_registers.registers[7][6] ),
    .S0(net608),
    .S1(net587),
    .X(_02351_));
 sky130_fd_sc_hd__mux4_1 _12024_ (.A0(\core_pipeline.pipeline_registers.registers[0][6] ),
    .A1(\core_pipeline.pipeline_registers.registers[1][6] ),
    .A2(\core_pipeline.pipeline_registers.registers[2][6] ),
    .A3(\core_pipeline.pipeline_registers.registers[3][6] ),
    .S0(net608),
    .S1(net587),
    .X(_02352_));
 sky130_fd_sc_hd__mux4_1 _12025_ (.A0(\core_pipeline.pipeline_registers.registers[20][6] ),
    .A1(\core_pipeline.pipeline_registers.registers[21][6] ),
    .A2(\core_pipeline.pipeline_registers.registers[22][6] ),
    .A3(\core_pipeline.pipeline_registers.registers[23][6] ),
    .S0(net615),
    .S1(net592),
    .X(_02353_));
 sky130_fd_sc_hd__mux4_1 _12026_ (.A0(\core_pipeline.pipeline_registers.registers[16][6] ),
    .A1(\core_pipeline.pipeline_registers.registers[17][6] ),
    .A2(\core_pipeline.pipeline_registers.registers[18][6] ),
    .A3(\core_pipeline.pipeline_registers.registers[19][6] ),
    .S0(net623),
    .S1(net592),
    .X(_02354_));
 sky130_fd_sc_hd__mux2_1 _12027_ (.A0(_02351_),
    .A1(_02352_),
    .S(net473),
    .X(_02355_));
 sky130_fd_sc_hd__mux4_1 _12028_ (.A0(\core_pipeline.pipeline_registers.registers[8][6] ),
    .A1(\core_pipeline.pipeline_registers.registers[9][6] ),
    .A2(\core_pipeline.pipeline_registers.registers[10][6] ),
    .A3(\core_pipeline.pipeline_registers.registers[11][6] ),
    .S0(net615),
    .S1(net592),
    .X(_02356_));
 sky130_fd_sc_hd__mux4_1 _12029_ (.A0(\core_pipeline.pipeline_registers.registers[12][6] ),
    .A1(\core_pipeline.pipeline_registers.registers[13][6] ),
    .A2(\core_pipeline.pipeline_registers.registers[14][6] ),
    .A3(\core_pipeline.pipeline_registers.registers[15][6] ),
    .S0(net608),
    .S1(net587),
    .X(_02357_));
 sky130_fd_sc_hd__or2_1 _12030_ (.A(net473),
    .B(_02357_),
    .X(_02358_));
 sky130_fd_sc_hd__o21a_1 _12031_ (.A1(net579),
    .A2(_02356_),
    .B1(net573),
    .X(_02359_));
 sky130_fd_sc_hd__a221o_1 _12032_ (.A1(net470),
    .A2(_02355_),
    .B1(_02358_),
    .B2(_02359_),
    .C1(net568),
    .X(_02360_));
 sky130_fd_sc_hd__mux2_1 _12033_ (.A0(\core_pipeline.pipeline_registers.registers[30][6] ),
    .A1(\core_pipeline.pipeline_registers.registers[31][6] ),
    .S(net615),
    .X(_02361_));
 sky130_fd_sc_hd__and2_1 _12034_ (.A(net592),
    .B(_02361_),
    .X(_02362_));
 sky130_fd_sc_hd__mux2_1 _12035_ (.A0(\core_pipeline.pipeline_registers.registers[28][6] ),
    .A1(\core_pipeline.pipeline_registers.registers[29][6] ),
    .S(net615),
    .X(_02363_));
 sky130_fd_sc_hd__a21o_1 _12036_ (.A1(net484),
    .A2(_02363_),
    .B1(net477),
    .X(_02364_));
 sky130_fd_sc_hd__mux2_1 _12037_ (.A0(\core_pipeline.pipeline_registers.registers[26][6] ),
    .A1(\core_pipeline.pipeline_registers.registers[27][6] ),
    .S(net615),
    .X(_02365_));
 sky130_fd_sc_hd__and2_1 _12038_ (.A(net592),
    .B(_02365_),
    .X(_02366_));
 sky130_fd_sc_hd__mux2_1 _12039_ (.A0(\core_pipeline.pipeline_registers.registers[24][6] ),
    .A1(\core_pipeline.pipeline_registers.registers[25][6] ),
    .S(net615),
    .X(_02367_));
 sky130_fd_sc_hd__a21o_1 _12040_ (.A1(net484),
    .A2(_02367_),
    .B1(net579),
    .X(_02368_));
 sky130_fd_sc_hd__o221a_1 _12041_ (.A1(_02362_),
    .A2(_02364_),
    .B1(_02366_),
    .B2(_02368_),
    .C1(net573),
    .X(_02369_));
 sky130_fd_sc_hd__mux2_1 _12042_ (.A0(_02353_),
    .A1(_02354_),
    .S(net477),
    .X(_02370_));
 sky130_fd_sc_hd__a211o_1 _12043_ (.A1(net470),
    .A2(_02370_),
    .B1(_02369_),
    .C1(net466),
    .X(_02371_));
 sky130_fd_sc_hd__and3_2 _12044_ (.A(net144),
    .B(_02360_),
    .C(_02371_),
    .X(_02372_));
 sky130_fd_sc_hd__a21o_1 _12045_ (.A1(\core_pipeline.decode_to_execute_rs1_data[6] ),
    .A2(net125),
    .B1(_02372_),
    .X(_01927_));
 sky130_fd_sc_hd__mux4_1 _12046_ (.A0(\core_pipeline.pipeline_registers.registers[4][7] ),
    .A1(\core_pipeline.pipeline_registers.registers[5][7] ),
    .A2(\core_pipeline.pipeline_registers.registers[6][7] ),
    .A3(\core_pipeline.pipeline_registers.registers[7][7] ),
    .S0(net603),
    .S1(net582),
    .X(_02373_));
 sky130_fd_sc_hd__mux4_1 _12047_ (.A0(\core_pipeline.pipeline_registers.registers[0][7] ),
    .A1(\core_pipeline.pipeline_registers.registers[1][7] ),
    .A2(\core_pipeline.pipeline_registers.registers[2][7] ),
    .A3(\core_pipeline.pipeline_registers.registers[3][7] ),
    .S0(net603),
    .S1(net582),
    .X(_02374_));
 sky130_fd_sc_hd__mux4_1 _12048_ (.A0(\core_pipeline.pipeline_registers.registers[20][7] ),
    .A1(\core_pipeline.pipeline_registers.registers[21][7] ),
    .A2(\core_pipeline.pipeline_registers.registers[22][7] ),
    .A3(\core_pipeline.pipeline_registers.registers[23][7] ),
    .S0(net609),
    .S1(net586),
    .X(_02375_));
 sky130_fd_sc_hd__mux4_1 _12049_ (.A0(\core_pipeline.pipeline_registers.registers[16][7] ),
    .A1(\core_pipeline.pipeline_registers.registers[17][7] ),
    .A2(\core_pipeline.pipeline_registers.registers[18][7] ),
    .A3(\core_pipeline.pipeline_registers.registers[19][7] ),
    .S0(net609),
    .S1(net588),
    .X(_02376_));
 sky130_fd_sc_hd__mux2_1 _12050_ (.A0(_02373_),
    .A1(_02374_),
    .S(net472),
    .X(_02377_));
 sky130_fd_sc_hd__mux4_1 _12051_ (.A0(\core_pipeline.pipeline_registers.registers[8][7] ),
    .A1(\core_pipeline.pipeline_registers.registers[9][7] ),
    .A2(\core_pipeline.pipeline_registers.registers[10][7] ),
    .A3(\core_pipeline.pipeline_registers.registers[11][7] ),
    .S0(net603),
    .S1(net582),
    .X(_02378_));
 sky130_fd_sc_hd__mux4_1 _12052_ (.A0(\core_pipeline.pipeline_registers.registers[12][7] ),
    .A1(\core_pipeline.pipeline_registers.registers[13][7] ),
    .A2(\core_pipeline.pipeline_registers.registers[14][7] ),
    .A3(\core_pipeline.pipeline_registers.registers[15][7] ),
    .S0(net603),
    .S1(net582),
    .X(_02379_));
 sky130_fd_sc_hd__or2_1 _12053_ (.A(net472),
    .B(_02379_),
    .X(_02380_));
 sky130_fd_sc_hd__o21a_1 _12054_ (.A1(net576),
    .A2(_02378_),
    .B1(net570),
    .X(_02381_));
 sky130_fd_sc_hd__a221o_4 _12055_ (.A1(net468),
    .A2(_02377_),
    .B1(_02380_),
    .B2(_02381_),
    .C1(net567),
    .X(_02382_));
 sky130_fd_sc_hd__mux2_1 _12056_ (.A0(\core_pipeline.pipeline_registers.registers[30][7] ),
    .A1(\core_pipeline.pipeline_registers.registers[31][7] ),
    .S(net610),
    .X(_02383_));
 sky130_fd_sc_hd__and2_1 _12057_ (.A(net588),
    .B(_02383_),
    .X(_02384_));
 sky130_fd_sc_hd__mux2_1 _12058_ (.A0(\core_pipeline.pipeline_registers.registers[28][7] ),
    .A1(\core_pipeline.pipeline_registers.registers[29][7] ),
    .S(net609),
    .X(_02385_));
 sky130_fd_sc_hd__a21o_1 _12059_ (.A1(net482),
    .A2(_02385_),
    .B1(net473),
    .X(_02386_));
 sky130_fd_sc_hd__mux2_1 _12060_ (.A0(\core_pipeline.pipeline_registers.registers[26][7] ),
    .A1(\core_pipeline.pipeline_registers.registers[27][7] ),
    .S(net609),
    .X(_02387_));
 sky130_fd_sc_hd__and2_1 _12061_ (.A(net589),
    .B(_02387_),
    .X(_02388_));
 sky130_fd_sc_hd__mux2_1 _12062_ (.A0(\core_pipeline.pipeline_registers.registers[24][7] ),
    .A1(\core_pipeline.pipeline_registers.registers[25][7] ),
    .S(net610),
    .X(_02389_));
 sky130_fd_sc_hd__a21o_1 _12063_ (.A1(net482),
    .A2(_02389_),
    .B1(net577),
    .X(_02390_));
 sky130_fd_sc_hd__o221a_1 _12064_ (.A1(_02384_),
    .A2(_02386_),
    .B1(_02388_),
    .B2(_02390_),
    .C1(net571),
    .X(_02391_));
 sky130_fd_sc_hd__mux2_1 _12065_ (.A0(_02375_),
    .A1(_02376_),
    .S(net473),
    .X(_02392_));
 sky130_fd_sc_hd__a211o_1 _12066_ (.A1(net468),
    .A2(_02392_),
    .B1(_02391_),
    .C1(net467),
    .X(_02393_));
 sky130_fd_sc_hd__and3_1 _12067_ (.A(net144),
    .B(_02382_),
    .C(_02393_),
    .X(_02394_));
 sky130_fd_sc_hd__a21o_1 _12068_ (.A1(\core_pipeline.decode_to_execute_rs1_data[7] ),
    .A2(net121),
    .B1(_02394_),
    .X(_01928_));
 sky130_fd_sc_hd__mux4_1 _12069_ (.A0(\core_pipeline.pipeline_registers.registers[4][8] ),
    .A1(\core_pipeline.pipeline_registers.registers[5][8] ),
    .A2(\core_pipeline.pipeline_registers.registers[6][8] ),
    .A3(\core_pipeline.pipeline_registers.registers[7][8] ),
    .S0(net611),
    .S1(net587),
    .X(_02395_));
 sky130_fd_sc_hd__mux4_1 _12070_ (.A0(\core_pipeline.pipeline_registers.registers[0][8] ),
    .A1(\core_pipeline.pipeline_registers.registers[1][8] ),
    .A2(\core_pipeline.pipeline_registers.registers[2][8] ),
    .A3(\core_pipeline.pipeline_registers.registers[3][8] ),
    .S0(net611),
    .S1(net587),
    .X(_02396_));
 sky130_fd_sc_hd__mux4_1 _12071_ (.A0(\core_pipeline.pipeline_registers.registers[20][8] ),
    .A1(\core_pipeline.pipeline_registers.registers[21][8] ),
    .A2(\core_pipeline.pipeline_registers.registers[22][8] ),
    .A3(\core_pipeline.pipeline_registers.registers[23][8] ),
    .S0(net608),
    .S1(net586),
    .X(_02397_));
 sky130_fd_sc_hd__mux4_1 _12072_ (.A0(\core_pipeline.pipeline_registers.registers[16][8] ),
    .A1(\core_pipeline.pipeline_registers.registers[17][8] ),
    .A2(\core_pipeline.pipeline_registers.registers[18][8] ),
    .A3(\core_pipeline.pipeline_registers.registers[19][8] ),
    .S0(net608),
    .S1(net586),
    .X(_02398_));
 sky130_fd_sc_hd__mux2_1 _12073_ (.A0(_02395_),
    .A1(_02396_),
    .S(net473),
    .X(_02399_));
 sky130_fd_sc_hd__mux4_1 _12074_ (.A0(\core_pipeline.pipeline_registers.registers[8][8] ),
    .A1(\core_pipeline.pipeline_registers.registers[9][8] ),
    .A2(\core_pipeline.pipeline_registers.registers[10][8] ),
    .A3(\core_pipeline.pipeline_registers.registers[11][8] ),
    .S0(net608),
    .S1(net587),
    .X(_02400_));
 sky130_fd_sc_hd__mux4_1 _12075_ (.A0(\core_pipeline.pipeline_registers.registers[12][8] ),
    .A1(\core_pipeline.pipeline_registers.registers[13][8] ),
    .A2(\core_pipeline.pipeline_registers.registers[14][8] ),
    .A3(\core_pipeline.pipeline_registers.registers[15][8] ),
    .S0(net611),
    .S1(net587),
    .X(_02401_));
 sky130_fd_sc_hd__or2_1 _12076_ (.A(net473),
    .B(_02401_),
    .X(_02402_));
 sky130_fd_sc_hd__o21a_1 _12077_ (.A1(net577),
    .A2(_02400_),
    .B1(net571),
    .X(_02403_));
 sky130_fd_sc_hd__a221o_1 _12078_ (.A1(net468),
    .A2(_02399_),
    .B1(_02402_),
    .B2(_02403_),
    .C1(net567),
    .X(_02404_));
 sky130_fd_sc_hd__mux2_1 _12079_ (.A0(\core_pipeline.pipeline_registers.registers[30][8] ),
    .A1(\core_pipeline.pipeline_registers.registers[31][8] ),
    .S(net608),
    .X(_02405_));
 sky130_fd_sc_hd__and2_1 _12080_ (.A(net587),
    .B(_02405_),
    .X(_02406_));
 sky130_fd_sc_hd__mux2_1 _12081_ (.A0(\core_pipeline.pipeline_registers.registers[28][8] ),
    .A1(\core_pipeline.pipeline_registers.registers[29][8] ),
    .S(net607),
    .X(_02407_));
 sky130_fd_sc_hd__a21o_1 _12082_ (.A1(net482),
    .A2(_02407_),
    .B1(net473),
    .X(_02408_));
 sky130_fd_sc_hd__mux2_1 _12083_ (.A0(\core_pipeline.pipeline_registers.registers[26][8] ),
    .A1(\core_pipeline.pipeline_registers.registers[27][8] ),
    .S(net607),
    .X(_02409_));
 sky130_fd_sc_hd__and2_1 _12084_ (.A(net586),
    .B(_02409_),
    .X(_02410_));
 sky130_fd_sc_hd__mux2_1 _12085_ (.A0(\core_pipeline.pipeline_registers.registers[24][8] ),
    .A1(\core_pipeline.pipeline_registers.registers[25][8] ),
    .S(net607),
    .X(_02411_));
 sky130_fd_sc_hd__a21o_1 _12086_ (.A1(net482),
    .A2(_02411_),
    .B1(net577),
    .X(_02412_));
 sky130_fd_sc_hd__o221a_1 _12087_ (.A1(_02406_),
    .A2(_02408_),
    .B1(_02410_),
    .B2(_02412_),
    .C1(net571),
    .X(_02413_));
 sky130_fd_sc_hd__mux2_1 _12088_ (.A0(_02397_),
    .A1(_02398_),
    .S(net473),
    .X(_02414_));
 sky130_fd_sc_hd__a211o_1 _12089_ (.A1(net468),
    .A2(_02414_),
    .B1(_02413_),
    .C1(net467),
    .X(_02415_));
 sky130_fd_sc_hd__and3_1 _12090_ (.A(net144),
    .B(_02404_),
    .C(_02415_),
    .X(_02416_));
 sky130_fd_sc_hd__a21o_1 _12091_ (.A1(\core_pipeline.decode_to_execute_rs1_data[8] ),
    .A2(net124),
    .B1(_02416_),
    .X(_01929_));
 sky130_fd_sc_hd__mux4_1 _12092_ (.A0(\core_pipeline.pipeline_registers.registers[4][9] ),
    .A1(\core_pipeline.pipeline_registers.registers[5][9] ),
    .A2(\core_pipeline.pipeline_registers.registers[6][9] ),
    .A3(\core_pipeline.pipeline_registers.registers[7][9] ),
    .S0(net606),
    .S1(net584),
    .X(_02417_));
 sky130_fd_sc_hd__mux4_1 _12093_ (.A0(\core_pipeline.pipeline_registers.registers[0][9] ),
    .A1(\core_pipeline.pipeline_registers.registers[1][9] ),
    .A2(\core_pipeline.pipeline_registers.registers[2][9] ),
    .A3(\core_pipeline.pipeline_registers.registers[3][9] ),
    .S0(net606),
    .S1(net584),
    .X(_02418_));
 sky130_fd_sc_hd__mux4_1 _12094_ (.A0(\core_pipeline.pipeline_registers.registers[20][9] ),
    .A1(\core_pipeline.pipeline_registers.registers[21][9] ),
    .A2(\core_pipeline.pipeline_registers.registers[22][9] ),
    .A3(\core_pipeline.pipeline_registers.registers[23][9] ),
    .S0(net605),
    .S1(net585),
    .X(_02419_));
 sky130_fd_sc_hd__mux4_1 _12095_ (.A0(\core_pipeline.pipeline_registers.registers[16][9] ),
    .A1(\core_pipeline.pipeline_registers.registers[17][9] ),
    .A2(\core_pipeline.pipeline_registers.registers[18][9] ),
    .A3(\core_pipeline.pipeline_registers.registers[19][9] ),
    .S0(net605),
    .S1(net585),
    .X(_02420_));
 sky130_fd_sc_hd__mux2_1 _12096_ (.A0(_02417_),
    .A1(_02418_),
    .S(net474),
    .X(_02421_));
 sky130_fd_sc_hd__mux4_1 _12097_ (.A0(\core_pipeline.pipeline_registers.registers[8][9] ),
    .A1(\core_pipeline.pipeline_registers.registers[9][9] ),
    .A2(\core_pipeline.pipeline_registers.registers[10][9] ),
    .A3(\core_pipeline.pipeline_registers.registers[11][9] ),
    .S0(net606),
    .S1(net584),
    .X(_02422_));
 sky130_fd_sc_hd__mux4_1 _12098_ (.A0(\core_pipeline.pipeline_registers.registers[12][9] ),
    .A1(\core_pipeline.pipeline_registers.registers[13][9] ),
    .A2(\core_pipeline.pipeline_registers.registers[14][9] ),
    .A3(\core_pipeline.pipeline_registers.registers[15][9] ),
    .S0(net606),
    .S1(net584),
    .X(_02423_));
 sky130_fd_sc_hd__or2_1 _12099_ (.A(net472),
    .B(_02423_),
    .X(_02424_));
 sky130_fd_sc_hd__o21a_1 _12100_ (.A1(net576),
    .A2(_02422_),
    .B1(net570),
    .X(_02425_));
 sky130_fd_sc_hd__a221o_1 _12101_ (.A1(net468),
    .A2(_02421_),
    .B1(_02424_),
    .B2(_02425_),
    .C1(net567),
    .X(_02426_));
 sky130_fd_sc_hd__mux2_1 _12102_ (.A0(\core_pipeline.pipeline_registers.registers[30][9] ),
    .A1(\core_pipeline.pipeline_registers.registers[31][9] ),
    .S(net609),
    .X(_02427_));
 sky130_fd_sc_hd__and2_1 _12103_ (.A(net585),
    .B(_02427_),
    .X(_02428_));
 sky130_fd_sc_hd__mux2_1 _12104_ (.A0(\core_pipeline.pipeline_registers.registers[28][9] ),
    .A1(\core_pipeline.pipeline_registers.registers[29][9] ),
    .S(net605),
    .X(_02429_));
 sky130_fd_sc_hd__a21o_1 _12105_ (.A1(net483),
    .A2(_02429_),
    .B1(net472),
    .X(_02430_));
 sky130_fd_sc_hd__mux2_1 _12106_ (.A0(\core_pipeline.pipeline_registers.registers[26][9] ),
    .A1(\core_pipeline.pipeline_registers.registers[27][9] ),
    .S(net605),
    .X(_02431_));
 sky130_fd_sc_hd__and2_1 _12107_ (.A(net585),
    .B(_02431_),
    .X(_02432_));
 sky130_fd_sc_hd__mux2_1 _12108_ (.A0(\core_pipeline.pipeline_registers.registers[24][9] ),
    .A1(\core_pipeline.pipeline_registers.registers[25][9] ),
    .S(net605),
    .X(_02433_));
 sky130_fd_sc_hd__a21o_1 _12109_ (.A1(net482),
    .A2(_02433_),
    .B1(net576),
    .X(_02434_));
 sky130_fd_sc_hd__o221a_1 _12110_ (.A1(_02428_),
    .A2(_02430_),
    .B1(_02432_),
    .B2(_02434_),
    .C1(net570),
    .X(_02435_));
 sky130_fd_sc_hd__mux2_1 _12111_ (.A0(_02419_),
    .A1(_02420_),
    .S(net472),
    .X(_02436_));
 sky130_fd_sc_hd__a211o_1 _12112_ (.A1(net468),
    .A2(_02436_),
    .B1(_02435_),
    .C1(net467),
    .X(_02437_));
 sky130_fd_sc_hd__and3_1 _12113_ (.A(net144),
    .B(_02426_),
    .C(_02437_),
    .X(_02438_));
 sky130_fd_sc_hd__a21o_1 _12114_ (.A1(\core_pipeline.decode_to_execute_rs1_data[9] ),
    .A2(net121),
    .B1(_02438_),
    .X(_01930_));
 sky130_fd_sc_hd__mux4_1 _12115_ (.A0(\core_pipeline.pipeline_registers.registers[4][10] ),
    .A1(\core_pipeline.pipeline_registers.registers[5][10] ),
    .A2(\core_pipeline.pipeline_registers.registers[6][10] ),
    .A3(\core_pipeline.pipeline_registers.registers[7][10] ),
    .S0(net612),
    .S1(net590),
    .X(_02439_));
 sky130_fd_sc_hd__mux4_1 _12116_ (.A0(\core_pipeline.pipeline_registers.registers[0][10] ),
    .A1(\core_pipeline.pipeline_registers.registers[1][10] ),
    .A2(\core_pipeline.pipeline_registers.registers[2][10] ),
    .A3(\core_pipeline.pipeline_registers.registers[3][10] ),
    .S0(net614),
    .S1(net590),
    .X(_02440_));
 sky130_fd_sc_hd__mux4_1 _12117_ (.A0(\core_pipeline.pipeline_registers.registers[20][10] ),
    .A1(\core_pipeline.pipeline_registers.registers[21][10] ),
    .A2(\core_pipeline.pipeline_registers.registers[22][10] ),
    .A3(\core_pipeline.pipeline_registers.registers[23][10] ),
    .S0(net606),
    .S1(net584),
    .X(_02441_));
 sky130_fd_sc_hd__mux4_1 _12118_ (.A0(\core_pipeline.pipeline_registers.registers[16][10] ),
    .A1(\core_pipeline.pipeline_registers.registers[17][10] ),
    .A2(\core_pipeline.pipeline_registers.registers[18][10] ),
    .A3(\core_pipeline.pipeline_registers.registers[19][10] ),
    .S0(net606),
    .S1(net584),
    .X(_02442_));
 sky130_fd_sc_hd__mux2_1 _12119_ (.A0(_02439_),
    .A1(_02440_),
    .S(net475),
    .X(_02443_));
 sky130_fd_sc_hd__mux4_1 _12120_ (.A0(\core_pipeline.pipeline_registers.registers[8][10] ),
    .A1(\core_pipeline.pipeline_registers.registers[9][10] ),
    .A2(\core_pipeline.pipeline_registers.registers[10][10] ),
    .A3(\core_pipeline.pipeline_registers.registers[11][10] ),
    .S0(net612),
    .S1(net590),
    .X(_02444_));
 sky130_fd_sc_hd__mux4_1 _12121_ (.A0(\core_pipeline.pipeline_registers.registers[12][10] ),
    .A1(\core_pipeline.pipeline_registers.registers[13][10] ),
    .A2(\core_pipeline.pipeline_registers.registers[14][10] ),
    .A3(\core_pipeline.pipeline_registers.registers[15][10] ),
    .S0(net612),
    .S1(net590),
    .X(_02445_));
 sky130_fd_sc_hd__or2_1 _12122_ (.A(net475),
    .B(_02445_),
    .X(_02446_));
 sky130_fd_sc_hd__o21a_1 _12123_ (.A1(net578),
    .A2(_02444_),
    .B1(net572),
    .X(_02447_));
 sky130_fd_sc_hd__a221o_1 _12124_ (.A1(net469),
    .A2(_02443_),
    .B1(_02446_),
    .B2(_02447_),
    .C1(net567),
    .X(_02448_));
 sky130_fd_sc_hd__mux2_1 _12125_ (.A0(\core_pipeline.pipeline_registers.registers[30][10] ),
    .A1(\core_pipeline.pipeline_registers.registers[31][10] ),
    .S(net605),
    .X(_02449_));
 sky130_fd_sc_hd__and2_1 _12126_ (.A(net585),
    .B(_02449_),
    .X(_02450_));
 sky130_fd_sc_hd__mux2_1 _12127_ (.A0(\core_pipeline.pipeline_registers.registers[28][10] ),
    .A1(\core_pipeline.pipeline_registers.registers[29][10] ),
    .S(net605),
    .X(_02451_));
 sky130_fd_sc_hd__a21o_1 _12128_ (.A1(net483),
    .A2(_02451_),
    .B1(net475),
    .X(_02452_));
 sky130_fd_sc_hd__mux2_1 _12129_ (.A0(\core_pipeline.pipeline_registers.registers[26][10] ),
    .A1(\core_pipeline.pipeline_registers.registers[27][10] ),
    .S(net605),
    .X(_02453_));
 sky130_fd_sc_hd__and2_1 _12130_ (.A(net585),
    .B(_02453_),
    .X(_02454_));
 sky130_fd_sc_hd__mux2_1 _12131_ (.A0(\core_pipeline.pipeline_registers.registers[24][10] ),
    .A1(\core_pipeline.pipeline_registers.registers[25][10] ),
    .S(net605),
    .X(_02455_));
 sky130_fd_sc_hd__a21o_1 _12132_ (.A1(net483),
    .A2(_02455_),
    .B1(net576),
    .X(_02456_));
 sky130_fd_sc_hd__o221a_1 _12133_ (.A1(_02450_),
    .A2(_02452_),
    .B1(_02454_),
    .B2(_02456_),
    .C1(net570),
    .X(_02457_));
 sky130_fd_sc_hd__mux2_1 _12134_ (.A0(_02441_),
    .A1(_02442_),
    .S(net475),
    .X(_02458_));
 sky130_fd_sc_hd__a211o_1 _12135_ (.A1(net469),
    .A2(_02458_),
    .B1(_02457_),
    .C1(net467),
    .X(_02459_));
 sky130_fd_sc_hd__and3_1 _12136_ (.A(net139),
    .B(_02448_),
    .C(_02459_),
    .X(_02460_));
 sky130_fd_sc_hd__a21o_1 _12137_ (.A1(\core_pipeline.decode_to_execute_rs1_data[10] ),
    .A2(net122),
    .B1(_02460_),
    .X(_01931_));
 sky130_fd_sc_hd__mux4_1 _12138_ (.A0(\core_pipeline.pipeline_registers.registers[4][11] ),
    .A1(\core_pipeline.pipeline_registers.registers[5][11] ),
    .A2(\core_pipeline.pipeline_registers.registers[6][11] ),
    .A3(\core_pipeline.pipeline_registers.registers[7][11] ),
    .S0(net606),
    .S1(net584),
    .X(_02461_));
 sky130_fd_sc_hd__mux4_1 _12139_ (.A0(\core_pipeline.pipeline_registers.registers[0][11] ),
    .A1(\core_pipeline.pipeline_registers.registers[1][11] ),
    .A2(\core_pipeline.pipeline_registers.registers[2][11] ),
    .A3(\core_pipeline.pipeline_registers.registers[3][11] ),
    .S0(net606),
    .S1(net584),
    .X(_02462_));
 sky130_fd_sc_hd__mux4_1 _12140_ (.A0(\core_pipeline.pipeline_registers.registers[20][11] ),
    .A1(\core_pipeline.pipeline_registers.registers[21][11] ),
    .A2(\core_pipeline.pipeline_registers.registers[22][11] ),
    .A3(\core_pipeline.pipeline_registers.registers[23][11] ),
    .S0(net604),
    .S1(net582),
    .X(_02463_));
 sky130_fd_sc_hd__mux4_1 _12141_ (.A0(\core_pipeline.pipeline_registers.registers[16][11] ),
    .A1(\core_pipeline.pipeline_registers.registers[17][11] ),
    .A2(\core_pipeline.pipeline_registers.registers[18][11] ),
    .A3(\core_pipeline.pipeline_registers.registers[19][11] ),
    .S0(net604),
    .S1(net583),
    .X(_02464_));
 sky130_fd_sc_hd__mux2_1 _12142_ (.A0(_02461_),
    .A1(_02462_),
    .S(net474),
    .X(_02465_));
 sky130_fd_sc_hd__mux4_1 _12143_ (.A0(\core_pipeline.pipeline_registers.registers[8][11] ),
    .A1(\core_pipeline.pipeline_registers.registers[9][11] ),
    .A2(\core_pipeline.pipeline_registers.registers[10][11] ),
    .A3(\core_pipeline.pipeline_registers.registers[11][11] ),
    .S0(net603),
    .S1(net582),
    .X(_02466_));
 sky130_fd_sc_hd__mux4_1 _12144_ (.A0(\core_pipeline.pipeline_registers.registers[12][11] ),
    .A1(\core_pipeline.pipeline_registers.registers[13][11] ),
    .A2(\core_pipeline.pipeline_registers.registers[14][11] ),
    .A3(\core_pipeline.pipeline_registers.registers[15][11] ),
    .S0(net603),
    .S1(net582),
    .X(_02467_));
 sky130_fd_sc_hd__or2_1 _12145_ (.A(net474),
    .B(_02467_),
    .X(_02468_));
 sky130_fd_sc_hd__o21a_1 _12146_ (.A1(net576),
    .A2(_02466_),
    .B1(net570),
    .X(_02469_));
 sky130_fd_sc_hd__a221o_2 _12147_ (.A1(net468),
    .A2(_02465_),
    .B1(_02468_),
    .B2(_02469_),
    .C1(net567),
    .X(_02470_));
 sky130_fd_sc_hd__mux2_1 _12148_ (.A0(\core_pipeline.pipeline_registers.registers[30][11] ),
    .A1(\core_pipeline.pipeline_registers.registers[31][11] ),
    .S(net607),
    .X(_02471_));
 sky130_fd_sc_hd__and2_1 _12149_ (.A(net586),
    .B(_02471_),
    .X(_02472_));
 sky130_fd_sc_hd__mux2_1 _12150_ (.A0(\core_pipeline.pipeline_registers.registers[28][11] ),
    .A1(\core_pipeline.pipeline_registers.registers[29][11] ),
    .S(net607),
    .X(_02473_));
 sky130_fd_sc_hd__a21o_1 _12151_ (.A1(net482),
    .A2(_02473_),
    .B1(net473),
    .X(_02474_));
 sky130_fd_sc_hd__mux2_1 _12152_ (.A0(\core_pipeline.pipeline_registers.registers[26][11] ),
    .A1(\core_pipeline.pipeline_registers.registers[27][11] ),
    .S(net607),
    .X(_02475_));
 sky130_fd_sc_hd__and2_1 _12153_ (.A(net586),
    .B(_02475_),
    .X(_02476_));
 sky130_fd_sc_hd__mux2_1 _12154_ (.A0(\core_pipeline.pipeline_registers.registers[24][11] ),
    .A1(\core_pipeline.pipeline_registers.registers[25][11] ),
    .S(net603),
    .X(_02477_));
 sky130_fd_sc_hd__a21o_1 _12155_ (.A1(net482),
    .A2(_02477_),
    .B1(net576),
    .X(_02478_));
 sky130_fd_sc_hd__o221a_1 _12156_ (.A1(_02472_),
    .A2(_02474_),
    .B1(_02476_),
    .B2(_02478_),
    .C1(net571),
    .X(_02479_));
 sky130_fd_sc_hd__mux2_1 _12157_ (.A0(_02463_),
    .A1(_02464_),
    .S(net472),
    .X(_02480_));
 sky130_fd_sc_hd__a211o_1 _12158_ (.A1(net468),
    .A2(_02480_),
    .B1(_02479_),
    .C1(net467),
    .X(_02481_));
 sky130_fd_sc_hd__and3_1 _12159_ (.A(net144),
    .B(_02470_),
    .C(_02481_),
    .X(_02482_));
 sky130_fd_sc_hd__a21o_1 _12160_ (.A1(\core_pipeline.decode_to_execute_rs1_data[11] ),
    .A2(net121),
    .B1(_02482_),
    .X(_01932_));
 sky130_fd_sc_hd__mux4_1 _12161_ (.A0(\core_pipeline.pipeline_registers.registers[4][12] ),
    .A1(\core_pipeline.pipeline_registers.registers[5][12] ),
    .A2(\core_pipeline.pipeline_registers.registers[6][12] ),
    .A3(\core_pipeline.pipeline_registers.registers[7][12] ),
    .S0(net609),
    .S1(net586),
    .X(_02483_));
 sky130_fd_sc_hd__mux4_1 _12162_ (.A0(\core_pipeline.pipeline_registers.registers[0][12] ),
    .A1(\core_pipeline.pipeline_registers.registers[1][12] ),
    .A2(\core_pipeline.pipeline_registers.registers[2][12] ),
    .A3(\core_pipeline.pipeline_registers.registers[3][12] ),
    .S0(net609),
    .S1(net588),
    .X(_02484_));
 sky130_fd_sc_hd__mux4_1 _12163_ (.A0(\core_pipeline.pipeline_registers.registers[20][12] ),
    .A1(\core_pipeline.pipeline_registers.registers[21][12] ),
    .A2(\core_pipeline.pipeline_registers.registers[22][12] ),
    .A3(\core_pipeline.pipeline_registers.registers[23][12] ),
    .S0(net609),
    .S1(net588),
    .X(_02485_));
 sky130_fd_sc_hd__mux4_1 _12164_ (.A0(\core_pipeline.pipeline_registers.registers[16][12] ),
    .A1(\core_pipeline.pipeline_registers.registers[17][12] ),
    .A2(\core_pipeline.pipeline_registers.registers[18][12] ),
    .A3(\core_pipeline.pipeline_registers.registers[19][12] ),
    .S0(net609),
    .S1(net588),
    .X(_02486_));
 sky130_fd_sc_hd__mux2_1 _12165_ (.A0(_02483_),
    .A1(_02484_),
    .S(net474),
    .X(_02487_));
 sky130_fd_sc_hd__mux4_1 _12166_ (.A0(\core_pipeline.pipeline_registers.registers[8][12] ),
    .A1(\core_pipeline.pipeline_registers.registers[9][12] ),
    .A2(\core_pipeline.pipeline_registers.registers[10][12] ),
    .A3(\core_pipeline.pipeline_registers.registers[11][12] ),
    .S0(net605),
    .S1(net585),
    .X(_02488_));
 sky130_fd_sc_hd__mux4_1 _12167_ (.A0(\core_pipeline.pipeline_registers.registers[12][12] ),
    .A1(\core_pipeline.pipeline_registers.registers[13][12] ),
    .A2(\core_pipeline.pipeline_registers.registers[14][12] ),
    .A3(\core_pipeline.pipeline_registers.registers[15][12] ),
    .S0(net603),
    .S1(net583),
    .X(_02489_));
 sky130_fd_sc_hd__or2_1 _12168_ (.A(net474),
    .B(_02489_),
    .X(_02490_));
 sky130_fd_sc_hd__o21a_1 _12169_ (.A1(net576),
    .A2(_02488_),
    .B1(net570),
    .X(_02491_));
 sky130_fd_sc_hd__a221o_1 _12170_ (.A1(net469),
    .A2(_02487_),
    .B1(_02490_),
    .B2(_02491_),
    .C1(net567),
    .X(_02492_));
 sky130_fd_sc_hd__mux2_1 _12171_ (.A0(\core_pipeline.pipeline_registers.registers[30][12] ),
    .A1(\core_pipeline.pipeline_registers.registers[31][12] ),
    .S(net609),
    .X(_02493_));
 sky130_fd_sc_hd__and2_1 _12172_ (.A(net588),
    .B(_02493_),
    .X(_02494_));
 sky130_fd_sc_hd__mux2_1 _12173_ (.A0(\core_pipeline.pipeline_registers.registers[28][12] ),
    .A1(\core_pipeline.pipeline_registers.registers[29][12] ),
    .S(net609),
    .X(_02495_));
 sky130_fd_sc_hd__a21o_1 _12174_ (.A1(net483),
    .A2(_02495_),
    .B1(net476),
    .X(_02496_));
 sky130_fd_sc_hd__mux2_1 _12175_ (.A0(\core_pipeline.pipeline_registers.registers[26][12] ),
    .A1(\core_pipeline.pipeline_registers.registers[27][12] ),
    .S(net609),
    .X(_02497_));
 sky130_fd_sc_hd__and2_1 _12176_ (.A(net588),
    .B(_02497_),
    .X(_02498_));
 sky130_fd_sc_hd__mux2_1 _12177_ (.A0(\core_pipeline.pipeline_registers.registers[24][12] ),
    .A1(\core_pipeline.pipeline_registers.registers[25][12] ),
    .S(net609),
    .X(_02499_));
 sky130_fd_sc_hd__a21o_1 _12178_ (.A1(net483),
    .A2(_02499_),
    .B1(net577),
    .X(_02500_));
 sky130_fd_sc_hd__o221a_1 _12179_ (.A1(_02494_),
    .A2(_02496_),
    .B1(_02498_),
    .B2(_02500_),
    .C1(net571),
    .X(_02501_));
 sky130_fd_sc_hd__mux2_1 _12180_ (.A0(_02485_),
    .A1(_02486_),
    .S(net476),
    .X(_02502_));
 sky130_fd_sc_hd__a211o_1 _12181_ (.A1(net469),
    .A2(_02502_),
    .B1(_02501_),
    .C1(net467),
    .X(_02503_));
 sky130_fd_sc_hd__and3_1 _12182_ (.A(net144),
    .B(_02492_),
    .C(_02503_),
    .X(_02504_));
 sky130_fd_sc_hd__a21o_1 _12183_ (.A1(\core_pipeline.decode_to_execute_rs1_data[12] ),
    .A2(net121),
    .B1(_02504_),
    .X(_01933_));
 sky130_fd_sc_hd__mux4_1 _12184_ (.A0(\core_pipeline.pipeline_registers.registers[4][13] ),
    .A1(\core_pipeline.pipeline_registers.registers[5][13] ),
    .A2(\core_pipeline.pipeline_registers.registers[6][13] ),
    .A3(\core_pipeline.pipeline_registers.registers[7][13] ),
    .S0(net612),
    .S1(net590),
    .X(_02505_));
 sky130_fd_sc_hd__mux4_1 _12185_ (.A0(\core_pipeline.pipeline_registers.registers[0][13] ),
    .A1(\core_pipeline.pipeline_registers.registers[1][13] ),
    .A2(\core_pipeline.pipeline_registers.registers[2][13] ),
    .A3(\core_pipeline.pipeline_registers.registers[3][13] ),
    .S0(net612),
    .S1(net590),
    .X(_02506_));
 sky130_fd_sc_hd__mux4_1 _12186_ (.A0(\core_pipeline.pipeline_registers.registers[20][13] ),
    .A1(\core_pipeline.pipeline_registers.registers[21][13] ),
    .A2(\core_pipeline.pipeline_registers.registers[22][13] ),
    .A3(\core_pipeline.pipeline_registers.registers[23][13] ),
    .S0(net606),
    .S1(net584),
    .X(_02507_));
 sky130_fd_sc_hd__mux4_1 _12187_ (.A0(\core_pipeline.pipeline_registers.registers[16][13] ),
    .A1(\core_pipeline.pipeline_registers.registers[17][13] ),
    .A2(\core_pipeline.pipeline_registers.registers[18][13] ),
    .A3(\core_pipeline.pipeline_registers.registers[19][13] ),
    .S0(net612),
    .S1(net584),
    .X(_02508_));
 sky130_fd_sc_hd__mux2_1 _12188_ (.A0(_02505_),
    .A1(_02506_),
    .S(net475),
    .X(_02509_));
 sky130_fd_sc_hd__mux4_1 _12189_ (.A0(\core_pipeline.pipeline_registers.registers[8][13] ),
    .A1(\core_pipeline.pipeline_registers.registers[9][13] ),
    .A2(\core_pipeline.pipeline_registers.registers[10][13] ),
    .A3(\core_pipeline.pipeline_registers.registers[11][13] ),
    .S0(net606),
    .S1(net585),
    .X(_02510_));
 sky130_fd_sc_hd__mux4_1 _12190_ (.A0(\core_pipeline.pipeline_registers.registers[12][13] ),
    .A1(\core_pipeline.pipeline_registers.registers[13][13] ),
    .A2(\core_pipeline.pipeline_registers.registers[14][13] ),
    .A3(\core_pipeline.pipeline_registers.registers[15][13] ),
    .S0(net612),
    .S1(net584),
    .X(_02511_));
 sky130_fd_sc_hd__or2_1 _12191_ (.A(net475),
    .B(_02511_),
    .X(_02512_));
 sky130_fd_sc_hd__o21a_1 _12192_ (.A1(net576),
    .A2(_02510_),
    .B1(net570),
    .X(_02513_));
 sky130_fd_sc_hd__a221o_1 _12193_ (.A1(net469),
    .A2(_02509_),
    .B1(_02512_),
    .B2(_02513_),
    .C1(net567),
    .X(_02514_));
 sky130_fd_sc_hd__mux2_1 _12194_ (.A0(\core_pipeline.pipeline_registers.registers[30][13] ),
    .A1(\core_pipeline.pipeline_registers.registers[31][13] ),
    .S(net613),
    .X(_02515_));
 sky130_fd_sc_hd__and2_1 _12195_ (.A(net585),
    .B(_02515_),
    .X(_02516_));
 sky130_fd_sc_hd__mux2_1 _12196_ (.A0(\core_pipeline.pipeline_registers.registers[28][13] ),
    .A1(\core_pipeline.pipeline_registers.registers[29][13] ),
    .S(net613),
    .X(_02517_));
 sky130_fd_sc_hd__a21o_1 _12197_ (.A1(net483),
    .A2(_02517_),
    .B1(net475),
    .X(_02518_));
 sky130_fd_sc_hd__mux2_1 _12198_ (.A0(\core_pipeline.pipeline_registers.registers[26][13] ),
    .A1(\core_pipeline.pipeline_registers.registers[27][13] ),
    .S(net605),
    .X(_02519_));
 sky130_fd_sc_hd__and2_1 _12199_ (.A(net585),
    .B(_02519_),
    .X(_02520_));
 sky130_fd_sc_hd__mux2_1 _12200_ (.A0(\core_pipeline.pipeline_registers.registers[24][13] ),
    .A1(\core_pipeline.pipeline_registers.registers[25][13] ),
    .S(net613),
    .X(_02521_));
 sky130_fd_sc_hd__a21o_1 _12201_ (.A1(net483),
    .A2(_02521_),
    .B1(net576),
    .X(_02522_));
 sky130_fd_sc_hd__o221a_1 _12202_ (.A1(_02516_),
    .A2(_02518_),
    .B1(_02520_),
    .B2(_02522_),
    .C1(net570),
    .X(_02523_));
 sky130_fd_sc_hd__mux2_1 _12203_ (.A0(_02507_),
    .A1(_02508_),
    .S(net475),
    .X(_02524_));
 sky130_fd_sc_hd__a211o_1 _12204_ (.A1(net469),
    .A2(_02524_),
    .B1(_02523_),
    .C1(net467),
    .X(_02525_));
 sky130_fd_sc_hd__and3_1 _12205_ (.A(net139),
    .B(_02514_),
    .C(_02525_),
    .X(_02526_));
 sky130_fd_sc_hd__a21o_1 _12206_ (.A1(\core_pipeline.decode_to_execute_rs1_data[13] ),
    .A2(net122),
    .B1(_02526_),
    .X(_01934_));
 sky130_fd_sc_hd__mux4_1 _12207_ (.A0(\core_pipeline.pipeline_registers.registers[4][14] ),
    .A1(\core_pipeline.pipeline_registers.registers[5][14] ),
    .A2(\core_pipeline.pipeline_registers.registers[6][14] ),
    .A3(\core_pipeline.pipeline_registers.registers[7][14] ),
    .S0(net612),
    .S1(net590),
    .X(_02527_));
 sky130_fd_sc_hd__mux4_1 _12208_ (.A0(\core_pipeline.pipeline_registers.registers[0][14] ),
    .A1(\core_pipeline.pipeline_registers.registers[1][14] ),
    .A2(\core_pipeline.pipeline_registers.registers[2][14] ),
    .A3(\core_pipeline.pipeline_registers.registers[3][14] ),
    .S0(net614),
    .S1(net590),
    .X(_02528_));
 sky130_fd_sc_hd__mux4_1 _12209_ (.A0(\core_pipeline.pipeline_registers.registers[20][14] ),
    .A1(\core_pipeline.pipeline_registers.registers[21][14] ),
    .A2(\core_pipeline.pipeline_registers.registers[22][14] ),
    .A3(\core_pipeline.pipeline_registers.registers[23][14] ),
    .S0(net606),
    .S1(net584),
    .X(_02529_));
 sky130_fd_sc_hd__mux4_1 _12210_ (.A0(\core_pipeline.pipeline_registers.registers[16][14] ),
    .A1(\core_pipeline.pipeline_registers.registers[17][14] ),
    .A2(\core_pipeline.pipeline_registers.registers[18][14] ),
    .A3(\core_pipeline.pipeline_registers.registers[19][14] ),
    .S0(net606),
    .S1(net584),
    .X(_02530_));
 sky130_fd_sc_hd__mux2_1 _12211_ (.A0(_02527_),
    .A1(_02528_),
    .S(net475),
    .X(_02531_));
 sky130_fd_sc_hd__mux4_1 _12212_ (.A0(\core_pipeline.pipeline_registers.registers[8][14] ),
    .A1(\core_pipeline.pipeline_registers.registers[9][14] ),
    .A2(\core_pipeline.pipeline_registers.registers[10][14] ),
    .A3(\core_pipeline.pipeline_registers.registers[11][14] ),
    .S0(net612),
    .S1(net590),
    .X(_02532_));
 sky130_fd_sc_hd__mux4_1 _12213_ (.A0(\core_pipeline.pipeline_registers.registers[12][14] ),
    .A1(\core_pipeline.pipeline_registers.registers[13][14] ),
    .A2(\core_pipeline.pipeline_registers.registers[14][14] ),
    .A3(\core_pipeline.pipeline_registers.registers[15][14] ),
    .S0(net612),
    .S1(net590),
    .X(_02533_));
 sky130_fd_sc_hd__or2_1 _12214_ (.A(net476),
    .B(_02533_),
    .X(_02534_));
 sky130_fd_sc_hd__o21a_1 _12215_ (.A1(net578),
    .A2(_02532_),
    .B1(net572),
    .X(_02535_));
 sky130_fd_sc_hd__a221o_1 _12216_ (.A1(net469),
    .A2(_02531_),
    .B1(_02534_),
    .B2(_02535_),
    .C1(net569),
    .X(_02536_));
 sky130_fd_sc_hd__mux2_1 _12217_ (.A0(\core_pipeline.pipeline_registers.registers[30][14] ),
    .A1(\core_pipeline.pipeline_registers.registers[31][14] ),
    .S(net605),
    .X(_02537_));
 sky130_fd_sc_hd__and2_1 _12218_ (.A(net585),
    .B(_02537_),
    .X(_02538_));
 sky130_fd_sc_hd__mux2_1 _12219_ (.A0(\core_pipeline.pipeline_registers.registers[28][14] ),
    .A1(\core_pipeline.pipeline_registers.registers[29][14] ),
    .S(net605),
    .X(_02539_));
 sky130_fd_sc_hd__a21o_1 _12220_ (.A1(net483),
    .A2(_02539_),
    .B1(net474),
    .X(_02540_));
 sky130_fd_sc_hd__mux2_1 _12221_ (.A0(\core_pipeline.pipeline_registers.registers[26][14] ),
    .A1(\core_pipeline.pipeline_registers.registers[27][14] ),
    .S(net605),
    .X(_02541_));
 sky130_fd_sc_hd__and2_1 _12222_ (.A(net585),
    .B(_02541_),
    .X(_02542_));
 sky130_fd_sc_hd__mux2_1 _12223_ (.A0(\core_pipeline.pipeline_registers.registers[24][14] ),
    .A1(\core_pipeline.pipeline_registers.registers[25][14] ),
    .S(net605),
    .X(_02543_));
 sky130_fd_sc_hd__a21o_1 _12224_ (.A1(net483),
    .A2(_02543_),
    .B1(net576),
    .X(_02544_));
 sky130_fd_sc_hd__o221a_1 _12225_ (.A1(_02538_),
    .A2(_02540_),
    .B1(_02542_),
    .B2(_02544_),
    .C1(net570),
    .X(_02545_));
 sky130_fd_sc_hd__mux2_1 _12226_ (.A0(_02529_),
    .A1(_02530_),
    .S(net472),
    .X(_02546_));
 sky130_fd_sc_hd__a211o_2 _12227_ (.A1(net468),
    .A2(_02546_),
    .B1(_02545_),
    .C1(net467),
    .X(_02547_));
 sky130_fd_sc_hd__and3_1 _12228_ (.A(net140),
    .B(_02536_),
    .C(_02547_),
    .X(_02548_));
 sky130_fd_sc_hd__a21o_1 _12229_ (.A1(\core_pipeline.decode_to_execute_rs1_data[14] ),
    .A2(net122),
    .B1(_02548_),
    .X(_01935_));
 sky130_fd_sc_hd__mux4_1 _12230_ (.A0(\core_pipeline.pipeline_registers.registers[4][15] ),
    .A1(\core_pipeline.pipeline_registers.registers[5][15] ),
    .A2(\core_pipeline.pipeline_registers.registers[6][15] ),
    .A3(\core_pipeline.pipeline_registers.registers[7][15] ),
    .S0(net613),
    .S1(net591),
    .X(_02549_));
 sky130_fd_sc_hd__mux4_1 _12231_ (.A0(\core_pipeline.pipeline_registers.registers[0][15] ),
    .A1(\core_pipeline.pipeline_registers.registers[1][15] ),
    .A2(\core_pipeline.pipeline_registers.registers[2][15] ),
    .A3(\core_pipeline.pipeline_registers.registers[3][15] ),
    .S0(net613),
    .S1(net591),
    .X(_02550_));
 sky130_fd_sc_hd__mux4_1 _12232_ (.A0(\core_pipeline.pipeline_registers.registers[20][15] ),
    .A1(\core_pipeline.pipeline_registers.registers[21][15] ),
    .A2(\core_pipeline.pipeline_registers.registers[22][15] ),
    .A3(\core_pipeline.pipeline_registers.registers[23][15] ),
    .S0(net613),
    .S1(net590),
    .X(_02551_));
 sky130_fd_sc_hd__mux4_1 _12233_ (.A0(\core_pipeline.pipeline_registers.registers[16][15] ),
    .A1(\core_pipeline.pipeline_registers.registers[17][15] ),
    .A2(\core_pipeline.pipeline_registers.registers[18][15] ),
    .A3(\core_pipeline.pipeline_registers.registers[19][15] ),
    .S0(net613),
    .S1(net591),
    .X(_02552_));
 sky130_fd_sc_hd__mux2_1 _12234_ (.A0(_02549_),
    .A1(_02550_),
    .S(net476),
    .X(_02553_));
 sky130_fd_sc_hd__mux4_1 _12235_ (.A0(\core_pipeline.pipeline_registers.registers[8][15] ),
    .A1(\core_pipeline.pipeline_registers.registers[9][15] ),
    .A2(\core_pipeline.pipeline_registers.registers[10][15] ),
    .A3(\core_pipeline.pipeline_registers.registers[11][15] ),
    .S0(net613),
    .S1(net591),
    .X(_02554_));
 sky130_fd_sc_hd__mux4_1 _12236_ (.A0(\core_pipeline.pipeline_registers.registers[12][15] ),
    .A1(\core_pipeline.pipeline_registers.registers[13][15] ),
    .A2(\core_pipeline.pipeline_registers.registers[14][15] ),
    .A3(\core_pipeline.pipeline_registers.registers[15][15] ),
    .S0(net613),
    .S1(net591),
    .X(_02555_));
 sky130_fd_sc_hd__or2_1 _12237_ (.A(net476),
    .B(_02555_),
    .X(_02556_));
 sky130_fd_sc_hd__o21a_1 _12238_ (.A1(net578),
    .A2(_02554_),
    .B1(net572),
    .X(_02557_));
 sky130_fd_sc_hd__a221o_1 _12239_ (.A1(net469),
    .A2(_02553_),
    .B1(_02556_),
    .B2(_02557_),
    .C1(net567),
    .X(_02558_));
 sky130_fd_sc_hd__mux2_1 _12240_ (.A0(\core_pipeline.pipeline_registers.registers[30][15] ),
    .A1(\core_pipeline.pipeline_registers.registers[31][15] ),
    .S(net609),
    .X(_02559_));
 sky130_fd_sc_hd__and2_1 _12241_ (.A(net588),
    .B(_02559_),
    .X(_02560_));
 sky130_fd_sc_hd__mux2_1 _12242_ (.A0(\core_pipeline.pipeline_registers.registers[28][15] ),
    .A1(\core_pipeline.pipeline_registers.registers[29][15] ),
    .S(net609),
    .X(_02561_));
 sky130_fd_sc_hd__a21o_1 _12243_ (.A1(net483),
    .A2(_02561_),
    .B1(net475),
    .X(_02562_));
 sky130_fd_sc_hd__mux2_1 _12244_ (.A0(\core_pipeline.pipeline_registers.registers[26][15] ),
    .A1(\core_pipeline.pipeline_registers.registers[27][15] ),
    .S(net609),
    .X(_02563_));
 sky130_fd_sc_hd__and2_1 _12245_ (.A(net588),
    .B(_02563_),
    .X(_02564_));
 sky130_fd_sc_hd__mux2_1 _12246_ (.A0(\core_pipeline.pipeline_registers.registers[24][15] ),
    .A1(\core_pipeline.pipeline_registers.registers[25][15] ),
    .S(net609),
    .X(_02565_));
 sky130_fd_sc_hd__a21o_1 _12247_ (.A1(net483),
    .A2(_02565_),
    .B1(net577),
    .X(_02566_));
 sky130_fd_sc_hd__o221a_1 _12248_ (.A1(_02560_),
    .A2(_02562_),
    .B1(_02564_),
    .B2(_02566_),
    .C1(net571),
    .X(_02567_));
 sky130_fd_sc_hd__mux2_1 _12249_ (.A0(_02551_),
    .A1(_02552_),
    .S(net476),
    .X(_02568_));
 sky130_fd_sc_hd__a211o_1 _12250_ (.A1(net469),
    .A2(_02568_),
    .B1(_02567_),
    .C1(net467),
    .X(_02569_));
 sky130_fd_sc_hd__and3_1 _12251_ (.A(net140),
    .B(_02558_),
    .C(_02569_),
    .X(_02570_));
 sky130_fd_sc_hd__a21o_1 _12252_ (.A1(\core_pipeline.decode_to_execute_rs1_data[15] ),
    .A2(net122),
    .B1(_02570_),
    .X(_01936_));
 sky130_fd_sc_hd__mux4_1 _12253_ (.A0(\core_pipeline.pipeline_registers.registers[4][16] ),
    .A1(\core_pipeline.pipeline_registers.registers[5][16] ),
    .A2(\core_pipeline.pipeline_registers.registers[6][16] ),
    .A3(\core_pipeline.pipeline_registers.registers[7][16] ),
    .S0(net603),
    .S1(net582),
    .X(_02571_));
 sky130_fd_sc_hd__mux4_1 _12254_ (.A0(\core_pipeline.pipeline_registers.registers[0][16] ),
    .A1(\core_pipeline.pipeline_registers.registers[1][16] ),
    .A2(\core_pipeline.pipeline_registers.registers[2][16] ),
    .A3(\core_pipeline.pipeline_registers.registers[3][16] ),
    .S0(net604),
    .S1(net583),
    .X(_02572_));
 sky130_fd_sc_hd__mux4_1 _12255_ (.A0(\core_pipeline.pipeline_registers.registers[20][16] ),
    .A1(\core_pipeline.pipeline_registers.registers[21][16] ),
    .A2(\core_pipeline.pipeline_registers.registers[22][16] ),
    .A3(\core_pipeline.pipeline_registers.registers[23][16] ),
    .S0(net607),
    .S1(net586),
    .X(_02573_));
 sky130_fd_sc_hd__mux4_1 _12256_ (.A0(\core_pipeline.pipeline_registers.registers[16][16] ),
    .A1(\core_pipeline.pipeline_registers.registers[17][16] ),
    .A2(\core_pipeline.pipeline_registers.registers[18][16] ),
    .A3(\core_pipeline.pipeline_registers.registers[19][16] ),
    .S0(net607),
    .S1(net586),
    .X(_02574_));
 sky130_fd_sc_hd__mux2_1 _12257_ (.A0(_02571_),
    .A1(_02572_),
    .S(net472),
    .X(_02575_));
 sky130_fd_sc_hd__mux4_1 _12258_ (.A0(\core_pipeline.pipeline_registers.registers[8][16] ),
    .A1(\core_pipeline.pipeline_registers.registers[9][16] ),
    .A2(\core_pipeline.pipeline_registers.registers[10][16] ),
    .A3(\core_pipeline.pipeline_registers.registers[11][16] ),
    .S0(net604),
    .S1(net583),
    .X(_02576_));
 sky130_fd_sc_hd__mux4_1 _12259_ (.A0(\core_pipeline.pipeline_registers.registers[12][16] ),
    .A1(\core_pipeline.pipeline_registers.registers[13][16] ),
    .A2(\core_pipeline.pipeline_registers.registers[14][16] ),
    .A3(\core_pipeline.pipeline_registers.registers[15][16] ),
    .S0(net604),
    .S1(net583),
    .X(_02577_));
 sky130_fd_sc_hd__or2_1 _12260_ (.A(net472),
    .B(_02577_),
    .X(_02578_));
 sky130_fd_sc_hd__o21a_1 _12261_ (.A1(net576),
    .A2(_02576_),
    .B1(net570),
    .X(_02579_));
 sky130_fd_sc_hd__a221o_1 _12262_ (.A1(net468),
    .A2(_02575_),
    .B1(_02578_),
    .B2(_02579_),
    .C1(net567),
    .X(_02580_));
 sky130_fd_sc_hd__mux2_1 _12263_ (.A0(\core_pipeline.pipeline_registers.registers[30][16] ),
    .A1(\core_pipeline.pipeline_registers.registers[31][16] ),
    .S(net607),
    .X(_02581_));
 sky130_fd_sc_hd__and2_1 _12264_ (.A(net586),
    .B(_02581_),
    .X(_02582_));
 sky130_fd_sc_hd__mux2_1 _12265_ (.A0(\core_pipeline.pipeline_registers.registers[28][16] ),
    .A1(\core_pipeline.pipeline_registers.registers[29][16] ),
    .S(net607),
    .X(_02583_));
 sky130_fd_sc_hd__a21o_1 _12266_ (.A1(net482),
    .A2(_02583_),
    .B1(net473),
    .X(_02584_));
 sky130_fd_sc_hd__mux2_1 _12267_ (.A0(\core_pipeline.pipeline_registers.registers[26][16] ),
    .A1(\core_pipeline.pipeline_registers.registers[27][16] ),
    .S(net607),
    .X(_02585_));
 sky130_fd_sc_hd__and2_1 _12268_ (.A(net586),
    .B(_02585_),
    .X(_02586_));
 sky130_fd_sc_hd__mux2_1 _12269_ (.A0(\core_pipeline.pipeline_registers.registers[24][16] ),
    .A1(\core_pipeline.pipeline_registers.registers[25][16] ),
    .S(net607),
    .X(_02587_));
 sky130_fd_sc_hd__a21o_1 _12270_ (.A1(net482),
    .A2(_02587_),
    .B1(net577),
    .X(_02588_));
 sky130_fd_sc_hd__o221a_1 _12271_ (.A1(_02582_),
    .A2(_02584_),
    .B1(_02586_),
    .B2(_02588_),
    .C1(net571),
    .X(_02589_));
 sky130_fd_sc_hd__mux2_1 _12272_ (.A0(_02573_),
    .A1(_02574_),
    .S(net473),
    .X(_02590_));
 sky130_fd_sc_hd__a211o_1 _12273_ (.A1(net468),
    .A2(_02590_),
    .B1(_02589_),
    .C1(net467),
    .X(_02591_));
 sky130_fd_sc_hd__and3_2 _12274_ (.A(net144),
    .B(_02580_),
    .C(_02591_),
    .X(_02592_));
 sky130_fd_sc_hd__a21o_1 _12275_ (.A1(\core_pipeline.decode_to_execute_rs1_data[16] ),
    .A2(net124),
    .B1(_02592_),
    .X(_01937_));
 sky130_fd_sc_hd__mux4_1 _12276_ (.A0(\core_pipeline.pipeline_registers.registers[4][17] ),
    .A1(\core_pipeline.pipeline_registers.registers[5][17] ),
    .A2(\core_pipeline.pipeline_registers.registers[6][17] ),
    .A3(\core_pipeline.pipeline_registers.registers[7][17] ),
    .S0(net621),
    .S1(net598),
    .X(_02593_));
 sky130_fd_sc_hd__mux4_1 _12277_ (.A0(\core_pipeline.pipeline_registers.registers[0][17] ),
    .A1(\core_pipeline.pipeline_registers.registers[1][17] ),
    .A2(\core_pipeline.pipeline_registers.registers[2][17] ),
    .A3(\core_pipeline.pipeline_registers.registers[3][17] ),
    .S0(net621),
    .S1(net598),
    .X(_02594_));
 sky130_fd_sc_hd__mux4_1 _12278_ (.A0(\core_pipeline.pipeline_registers.registers[20][17] ),
    .A1(\core_pipeline.pipeline_registers.registers[21][17] ),
    .A2(\core_pipeline.pipeline_registers.registers[22][17] ),
    .A3(\core_pipeline.pipeline_registers.registers[23][17] ),
    .S0(net621),
    .S1(net598),
    .X(_02595_));
 sky130_fd_sc_hd__mux4_1 _12279_ (.A0(\core_pipeline.pipeline_registers.registers[16][17] ),
    .A1(\core_pipeline.pipeline_registers.registers[17][17] ),
    .A2(\core_pipeline.pipeline_registers.registers[18][17] ),
    .A3(\core_pipeline.pipeline_registers.registers[19][17] ),
    .S0(net622),
    .S1(net598),
    .X(_02596_));
 sky130_fd_sc_hd__mux2_1 _12280_ (.A0(_02593_),
    .A1(_02594_),
    .S(net478),
    .X(_02597_));
 sky130_fd_sc_hd__mux4_1 _12281_ (.A0(\core_pipeline.pipeline_registers.registers[8][17] ),
    .A1(\core_pipeline.pipeline_registers.registers[9][17] ),
    .A2(\core_pipeline.pipeline_registers.registers[10][17] ),
    .A3(\core_pipeline.pipeline_registers.registers[11][17] ),
    .S0(net617),
    .S1(net594),
    .X(_02598_));
 sky130_fd_sc_hd__mux4_1 _12282_ (.A0(\core_pipeline.pipeline_registers.registers[12][17] ),
    .A1(\core_pipeline.pipeline_registers.registers[13][17] ),
    .A2(\core_pipeline.pipeline_registers.registers[14][17] ),
    .A3(\core_pipeline.pipeline_registers.registers[15][17] ),
    .S0(net618),
    .S1(net595),
    .X(_02599_));
 sky130_fd_sc_hd__or2_1 _12283_ (.A(net477),
    .B(_02599_),
    .X(_02600_));
 sky130_fd_sc_hd__o21a_1 _12284_ (.A1(net579),
    .A2(_02598_),
    .B1(net573),
    .X(_02601_));
 sky130_fd_sc_hd__a221o_1 _12285_ (.A1(net470),
    .A2(_02597_),
    .B1(_02600_),
    .B2(_02601_),
    .C1(net568),
    .X(_02602_));
 sky130_fd_sc_hd__mux2_1 _12286_ (.A0(\core_pipeline.pipeline_registers.registers[30][17] ),
    .A1(\core_pipeline.pipeline_registers.registers[31][17] ),
    .S(net621),
    .X(_02603_));
 sky130_fd_sc_hd__and2_1 _12287_ (.A(net598),
    .B(_02603_),
    .X(_02604_));
 sky130_fd_sc_hd__mux2_1 _12288_ (.A0(\core_pipeline.pipeline_registers.registers[28][17] ),
    .A1(\core_pipeline.pipeline_registers.registers[29][17] ),
    .S(net621),
    .X(_02605_));
 sky130_fd_sc_hd__a21o_1 _12289_ (.A1(net484),
    .A2(_02605_),
    .B1(net478),
    .X(_02606_));
 sky130_fd_sc_hd__mux2_1 _12290_ (.A0(\core_pipeline.pipeline_registers.registers[26][17] ),
    .A1(\core_pipeline.pipeline_registers.registers[27][17] ),
    .S(net619),
    .X(_02607_));
 sky130_fd_sc_hd__and2_1 _12291_ (.A(net596),
    .B(_02607_),
    .X(_02608_));
 sky130_fd_sc_hd__mux2_1 _12292_ (.A0(\core_pipeline.pipeline_registers.registers[24][17] ),
    .A1(\core_pipeline.pipeline_registers.registers[25][17] ),
    .S(net621),
    .X(_02609_));
 sky130_fd_sc_hd__a21o_1 _12293_ (.A1(net484),
    .A2(_02609_),
    .B1(net579),
    .X(_02610_));
 sky130_fd_sc_hd__o221a_1 _12294_ (.A1(_02604_),
    .A2(_02606_),
    .B1(_02608_),
    .B2(_02610_),
    .C1(net573),
    .X(_02611_));
 sky130_fd_sc_hd__mux2_1 _12295_ (.A0(_02595_),
    .A1(_02596_),
    .S(net479),
    .X(_02612_));
 sky130_fd_sc_hd__a211o_1 _12296_ (.A1(net470),
    .A2(_02612_),
    .B1(_02611_),
    .C1(net466),
    .X(_02613_));
 sky130_fd_sc_hd__and3_1 _12297_ (.A(net148),
    .B(_02602_),
    .C(_02613_),
    .X(_02614_));
 sky130_fd_sc_hd__a21o_1 _12298_ (.A1(\core_pipeline.decode_to_execute_rs1_data[17] ),
    .A2(net131),
    .B1(_02614_),
    .X(_01938_));
 sky130_fd_sc_hd__mux4_1 _12299_ (.A0(\core_pipeline.pipeline_registers.registers[4][18] ),
    .A1(\core_pipeline.pipeline_registers.registers[5][18] ),
    .A2(\core_pipeline.pipeline_registers.registers[6][18] ),
    .A3(\core_pipeline.pipeline_registers.registers[7][18] ),
    .S0(net622),
    .S1(net598),
    .X(_02615_));
 sky130_fd_sc_hd__mux4_1 _12300_ (.A0(\core_pipeline.pipeline_registers.registers[0][18] ),
    .A1(\core_pipeline.pipeline_registers.registers[1][18] ),
    .A2(\core_pipeline.pipeline_registers.registers[2][18] ),
    .A3(\core_pipeline.pipeline_registers.registers[3][18] ),
    .S0(net622),
    .S1(net598),
    .X(_02616_));
 sky130_fd_sc_hd__mux4_1 _12301_ (.A0(\core_pipeline.pipeline_registers.registers[20][18] ),
    .A1(\core_pipeline.pipeline_registers.registers[21][18] ),
    .A2(\core_pipeline.pipeline_registers.registers[22][18] ),
    .A3(\core_pipeline.pipeline_registers.registers[23][18] ),
    .S0(net622),
    .S1(net598),
    .X(_02617_));
 sky130_fd_sc_hd__mux4_1 _12302_ (.A0(\core_pipeline.pipeline_registers.registers[16][18] ),
    .A1(\core_pipeline.pipeline_registers.registers[17][18] ),
    .A2(\core_pipeline.pipeline_registers.registers[18][18] ),
    .A3(\core_pipeline.pipeline_registers.registers[19][18] ),
    .S0(net621),
    .S1(net598),
    .X(_02618_));
 sky130_fd_sc_hd__mux2_1 _12303_ (.A0(_02615_),
    .A1(_02616_),
    .S(net479),
    .X(_02619_));
 sky130_fd_sc_hd__mux4_1 _12304_ (.A0(\core_pipeline.pipeline_registers.registers[8][18] ),
    .A1(\core_pipeline.pipeline_registers.registers[9][18] ),
    .A2(\core_pipeline.pipeline_registers.registers[10][18] ),
    .A3(\core_pipeline.pipeline_registers.registers[11][18] ),
    .S0(net620),
    .S1(net596),
    .X(_02620_));
 sky130_fd_sc_hd__mux4_1 _12305_ (.A0(\core_pipeline.pipeline_registers.registers[12][18] ),
    .A1(\core_pipeline.pipeline_registers.registers[13][18] ),
    .A2(\core_pipeline.pipeline_registers.registers[14][18] ),
    .A3(\core_pipeline.pipeline_registers.registers[15][18] ),
    .S0(net620),
    .S1(net596),
    .X(_02621_));
 sky130_fd_sc_hd__or2_1 _12306_ (.A(net478),
    .B(_02621_),
    .X(_02622_));
 sky130_fd_sc_hd__o21a_1 _12307_ (.A1(net580),
    .A2(_02620_),
    .B1(net574),
    .X(_02623_));
 sky130_fd_sc_hd__a221o_2 _12308_ (.A1(net470),
    .A2(_02619_),
    .B1(_02622_),
    .B2(_02623_),
    .C1(net568),
    .X(_02624_));
 sky130_fd_sc_hd__mux2_1 _12309_ (.A0(\core_pipeline.pipeline_registers.registers[30][18] ),
    .A1(\core_pipeline.pipeline_registers.registers[31][18] ),
    .S(net621),
    .X(_02625_));
 sky130_fd_sc_hd__and2_1 _12310_ (.A(net598),
    .B(_02625_),
    .X(_02626_));
 sky130_fd_sc_hd__mux2_1 _12311_ (.A0(\core_pipeline.pipeline_registers.registers[28][18] ),
    .A1(\core_pipeline.pipeline_registers.registers[29][18] ),
    .S(net621),
    .X(_02627_));
 sky130_fd_sc_hd__a21o_1 _12312_ (.A1(net484),
    .A2(_02627_),
    .B1(net478),
    .X(_02628_));
 sky130_fd_sc_hd__mux2_1 _12313_ (.A0(\core_pipeline.pipeline_registers.registers[26][18] ),
    .A1(\core_pipeline.pipeline_registers.registers[27][18] ),
    .S(net621),
    .X(_02629_));
 sky130_fd_sc_hd__and2_1 _12314_ (.A(net598),
    .B(_02629_),
    .X(_02630_));
 sky130_fd_sc_hd__mux2_1 _12315_ (.A0(\core_pipeline.pipeline_registers.registers[24][18] ),
    .A1(\core_pipeline.pipeline_registers.registers[25][18] ),
    .S(net621),
    .X(_02631_));
 sky130_fd_sc_hd__a21o_1 _12316_ (.A1(net484),
    .A2(_02631_),
    .B1(net580),
    .X(_02632_));
 sky130_fd_sc_hd__o221a_1 _12317_ (.A1(_02626_),
    .A2(_02628_),
    .B1(_02630_),
    .B2(_02632_),
    .C1(net574),
    .X(_02633_));
 sky130_fd_sc_hd__mux2_1 _12318_ (.A0(_02617_),
    .A1(_02618_),
    .S(net478),
    .X(_02634_));
 sky130_fd_sc_hd__a211o_1 _12319_ (.A1(net470),
    .A2(_02634_),
    .B1(_02633_),
    .C1(net466),
    .X(_02635_));
 sky130_fd_sc_hd__and3_1 _12320_ (.A(net148),
    .B(_02624_),
    .C(_02635_),
    .X(_02636_));
 sky130_fd_sc_hd__a21o_1 _12321_ (.A1(\core_pipeline.decode_to_execute_rs1_data[18] ),
    .A2(net135),
    .B1(_02636_),
    .X(_01939_));
 sky130_fd_sc_hd__mux4_1 _12322_ (.A0(\core_pipeline.pipeline_registers.registers[4][19] ),
    .A1(\core_pipeline.pipeline_registers.registers[5][19] ),
    .A2(\core_pipeline.pipeline_registers.registers[6][19] ),
    .A3(\core_pipeline.pipeline_registers.registers[7][19] ),
    .S0(net619),
    .S1(net596),
    .X(_02637_));
 sky130_fd_sc_hd__mux4_1 _12323_ (.A0(\core_pipeline.pipeline_registers.registers[0][19] ),
    .A1(\core_pipeline.pipeline_registers.registers[1][19] ),
    .A2(\core_pipeline.pipeline_registers.registers[2][19] ),
    .A3(\core_pipeline.pipeline_registers.registers[3][19] ),
    .S0(net619),
    .S1(net596),
    .X(_02638_));
 sky130_fd_sc_hd__mux4_1 _12324_ (.A0(\core_pipeline.pipeline_registers.registers[20][19] ),
    .A1(\core_pipeline.pipeline_registers.registers[21][19] ),
    .A2(\core_pipeline.pipeline_registers.registers[22][19] ),
    .A3(\core_pipeline.pipeline_registers.registers[23][19] ),
    .S0(net619),
    .S1(net596),
    .X(_02639_));
 sky130_fd_sc_hd__mux4_1 _12325_ (.A0(\core_pipeline.pipeline_registers.registers[16][19] ),
    .A1(\core_pipeline.pipeline_registers.registers[17][19] ),
    .A2(\core_pipeline.pipeline_registers.registers[18][19] ),
    .A3(\core_pipeline.pipeline_registers.registers[19][19] ),
    .S0(net619),
    .S1(net596),
    .X(_02640_));
 sky130_fd_sc_hd__mux2_1 _12326_ (.A0(_02637_),
    .A1(_02638_),
    .S(net478),
    .X(_02641_));
 sky130_fd_sc_hd__mux4_1 _12327_ (.A0(\core_pipeline.pipeline_registers.registers[8][19] ),
    .A1(\core_pipeline.pipeline_registers.registers[9][19] ),
    .A2(\core_pipeline.pipeline_registers.registers[10][19] ),
    .A3(\core_pipeline.pipeline_registers.registers[11][19] ),
    .S0(net619),
    .S1(net596),
    .X(_02642_));
 sky130_fd_sc_hd__mux4_1 _12328_ (.A0(\core_pipeline.pipeline_registers.registers[12][19] ),
    .A1(\core_pipeline.pipeline_registers.registers[13][19] ),
    .A2(\core_pipeline.pipeline_registers.registers[14][19] ),
    .A3(\core_pipeline.pipeline_registers.registers[15][19] ),
    .S0(net619),
    .S1(net596),
    .X(_02643_));
 sky130_fd_sc_hd__or2_1 _12329_ (.A(net478),
    .B(_02643_),
    .X(_02644_));
 sky130_fd_sc_hd__o21a_1 _12330_ (.A1(net580),
    .A2(_02642_),
    .B1(net574),
    .X(_02645_));
 sky130_fd_sc_hd__a221o_1 _12331_ (.A1(net471),
    .A2(_02641_),
    .B1(_02644_),
    .B2(_02645_),
    .C1(net568),
    .X(_02646_));
 sky130_fd_sc_hd__mux2_1 _12332_ (.A0(\core_pipeline.pipeline_registers.registers[30][19] ),
    .A1(\core_pipeline.pipeline_registers.registers[31][19] ),
    .S(net620),
    .X(_02647_));
 sky130_fd_sc_hd__and2_1 _12333_ (.A(net596),
    .B(_02647_),
    .X(_02648_));
 sky130_fd_sc_hd__mux2_1 _12334_ (.A0(\core_pipeline.pipeline_registers.registers[28][19] ),
    .A1(\core_pipeline.pipeline_registers.registers[29][19] ),
    .S(net619),
    .X(_02649_));
 sky130_fd_sc_hd__a21o_1 _12335_ (.A1(net485),
    .A2(_02649_),
    .B1(net478),
    .X(_02650_));
 sky130_fd_sc_hd__mux2_1 _12336_ (.A0(\core_pipeline.pipeline_registers.registers[26][19] ),
    .A1(\core_pipeline.pipeline_registers.registers[27][19] ),
    .S(net619),
    .X(_02651_));
 sky130_fd_sc_hd__and2_1 _12337_ (.A(net596),
    .B(_02651_),
    .X(_02652_));
 sky130_fd_sc_hd__mux2_1 _12338_ (.A0(\core_pipeline.pipeline_registers.registers[24][19] ),
    .A1(\core_pipeline.pipeline_registers.registers[25][19] ),
    .S(net619),
    .X(_02653_));
 sky130_fd_sc_hd__a21o_1 _12339_ (.A1(net485),
    .A2(_02653_),
    .B1(net580),
    .X(_02654_));
 sky130_fd_sc_hd__o221a_1 _12340_ (.A1(_02648_),
    .A2(_02650_),
    .B1(_02652_),
    .B2(_02654_),
    .C1(net574),
    .X(_02655_));
 sky130_fd_sc_hd__mux2_1 _12341_ (.A0(_02639_),
    .A1(_02640_),
    .S(net478),
    .X(_02656_));
 sky130_fd_sc_hd__a211o_1 _12342_ (.A1(net471),
    .A2(_02656_),
    .B1(_02655_),
    .C1(net466),
    .X(_02657_));
 sky130_fd_sc_hd__and3_2 _12343_ (.A(net145),
    .B(_02646_),
    .C(_02657_),
    .X(_02658_));
 sky130_fd_sc_hd__a21o_1 _12344_ (.A1(\core_pipeline.decode_to_execute_rs1_data[19] ),
    .A2(net135),
    .B1(_02658_),
    .X(_01940_));
 sky130_fd_sc_hd__mux4_1 _12345_ (.A0(\core_pipeline.pipeline_registers.registers[4][20] ),
    .A1(\core_pipeline.pipeline_registers.registers[5][20] ),
    .A2(\core_pipeline.pipeline_registers.registers[6][20] ),
    .A3(\core_pipeline.pipeline_registers.registers[7][20] ),
    .S0(net620),
    .S1(net597),
    .X(_02659_));
 sky130_fd_sc_hd__mux4_1 _12346_ (.A0(\core_pipeline.pipeline_registers.registers[0][20] ),
    .A1(\core_pipeline.pipeline_registers.registers[1][20] ),
    .A2(\core_pipeline.pipeline_registers.registers[2][20] ),
    .A3(\core_pipeline.pipeline_registers.registers[3][20] ),
    .S0(net620),
    .S1(net597),
    .X(_02660_));
 sky130_fd_sc_hd__mux4_1 _12347_ (.A0(\core_pipeline.pipeline_registers.registers[20][20] ),
    .A1(\core_pipeline.pipeline_registers.registers[21][20] ),
    .A2(\core_pipeline.pipeline_registers.registers[22][20] ),
    .A3(\core_pipeline.pipeline_registers.registers[23][20] ),
    .S0(net620),
    .S1(net597),
    .X(_02661_));
 sky130_fd_sc_hd__mux4_1 _12348_ (.A0(\core_pipeline.pipeline_registers.registers[16][20] ),
    .A1(\core_pipeline.pipeline_registers.registers[17][20] ),
    .A2(\core_pipeline.pipeline_registers.registers[18][20] ),
    .A3(\core_pipeline.pipeline_registers.registers[19][20] ),
    .S0(net620),
    .S1(net597),
    .X(_02662_));
 sky130_fd_sc_hd__mux2_1 _12349_ (.A0(_02659_),
    .A1(_02660_),
    .S(net478),
    .X(_02663_));
 sky130_fd_sc_hd__mux4_1 _12350_ (.A0(\core_pipeline.pipeline_registers.registers[8][20] ),
    .A1(\core_pipeline.pipeline_registers.registers[9][20] ),
    .A2(\core_pipeline.pipeline_registers.registers[10][20] ),
    .A3(\core_pipeline.pipeline_registers.registers[11][20] ),
    .S0(net620),
    .S1(net597),
    .X(_02664_));
 sky130_fd_sc_hd__mux4_1 _12351_ (.A0(\core_pipeline.pipeline_registers.registers[12][20] ),
    .A1(\core_pipeline.pipeline_registers.registers[13][20] ),
    .A2(\core_pipeline.pipeline_registers.registers[14][20] ),
    .A3(\core_pipeline.pipeline_registers.registers[15][20] ),
    .S0(net620),
    .S1(net597),
    .X(_02665_));
 sky130_fd_sc_hd__or2_1 _12352_ (.A(net478),
    .B(_02665_),
    .X(_02666_));
 sky130_fd_sc_hd__o21a_1 _12353_ (.A1(net580),
    .A2(_02664_),
    .B1(net574),
    .X(_02667_));
 sky130_fd_sc_hd__a221o_1 _12354_ (.A1(net470),
    .A2(_02663_),
    .B1(_02666_),
    .B2(_02667_),
    .C1(net568),
    .X(_02668_));
 sky130_fd_sc_hd__mux2_1 _12355_ (.A0(\core_pipeline.pipeline_registers.registers[30][20] ),
    .A1(\core_pipeline.pipeline_registers.registers[31][20] ),
    .S(net620),
    .X(_02669_));
 sky130_fd_sc_hd__and2_1 _12356_ (.A(net597),
    .B(_02669_),
    .X(_02670_));
 sky130_fd_sc_hd__mux2_1 _12357_ (.A0(\core_pipeline.pipeline_registers.registers[28][20] ),
    .A1(\core_pipeline.pipeline_registers.registers[29][20] ),
    .S(net620),
    .X(_02671_));
 sky130_fd_sc_hd__a21o_1 _12358_ (.A1(net484),
    .A2(_02671_),
    .B1(net478),
    .X(_02672_));
 sky130_fd_sc_hd__mux2_1 _12359_ (.A0(\core_pipeline.pipeline_registers.registers[26][20] ),
    .A1(\core_pipeline.pipeline_registers.registers[27][20] ),
    .S(net620),
    .X(_02673_));
 sky130_fd_sc_hd__and2_1 _12360_ (.A(net597),
    .B(_02673_),
    .X(_02674_));
 sky130_fd_sc_hd__mux2_1 _12361_ (.A0(\core_pipeline.pipeline_registers.registers[24][20] ),
    .A1(\core_pipeline.pipeline_registers.registers[25][20] ),
    .S(net620),
    .X(_02675_));
 sky130_fd_sc_hd__a21o_1 _12362_ (.A1(net484),
    .A2(_02675_),
    .B1(net580),
    .X(_02676_));
 sky130_fd_sc_hd__o221a_1 _12363_ (.A1(_02670_),
    .A2(_02672_),
    .B1(_02674_),
    .B2(_02676_),
    .C1(net574),
    .X(_02677_));
 sky130_fd_sc_hd__mux2_1 _12364_ (.A0(_02661_),
    .A1(_02662_),
    .S(net478),
    .X(_02678_));
 sky130_fd_sc_hd__a211o_1 _12365_ (.A1(net470),
    .A2(_02678_),
    .B1(_02677_),
    .C1(net466),
    .X(_02679_));
 sky130_fd_sc_hd__and3_1 _12366_ (.A(net145),
    .B(_02668_),
    .C(_02679_),
    .X(_02680_));
 sky130_fd_sc_hd__a21o_1 _12367_ (.A1(\core_pipeline.decode_to_execute_rs1_data[20] ),
    .A2(net135),
    .B1(_02680_),
    .X(_01941_));
 sky130_fd_sc_hd__mux4_1 _12368_ (.A0(\core_pipeline.pipeline_registers.registers[4][21] ),
    .A1(\core_pipeline.pipeline_registers.registers[5][21] ),
    .A2(\core_pipeline.pipeline_registers.registers[6][21] ),
    .A3(\core_pipeline.pipeline_registers.registers[7][21] ),
    .S0(net624),
    .S1(net601),
    .X(_02681_));
 sky130_fd_sc_hd__mux4_1 _12369_ (.A0(\core_pipeline.pipeline_registers.registers[0][21] ),
    .A1(\core_pipeline.pipeline_registers.registers[1][21] ),
    .A2(\core_pipeline.pipeline_registers.registers[2][21] ),
    .A3(\core_pipeline.pipeline_registers.registers[3][21] ),
    .S0(net624),
    .S1(net601),
    .X(_02682_));
 sky130_fd_sc_hd__mux4_1 _12370_ (.A0(\core_pipeline.pipeline_registers.registers[20][21] ),
    .A1(\core_pipeline.pipeline_registers.registers[21][21] ),
    .A2(\core_pipeline.pipeline_registers.registers[22][21] ),
    .A3(\core_pipeline.pipeline_registers.registers[23][21] ),
    .S0(net625),
    .S1(net601),
    .X(_02683_));
 sky130_fd_sc_hd__mux4_1 _12371_ (.A0(\core_pipeline.pipeline_registers.registers[16][21] ),
    .A1(\core_pipeline.pipeline_registers.registers[17][21] ),
    .A2(\core_pipeline.pipeline_registers.registers[18][21] ),
    .A3(\core_pipeline.pipeline_registers.registers[19][21] ),
    .S0(net624),
    .S1(net601),
    .X(_02684_));
 sky130_fd_sc_hd__mux2_1 _12372_ (.A0(_02681_),
    .A1(_02682_),
    .S(net479),
    .X(_02685_));
 sky130_fd_sc_hd__mux4_1 _12373_ (.A0(\core_pipeline.pipeline_registers.registers[8][21] ),
    .A1(\core_pipeline.pipeline_registers.registers[9][21] ),
    .A2(\core_pipeline.pipeline_registers.registers[10][21] ),
    .A3(\core_pipeline.pipeline_registers.registers[11][21] ),
    .S0(net625),
    .S1(net601),
    .X(_02686_));
 sky130_fd_sc_hd__mux4_1 _12374_ (.A0(\core_pipeline.pipeline_registers.registers[12][21] ),
    .A1(\core_pipeline.pipeline_registers.registers[13][21] ),
    .A2(\core_pipeline.pipeline_registers.registers[14][21] ),
    .A3(\core_pipeline.pipeline_registers.registers[15][21] ),
    .S0(net624),
    .S1(net602),
    .X(_02687_));
 sky130_fd_sc_hd__or2_1 _12375_ (.A(net479),
    .B(_02687_),
    .X(_02688_));
 sky130_fd_sc_hd__o21a_1 _12376_ (.A1(net581),
    .A2(_02686_),
    .B1(net575),
    .X(_02689_));
 sky130_fd_sc_hd__a221o_1 _12377_ (.A1(net471),
    .A2(_02685_),
    .B1(_02688_),
    .B2(_02689_),
    .C1(net569),
    .X(_02690_));
 sky130_fd_sc_hd__mux2_1 _12378_ (.A0(\core_pipeline.pipeline_registers.registers[30][21] ),
    .A1(\core_pipeline.pipeline_registers.registers[31][21] ),
    .S(net625),
    .X(_02691_));
 sky130_fd_sc_hd__and2_1 _12379_ (.A(net602),
    .B(_02691_),
    .X(_02692_));
 sky130_fd_sc_hd__mux2_1 _12380_ (.A0(\core_pipeline.pipeline_registers.registers[28][21] ),
    .A1(\core_pipeline.pipeline_registers.registers[29][21] ),
    .S(net625),
    .X(_02693_));
 sky130_fd_sc_hd__a21o_1 _12381_ (.A1(net485),
    .A2(_02693_),
    .B1(net479),
    .X(_02694_));
 sky130_fd_sc_hd__mux2_1 _12382_ (.A0(\core_pipeline.pipeline_registers.registers[26][21] ),
    .A1(\core_pipeline.pipeline_registers.registers[27][21] ),
    .S(net625),
    .X(_02695_));
 sky130_fd_sc_hd__and2_1 _12383_ (.A(net598),
    .B(_02695_),
    .X(_02696_));
 sky130_fd_sc_hd__mux2_1 _12384_ (.A0(\core_pipeline.pipeline_registers.registers[24][21] ),
    .A1(\core_pipeline.pipeline_registers.registers[25][21] ),
    .S(net621),
    .X(_02697_));
 sky130_fd_sc_hd__a21o_1 _12385_ (.A1(net485),
    .A2(_02697_),
    .B1(net580),
    .X(_02698_));
 sky130_fd_sc_hd__o221a_1 _12386_ (.A1(_02692_),
    .A2(_02694_),
    .B1(_02696_),
    .B2(_02698_),
    .C1(net575),
    .X(_02699_));
 sky130_fd_sc_hd__mux2_1 _12387_ (.A0(_02683_),
    .A1(_02684_),
    .S(net479),
    .X(_02700_));
 sky130_fd_sc_hd__a211o_1 _12388_ (.A1(net471),
    .A2(_02700_),
    .B1(_02699_),
    .C1(net466),
    .X(_02701_));
 sky130_fd_sc_hd__and3_1 _12389_ (.A(net146),
    .B(_02690_),
    .C(_02701_),
    .X(_02702_));
 sky130_fd_sc_hd__a21o_1 _12390_ (.A1(\core_pipeline.decode_to_execute_rs1_data[21] ),
    .A2(net134),
    .B1(_02702_),
    .X(_01942_));
 sky130_fd_sc_hd__mux4_1 _12391_ (.A0(\core_pipeline.pipeline_registers.registers[4][22] ),
    .A1(\core_pipeline.pipeline_registers.registers[5][22] ),
    .A2(\core_pipeline.pipeline_registers.registers[6][22] ),
    .A3(\core_pipeline.pipeline_registers.registers[7][22] ),
    .S0(net615),
    .S1(net592),
    .X(_02703_));
 sky130_fd_sc_hd__mux4_1 _12392_ (.A0(\core_pipeline.pipeline_registers.registers[0][22] ),
    .A1(\core_pipeline.pipeline_registers.registers[1][22] ),
    .A2(\core_pipeline.pipeline_registers.registers[2][22] ),
    .A3(\core_pipeline.pipeline_registers.registers[3][22] ),
    .S0(net615),
    .S1(net592),
    .X(_02704_));
 sky130_fd_sc_hd__mux4_1 _12393_ (.A0(\core_pipeline.pipeline_registers.registers[20][22] ),
    .A1(\core_pipeline.pipeline_registers.registers[21][22] ),
    .A2(\core_pipeline.pipeline_registers.registers[22][22] ),
    .A3(\core_pipeline.pipeline_registers.registers[23][22] ),
    .S0(net615),
    .S1(net592),
    .X(_02705_));
 sky130_fd_sc_hd__mux4_1 _12394_ (.A0(\core_pipeline.pipeline_registers.registers[16][22] ),
    .A1(\core_pipeline.pipeline_registers.registers[17][22] ),
    .A2(\core_pipeline.pipeline_registers.registers[18][22] ),
    .A3(\core_pipeline.pipeline_registers.registers[19][22] ),
    .S0(net615),
    .S1(net592),
    .X(_02706_));
 sky130_fd_sc_hd__mux2_1 _12395_ (.A0(_02703_),
    .A1(_02704_),
    .S(net477),
    .X(_02707_));
 sky130_fd_sc_hd__mux4_1 _12396_ (.A0(\core_pipeline.pipeline_registers.registers[8][22] ),
    .A1(\core_pipeline.pipeline_registers.registers[9][22] ),
    .A2(\core_pipeline.pipeline_registers.registers[10][22] ),
    .A3(\core_pipeline.pipeline_registers.registers[11][22] ),
    .S0(net615),
    .S1(net592),
    .X(_02708_));
 sky130_fd_sc_hd__mux4_1 _12397_ (.A0(\core_pipeline.pipeline_registers.registers[12][22] ),
    .A1(\core_pipeline.pipeline_registers.registers[13][22] ),
    .A2(\core_pipeline.pipeline_registers.registers[14][22] ),
    .A3(\core_pipeline.pipeline_registers.registers[15][22] ),
    .S0(net615),
    .S1(net592),
    .X(_02709_));
 sky130_fd_sc_hd__or2_1 _12398_ (.A(net477),
    .B(_02709_),
    .X(_02710_));
 sky130_fd_sc_hd__o21a_1 _12399_ (.A1(net579),
    .A2(_02708_),
    .B1(net573),
    .X(_02711_));
 sky130_fd_sc_hd__a221o_1 _12400_ (.A1(net470),
    .A2(_02707_),
    .B1(_02710_),
    .B2(_02711_),
    .C1(net568),
    .X(_02712_));
 sky130_fd_sc_hd__mux2_1 _12401_ (.A0(\core_pipeline.pipeline_registers.registers[30][22] ),
    .A1(\core_pipeline.pipeline_registers.registers[31][22] ),
    .S(net616),
    .X(_02713_));
 sky130_fd_sc_hd__and2_1 _12402_ (.A(net593),
    .B(_02713_),
    .X(_02714_));
 sky130_fd_sc_hd__mux2_1 _12403_ (.A0(\core_pipeline.pipeline_registers.registers[28][22] ),
    .A1(\core_pipeline.pipeline_registers.registers[29][22] ),
    .S(net616),
    .X(_02715_));
 sky130_fd_sc_hd__a21o_1 _12404_ (.A1(net484),
    .A2(_02715_),
    .B1(net481),
    .X(_02716_));
 sky130_fd_sc_hd__mux2_1 _12405_ (.A0(\core_pipeline.pipeline_registers.registers[26][22] ),
    .A1(\core_pipeline.pipeline_registers.registers[27][22] ),
    .S(net616),
    .X(_02717_));
 sky130_fd_sc_hd__and2_1 _12406_ (.A(net593),
    .B(_02717_),
    .X(_02718_));
 sky130_fd_sc_hd__mux2_1 _12407_ (.A0(\core_pipeline.pipeline_registers.registers[24][22] ),
    .A1(\core_pipeline.pipeline_registers.registers[25][22] ),
    .S(net616),
    .X(_02719_));
 sky130_fd_sc_hd__a21o_1 _12408_ (.A1(net484),
    .A2(_02719_),
    .B1(net579),
    .X(_02720_));
 sky130_fd_sc_hd__o221a_1 _12409_ (.A1(_02714_),
    .A2(_02716_),
    .B1(_02718_),
    .B2(_02720_),
    .C1(net573),
    .X(_02721_));
 sky130_fd_sc_hd__mux2_1 _12410_ (.A0(_02705_),
    .A1(_02706_),
    .S(net477),
    .X(_02722_));
 sky130_fd_sc_hd__a211o_1 _12411_ (.A1(net470),
    .A2(_02722_),
    .B1(_02721_),
    .C1(net466),
    .X(_02723_));
 sky130_fd_sc_hd__and3_1 _12412_ (.A(net145),
    .B(_02712_),
    .C(_02723_),
    .X(_02724_));
 sky130_fd_sc_hd__a21o_1 _12413_ (.A1(\core_pipeline.decode_to_execute_rs1_data[22] ),
    .A2(net131),
    .B1(_02724_),
    .X(_01943_));
 sky130_fd_sc_hd__mux4_1 _12414_ (.A0(\core_pipeline.pipeline_registers.registers[4][23] ),
    .A1(\core_pipeline.pipeline_registers.registers[5][23] ),
    .A2(\core_pipeline.pipeline_registers.registers[6][23] ),
    .A3(\core_pipeline.pipeline_registers.registers[7][23] ),
    .S0(net617),
    .S1(net594),
    .X(_02725_));
 sky130_fd_sc_hd__mux4_1 _12415_ (.A0(\core_pipeline.pipeline_registers.registers[0][23] ),
    .A1(\core_pipeline.pipeline_registers.registers[1][23] ),
    .A2(\core_pipeline.pipeline_registers.registers[2][23] ),
    .A3(\core_pipeline.pipeline_registers.registers[3][23] ),
    .S0(net617),
    .S1(net594),
    .X(_02726_));
 sky130_fd_sc_hd__mux4_1 _12416_ (.A0(\core_pipeline.pipeline_registers.registers[20][23] ),
    .A1(\core_pipeline.pipeline_registers.registers[21][23] ),
    .A2(\core_pipeline.pipeline_registers.registers[22][23] ),
    .A3(\core_pipeline.pipeline_registers.registers[23][23] ),
    .S0(net617),
    .S1(net594),
    .X(_02727_));
 sky130_fd_sc_hd__mux4_1 _12417_ (.A0(\core_pipeline.pipeline_registers.registers[16][23] ),
    .A1(\core_pipeline.pipeline_registers.registers[17][23] ),
    .A2(\core_pipeline.pipeline_registers.registers[18][23] ),
    .A3(\core_pipeline.pipeline_registers.registers[19][23] ),
    .S0(net617),
    .S1(net594),
    .X(_02728_));
 sky130_fd_sc_hd__mux2_1 _12418_ (.A0(_02725_),
    .A1(_02726_),
    .S(net480),
    .X(_02729_));
 sky130_fd_sc_hd__mux4_1 _12419_ (.A0(\core_pipeline.pipeline_registers.registers[8][23] ),
    .A1(\core_pipeline.pipeline_registers.registers[9][23] ),
    .A2(\core_pipeline.pipeline_registers.registers[10][23] ),
    .A3(\core_pipeline.pipeline_registers.registers[11][23] ),
    .S0(net617),
    .S1(net594),
    .X(_02730_));
 sky130_fd_sc_hd__mux4_1 _12420_ (.A0(\core_pipeline.pipeline_registers.registers[12][23] ),
    .A1(\core_pipeline.pipeline_registers.registers[13][23] ),
    .A2(\core_pipeline.pipeline_registers.registers[14][23] ),
    .A3(\core_pipeline.pipeline_registers.registers[15][23] ),
    .S0(net617),
    .S1(net594),
    .X(_02731_));
 sky130_fd_sc_hd__or2_1 _12421_ (.A(net480),
    .B(_02731_),
    .X(_02732_));
 sky130_fd_sc_hd__o21a_1 _12422_ (.A1(net579),
    .A2(_02730_),
    .B1(net573),
    .X(_02733_));
 sky130_fd_sc_hd__a221o_1 _12423_ (.A1(_03325_),
    .A2(_02729_),
    .B1(_02732_),
    .B2(_02733_),
    .C1(net568),
    .X(_02734_));
 sky130_fd_sc_hd__mux2_1 _12424_ (.A0(\core_pipeline.pipeline_registers.registers[30][23] ),
    .A1(\core_pipeline.pipeline_registers.registers[31][23] ),
    .S(net617),
    .X(_02735_));
 sky130_fd_sc_hd__and2_1 _12425_ (.A(net594),
    .B(_02735_),
    .X(_02736_));
 sky130_fd_sc_hd__mux2_1 _12426_ (.A0(\core_pipeline.pipeline_registers.registers[28][23] ),
    .A1(\core_pipeline.pipeline_registers.registers[29][23] ),
    .S(net617),
    .X(_02737_));
 sky130_fd_sc_hd__a21o_1 _12427_ (.A1(net485),
    .A2(_02737_),
    .B1(net480),
    .X(_02738_));
 sky130_fd_sc_hd__mux2_1 _12428_ (.A0(\core_pipeline.pipeline_registers.registers[26][23] ),
    .A1(\core_pipeline.pipeline_registers.registers[27][23] ),
    .S(net617),
    .X(_02739_));
 sky130_fd_sc_hd__and2_1 _12429_ (.A(net594),
    .B(_02739_),
    .X(_02740_));
 sky130_fd_sc_hd__mux2_1 _12430_ (.A0(\core_pipeline.pipeline_registers.registers[24][23] ),
    .A1(\core_pipeline.pipeline_registers.registers[25][23] ),
    .S(net617),
    .X(_02741_));
 sky130_fd_sc_hd__a21o_1 _12431_ (.A1(net485),
    .A2(_02741_),
    .B1(net579),
    .X(_02742_));
 sky130_fd_sc_hd__o221a_1 _12432_ (.A1(_02736_),
    .A2(_02738_),
    .B1(_02740_),
    .B2(_02742_),
    .C1(net573),
    .X(_02743_));
 sky130_fd_sc_hd__mux2_1 _12433_ (.A0(_02727_),
    .A1(_02728_),
    .S(net477),
    .X(_02744_));
 sky130_fd_sc_hd__a211o_1 _12434_ (.A1(net471),
    .A2(_02744_),
    .B1(_02743_),
    .C1(net466),
    .X(_02745_));
 sky130_fd_sc_hd__and3_1 _12435_ (.A(net145),
    .B(_02734_),
    .C(_02745_),
    .X(_02746_));
 sky130_fd_sc_hd__a21o_1 _12436_ (.A1(\core_pipeline.decode_to_execute_rs1_data[23] ),
    .A2(net130),
    .B1(_02746_),
    .X(_01944_));
 sky130_fd_sc_hd__mux4_1 _12437_ (.A0(\core_pipeline.pipeline_registers.registers[4][24] ),
    .A1(\core_pipeline.pipeline_registers.registers[5][24] ),
    .A2(\core_pipeline.pipeline_registers.registers[6][24] ),
    .A3(\core_pipeline.pipeline_registers.registers[7][24] ),
    .S0(net610),
    .S1(net588),
    .X(_02747_));
 sky130_fd_sc_hd__mux4_1 _12438_ (.A0(\core_pipeline.pipeline_registers.registers[0][24] ),
    .A1(\core_pipeline.pipeline_registers.registers[1][24] ),
    .A2(\core_pipeline.pipeline_registers.registers[2][24] ),
    .A3(\core_pipeline.pipeline_registers.registers[3][24] ),
    .S0(net610),
    .S1(net588),
    .X(_02748_));
 sky130_fd_sc_hd__mux4_1 _12439_ (.A0(\core_pipeline.pipeline_registers.registers[20][24] ),
    .A1(\core_pipeline.pipeline_registers.registers[21][24] ),
    .A2(\core_pipeline.pipeline_registers.registers[22][24] ),
    .A3(\core_pipeline.pipeline_registers.registers[23][24] ),
    .S0(net610),
    .S1(net588),
    .X(_02749_));
 sky130_fd_sc_hd__mux4_1 _12440_ (.A0(\core_pipeline.pipeline_registers.registers[16][24] ),
    .A1(\core_pipeline.pipeline_registers.registers[17][24] ),
    .A2(\core_pipeline.pipeline_registers.registers[18][24] ),
    .A3(\core_pipeline.pipeline_registers.registers[19][24] ),
    .S0(net610),
    .S1(net588),
    .X(_02750_));
 sky130_fd_sc_hd__mux2_1 _12441_ (.A0(_02747_),
    .A1(_02748_),
    .S(net476),
    .X(_02751_));
 sky130_fd_sc_hd__mux4_1 _12442_ (.A0(\core_pipeline.pipeline_registers.registers[8][24] ),
    .A1(\core_pipeline.pipeline_registers.registers[9][24] ),
    .A2(\core_pipeline.pipeline_registers.registers[10][24] ),
    .A3(\core_pipeline.pipeline_registers.registers[11][24] ),
    .S0(net610),
    .S1(net589),
    .X(_02752_));
 sky130_fd_sc_hd__mux4_1 _12443_ (.A0(\core_pipeline.pipeline_registers.registers[12][24] ),
    .A1(\core_pipeline.pipeline_registers.registers[13][24] ),
    .A2(\core_pipeline.pipeline_registers.registers[14][24] ),
    .A3(\core_pipeline.pipeline_registers.registers[15][24] ),
    .S0(net610),
    .S1(net588),
    .X(_02753_));
 sky130_fd_sc_hd__or2_1 _12444_ (.A(net473),
    .B(_02753_),
    .X(_02754_));
 sky130_fd_sc_hd__o21a_1 _12445_ (.A1(net577),
    .A2(_02752_),
    .B1(net571),
    .X(_02755_));
 sky130_fd_sc_hd__a221o_1 _12446_ (.A1(net469),
    .A2(_02751_),
    .B1(_02754_),
    .B2(_02755_),
    .C1(net567),
    .X(_02756_));
 sky130_fd_sc_hd__mux2_1 _12447_ (.A0(\core_pipeline.pipeline_registers.registers[30][24] ),
    .A1(\core_pipeline.pipeline_registers.registers[31][24] ),
    .S(net610),
    .X(_02757_));
 sky130_fd_sc_hd__and2_1 _12448_ (.A(net588),
    .B(_02757_),
    .X(_02758_));
 sky130_fd_sc_hd__mux2_1 _12449_ (.A0(\core_pipeline.pipeline_registers.registers[28][24] ),
    .A1(\core_pipeline.pipeline_registers.registers[29][24] ),
    .S(net610),
    .X(_02759_));
 sky130_fd_sc_hd__a21o_1 _12450_ (.A1(net483),
    .A2(_02759_),
    .B1(net476),
    .X(_02760_));
 sky130_fd_sc_hd__mux2_1 _12451_ (.A0(\core_pipeline.pipeline_registers.registers[26][24] ),
    .A1(\core_pipeline.pipeline_registers.registers[27][24] ),
    .S(net610),
    .X(_02761_));
 sky130_fd_sc_hd__and2_1 _12452_ (.A(net588),
    .B(_02761_),
    .X(_02762_));
 sky130_fd_sc_hd__mux2_1 _12453_ (.A0(\core_pipeline.pipeline_registers.registers[24][24] ),
    .A1(\core_pipeline.pipeline_registers.registers[25][24] ),
    .S(net610),
    .X(_02763_));
 sky130_fd_sc_hd__a21o_1 _12454_ (.A1(net483),
    .A2(_02763_),
    .B1(net577),
    .X(_02764_));
 sky130_fd_sc_hd__o221a_1 _12455_ (.A1(_02758_),
    .A2(_02760_),
    .B1(_02762_),
    .B2(_02764_),
    .C1(net571),
    .X(_02765_));
 sky130_fd_sc_hd__mux2_1 _12456_ (.A0(_02749_),
    .A1(_02750_),
    .S(net476),
    .X(_02766_));
 sky130_fd_sc_hd__a211o_1 _12457_ (.A1(net469),
    .A2(_02766_),
    .B1(_02765_),
    .C1(net467),
    .X(_02767_));
 sky130_fd_sc_hd__and3_1 _12458_ (.A(net144),
    .B(_02756_),
    .C(_02767_),
    .X(_02768_));
 sky130_fd_sc_hd__a21o_1 _12459_ (.A1(\core_pipeline.decode_to_execute_rs1_data[24] ),
    .A2(net124),
    .B1(_02768_),
    .X(_01945_));
 sky130_fd_sc_hd__mux4_1 _12460_ (.A0(\core_pipeline.pipeline_registers.registers[4][25] ),
    .A1(\core_pipeline.pipeline_registers.registers[5][25] ),
    .A2(\core_pipeline.pipeline_registers.registers[6][25] ),
    .A3(\core_pipeline.pipeline_registers.registers[7][25] ),
    .S0(net612),
    .S1(net584),
    .X(_02769_));
 sky130_fd_sc_hd__mux4_1 _12461_ (.A0(\core_pipeline.pipeline_registers.registers[0][25] ),
    .A1(\core_pipeline.pipeline_registers.registers[1][25] ),
    .A2(\core_pipeline.pipeline_registers.registers[2][25] ),
    .A3(\core_pipeline.pipeline_registers.registers[3][25] ),
    .S0(net612),
    .S1(net590),
    .X(_02770_));
 sky130_fd_sc_hd__mux4_1 _12462_ (.A0(\core_pipeline.pipeline_registers.registers[20][25] ),
    .A1(\core_pipeline.pipeline_registers.registers[21][25] ),
    .A2(\core_pipeline.pipeline_registers.registers[22][25] ),
    .A3(\core_pipeline.pipeline_registers.registers[23][25] ),
    .S0(net606),
    .S1(net584),
    .X(_02771_));
 sky130_fd_sc_hd__mux4_1 _12463_ (.A0(\core_pipeline.pipeline_registers.registers[16][25] ),
    .A1(\core_pipeline.pipeline_registers.registers[17][25] ),
    .A2(\core_pipeline.pipeline_registers.registers[18][25] ),
    .A3(\core_pipeline.pipeline_registers.registers[19][25] ),
    .S0(net606),
    .S1(net584),
    .X(_02772_));
 sky130_fd_sc_hd__mux2_1 _12464_ (.A0(_02769_),
    .A1(_02770_),
    .S(net475),
    .X(_02773_));
 sky130_fd_sc_hd__mux4_1 _12465_ (.A0(\core_pipeline.pipeline_registers.registers[8][25] ),
    .A1(\core_pipeline.pipeline_registers.registers[9][25] ),
    .A2(\core_pipeline.pipeline_registers.registers[10][25] ),
    .A3(\core_pipeline.pipeline_registers.registers[11][25] ),
    .S0(net606),
    .S1(net584),
    .X(_02774_));
 sky130_fd_sc_hd__mux4_1 _12466_ (.A0(\core_pipeline.pipeline_registers.registers[12][25] ),
    .A1(\core_pipeline.pipeline_registers.registers[13][25] ),
    .A2(\core_pipeline.pipeline_registers.registers[14][25] ),
    .A3(\core_pipeline.pipeline_registers.registers[15][25] ),
    .S0(net612),
    .S1(net590),
    .X(_02775_));
 sky130_fd_sc_hd__or2_1 _12467_ (.A(net475),
    .B(_02775_),
    .X(_02776_));
 sky130_fd_sc_hd__o21a_1 _12468_ (.A1(net577),
    .A2(_02774_),
    .B1(net570),
    .X(_02777_));
 sky130_fd_sc_hd__a221o_1 _12469_ (.A1(net469),
    .A2(_02773_),
    .B1(_02776_),
    .B2(_02777_),
    .C1(net569),
    .X(_02778_));
 sky130_fd_sc_hd__mux2_1 _12470_ (.A0(\core_pipeline.pipeline_registers.registers[30][25] ),
    .A1(\core_pipeline.pipeline_registers.registers[31][25] ),
    .S(net611),
    .X(_02779_));
 sky130_fd_sc_hd__and2_1 _12471_ (.A(net585),
    .B(_02779_),
    .X(_02780_));
 sky130_fd_sc_hd__mux2_1 _12472_ (.A0(\core_pipeline.pipeline_registers.registers[28][25] ),
    .A1(\core_pipeline.pipeline_registers.registers[29][25] ),
    .S(net606),
    .X(_02781_));
 sky130_fd_sc_hd__a21o_1 _12473_ (.A1(net483),
    .A2(_02781_),
    .B1(net475),
    .X(_02782_));
 sky130_fd_sc_hd__mux2_1 _12474_ (.A0(\core_pipeline.pipeline_registers.registers[26][25] ),
    .A1(\core_pipeline.pipeline_registers.registers[27][25] ),
    .S(net605),
    .X(_02783_));
 sky130_fd_sc_hd__and2_1 _12475_ (.A(net585),
    .B(_02783_),
    .X(_02784_));
 sky130_fd_sc_hd__mux2_1 _12476_ (.A0(\core_pipeline.pipeline_registers.registers[24][25] ),
    .A1(\core_pipeline.pipeline_registers.registers[25][25] ),
    .S(net605),
    .X(_02785_));
 sky130_fd_sc_hd__a21o_1 _12477_ (.A1(net483),
    .A2(_02785_),
    .B1(net576),
    .X(_02786_));
 sky130_fd_sc_hd__o221a_1 _12478_ (.A1(_02780_),
    .A2(_02782_),
    .B1(_02784_),
    .B2(_02786_),
    .C1(net570),
    .X(_02787_));
 sky130_fd_sc_hd__mux2_1 _12479_ (.A0(_02771_),
    .A1(_02772_),
    .S(net475),
    .X(_02788_));
 sky130_fd_sc_hd__a211o_1 _12480_ (.A1(net469),
    .A2(_02788_),
    .B1(_02787_),
    .C1(net467),
    .X(_02789_));
 sky130_fd_sc_hd__and3_1 _12481_ (.A(net139),
    .B(_02778_),
    .C(_02789_),
    .X(_02790_));
 sky130_fd_sc_hd__a21o_1 _12482_ (.A1(\core_pipeline.decode_to_execute_rs1_data[25] ),
    .A2(net121),
    .B1(_02790_),
    .X(_01946_));
 sky130_fd_sc_hd__mux4_1 _12483_ (.A0(\core_pipeline.pipeline_registers.registers[4][26] ),
    .A1(\core_pipeline.pipeline_registers.registers[5][26] ),
    .A2(\core_pipeline.pipeline_registers.registers[6][26] ),
    .A3(\core_pipeline.pipeline_registers.registers[7][26] ),
    .S0(net612),
    .S1(net590),
    .X(_02791_));
 sky130_fd_sc_hd__mux4_1 _12484_ (.A0(\core_pipeline.pipeline_registers.registers[0][26] ),
    .A1(\core_pipeline.pipeline_registers.registers[1][26] ),
    .A2(\core_pipeline.pipeline_registers.registers[2][26] ),
    .A3(\core_pipeline.pipeline_registers.registers[3][26] ),
    .S0(net612),
    .S1(net590),
    .X(_02792_));
 sky130_fd_sc_hd__mux4_1 _12485_ (.A0(\core_pipeline.pipeline_registers.registers[20][26] ),
    .A1(\core_pipeline.pipeline_registers.registers[21][26] ),
    .A2(\core_pipeline.pipeline_registers.registers[22][26] ),
    .A3(\core_pipeline.pipeline_registers.registers[23][26] ),
    .S0(net613),
    .S1(net591),
    .X(_02793_));
 sky130_fd_sc_hd__mux4_1 _12486_ (.A0(\core_pipeline.pipeline_registers.registers[16][26] ),
    .A1(\core_pipeline.pipeline_registers.registers[17][26] ),
    .A2(\core_pipeline.pipeline_registers.registers[18][26] ),
    .A3(\core_pipeline.pipeline_registers.registers[19][26] ),
    .S0(net613),
    .S1(net591),
    .X(_02794_));
 sky130_fd_sc_hd__mux2_1 _12487_ (.A0(_02791_),
    .A1(_02792_),
    .S(net475),
    .X(_02795_));
 sky130_fd_sc_hd__mux4_1 _12488_ (.A0(\core_pipeline.pipeline_registers.registers[8][26] ),
    .A1(\core_pipeline.pipeline_registers.registers[9][26] ),
    .A2(\core_pipeline.pipeline_registers.registers[10][26] ),
    .A3(\core_pipeline.pipeline_registers.registers[11][26] ),
    .S0(net612),
    .S1(net590),
    .X(_02796_));
 sky130_fd_sc_hd__mux4_1 _12489_ (.A0(\core_pipeline.pipeline_registers.registers[12][26] ),
    .A1(\core_pipeline.pipeline_registers.registers[13][26] ),
    .A2(\core_pipeline.pipeline_registers.registers[14][26] ),
    .A3(\core_pipeline.pipeline_registers.registers[15][26] ),
    .S0(net612),
    .S1(net590),
    .X(_02797_));
 sky130_fd_sc_hd__or2_1 _12490_ (.A(net475),
    .B(_02797_),
    .X(_02798_));
 sky130_fd_sc_hd__o21a_1 _12491_ (.A1(net578),
    .A2(_02796_),
    .B1(net572),
    .X(_02799_));
 sky130_fd_sc_hd__a221o_1 _12492_ (.A1(net469),
    .A2(_02795_),
    .B1(_02798_),
    .B2(_02799_),
    .C1(net567),
    .X(_02800_));
 sky130_fd_sc_hd__mux2_1 _12493_ (.A0(\core_pipeline.pipeline_registers.registers[30][26] ),
    .A1(\core_pipeline.pipeline_registers.registers[31][26] ),
    .S(net613),
    .X(_02801_));
 sky130_fd_sc_hd__and2_1 _12494_ (.A(net585),
    .B(_02801_),
    .X(_02802_));
 sky130_fd_sc_hd__mux2_1 _12495_ (.A0(\core_pipeline.pipeline_registers.registers[28][26] ),
    .A1(\core_pipeline.pipeline_registers.registers[29][26] ),
    .S(net613),
    .X(_02803_));
 sky130_fd_sc_hd__a21o_1 _12496_ (.A1(net482),
    .A2(_02803_),
    .B1(net475),
    .X(_02804_));
 sky130_fd_sc_hd__mux2_1 _12497_ (.A0(\core_pipeline.pipeline_registers.registers[26][26] ),
    .A1(\core_pipeline.pipeline_registers.registers[27][26] ),
    .S(net613),
    .X(_02805_));
 sky130_fd_sc_hd__and2_1 _12498_ (.A(net585),
    .B(_02805_),
    .X(_02806_));
 sky130_fd_sc_hd__mux2_1 _12499_ (.A0(\core_pipeline.pipeline_registers.registers[24][26] ),
    .A1(\core_pipeline.pipeline_registers.registers[25][26] ),
    .S(net613),
    .X(_02807_));
 sky130_fd_sc_hd__a21o_1 _12500_ (.A1(net482),
    .A2(_02807_),
    .B1(net576),
    .X(_02808_));
 sky130_fd_sc_hd__o221a_1 _12501_ (.A1(_02802_),
    .A2(_02804_),
    .B1(_02806_),
    .B2(_02808_),
    .C1(net570),
    .X(_02809_));
 sky130_fd_sc_hd__mux2_1 _12502_ (.A0(_02793_),
    .A1(_02794_),
    .S(net476),
    .X(_02810_));
 sky130_fd_sc_hd__a211o_1 _12503_ (.A1(net469),
    .A2(_02810_),
    .B1(_02809_),
    .C1(net467),
    .X(_02811_));
 sky130_fd_sc_hd__and3_1 _12504_ (.A(net140),
    .B(_02800_),
    .C(_02811_),
    .X(_02812_));
 sky130_fd_sc_hd__a21o_1 _12505_ (.A1(\core_pipeline.decode_to_execute_rs1_data[26] ),
    .A2(net122),
    .B1(_02812_),
    .X(_01947_));
 sky130_fd_sc_hd__mux4_1 _12506_ (.A0(\core_pipeline.pipeline_registers.registers[4][27] ),
    .A1(\core_pipeline.pipeline_registers.registers[5][27] ),
    .A2(\core_pipeline.pipeline_registers.registers[6][27] ),
    .A3(\core_pipeline.pipeline_registers.registers[7][27] ),
    .S0(net626),
    .S1(net601),
    .X(_02813_));
 sky130_fd_sc_hd__mux4_1 _12507_ (.A0(\core_pipeline.pipeline_registers.registers[0][27] ),
    .A1(\core_pipeline.pipeline_registers.registers[1][27] ),
    .A2(\core_pipeline.pipeline_registers.registers[2][27] ),
    .A3(\core_pipeline.pipeline_registers.registers[3][27] ),
    .S0(net624),
    .S1(net601),
    .X(_02814_));
 sky130_fd_sc_hd__mux4_1 _12508_ (.A0(\core_pipeline.pipeline_registers.registers[20][27] ),
    .A1(\core_pipeline.pipeline_registers.registers[21][27] ),
    .A2(\core_pipeline.pipeline_registers.registers[22][27] ),
    .A3(\core_pipeline.pipeline_registers.registers[23][27] ),
    .S0(net624),
    .S1(net601),
    .X(_02815_));
 sky130_fd_sc_hd__mux4_1 _12509_ (.A0(\core_pipeline.pipeline_registers.registers[16][27] ),
    .A1(\core_pipeline.pipeline_registers.registers[17][27] ),
    .A2(\core_pipeline.pipeline_registers.registers[18][27] ),
    .A3(\core_pipeline.pipeline_registers.registers[19][27] ),
    .S0(net624),
    .S1(net601),
    .X(_02816_));
 sky130_fd_sc_hd__mux2_1 _12510_ (.A0(_02813_),
    .A1(_02814_),
    .S(net479),
    .X(_02817_));
 sky130_fd_sc_hd__mux4_1 _12511_ (.A0(\core_pipeline.pipeline_registers.registers[8][27] ),
    .A1(\core_pipeline.pipeline_registers.registers[9][27] ),
    .A2(\core_pipeline.pipeline_registers.registers[10][27] ),
    .A3(\core_pipeline.pipeline_registers.registers[11][27] ),
    .S0(net624),
    .S1(net601),
    .X(_02818_));
 sky130_fd_sc_hd__mux4_1 _12512_ (.A0(\core_pipeline.pipeline_registers.registers[12][27] ),
    .A1(\core_pipeline.pipeline_registers.registers[13][27] ),
    .A2(\core_pipeline.pipeline_registers.registers[14][27] ),
    .A3(\core_pipeline.pipeline_registers.registers[15][27] ),
    .S0(net624),
    .S1(net601),
    .X(_02819_));
 sky130_fd_sc_hd__or2_1 _12513_ (.A(net479),
    .B(_02819_),
    .X(_02820_));
 sky130_fd_sc_hd__o21a_1 _12514_ (.A1(net581),
    .A2(_02818_),
    .B1(net575),
    .X(_02821_));
 sky130_fd_sc_hd__a221o_1 _12515_ (.A1(net471),
    .A2(_02817_),
    .B1(_02820_),
    .B2(_02821_),
    .C1(net569),
    .X(_02822_));
 sky130_fd_sc_hd__mux2_1 _12516_ (.A0(\core_pipeline.pipeline_registers.registers[30][27] ),
    .A1(\core_pipeline.pipeline_registers.registers[31][27] ),
    .S(net624),
    .X(_02823_));
 sky130_fd_sc_hd__and2_1 _12517_ (.A(net601),
    .B(_02823_),
    .X(_02824_));
 sky130_fd_sc_hd__mux2_1 _12518_ (.A0(\core_pipeline.pipeline_registers.registers[28][27] ),
    .A1(\core_pipeline.pipeline_registers.registers[29][27] ),
    .S(net625),
    .X(_02825_));
 sky130_fd_sc_hd__a21o_1 _12519_ (.A1(net485),
    .A2(_02825_),
    .B1(net479),
    .X(_02826_));
 sky130_fd_sc_hd__mux2_1 _12520_ (.A0(\core_pipeline.pipeline_registers.registers[26][27] ),
    .A1(\core_pipeline.pipeline_registers.registers[27][27] ),
    .S(net624),
    .X(_02827_));
 sky130_fd_sc_hd__and2_1 _12521_ (.A(net601),
    .B(_02827_),
    .X(_02828_));
 sky130_fd_sc_hd__mux2_1 _12522_ (.A0(\core_pipeline.pipeline_registers.registers[24][27] ),
    .A1(\core_pipeline.pipeline_registers.registers[25][27] ),
    .S(net624),
    .X(_02829_));
 sky130_fd_sc_hd__a21o_1 _12523_ (.A1(net485),
    .A2(_02829_),
    .B1(net581),
    .X(_02830_));
 sky130_fd_sc_hd__o221a_1 _12524_ (.A1(_02824_),
    .A2(_02826_),
    .B1(_02828_),
    .B2(_02830_),
    .C1(net575),
    .X(_02831_));
 sky130_fd_sc_hd__mux2_1 _12525_ (.A0(_02815_),
    .A1(_02816_),
    .S(net479),
    .X(_02832_));
 sky130_fd_sc_hd__a211o_1 _12526_ (.A1(net471),
    .A2(_02832_),
    .B1(_02831_),
    .C1(net466),
    .X(_02833_));
 sky130_fd_sc_hd__and3_1 _12527_ (.A(net146),
    .B(_02822_),
    .C(_02833_),
    .X(_02834_));
 sky130_fd_sc_hd__a21o_1 _12528_ (.A1(\core_pipeline.decode_to_execute_rs1_data[27] ),
    .A2(net134),
    .B1(_02834_),
    .X(_01948_));
 sky130_fd_sc_hd__mux4_1 _12529_ (.A0(\core_pipeline.pipeline_registers.registers[4][28] ),
    .A1(\core_pipeline.pipeline_registers.registers[5][28] ),
    .A2(\core_pipeline.pipeline_registers.registers[6][28] ),
    .A3(\core_pipeline.pipeline_registers.registers[7][28] ),
    .S0(net622),
    .S1(net599),
    .X(_02835_));
 sky130_fd_sc_hd__mux4_1 _12530_ (.A0(\core_pipeline.pipeline_registers.registers[0][28] ),
    .A1(\core_pipeline.pipeline_registers.registers[1][28] ),
    .A2(\core_pipeline.pipeline_registers.registers[2][28] ),
    .A3(\core_pipeline.pipeline_registers.registers[3][28] ),
    .S0(net622),
    .S1(net599),
    .X(_02836_));
 sky130_fd_sc_hd__mux4_1 _12531_ (.A0(\core_pipeline.pipeline_registers.registers[20][28] ),
    .A1(\core_pipeline.pipeline_registers.registers[21][28] ),
    .A2(\core_pipeline.pipeline_registers.registers[22][28] ),
    .A3(\core_pipeline.pipeline_registers.registers[23][28] ),
    .S0(net622),
    .S1(net599),
    .X(_02837_));
 sky130_fd_sc_hd__mux4_1 _12532_ (.A0(\core_pipeline.pipeline_registers.registers[16][28] ),
    .A1(\core_pipeline.pipeline_registers.registers[17][28] ),
    .A2(\core_pipeline.pipeline_registers.registers[18][28] ),
    .A3(\core_pipeline.pipeline_registers.registers[19][28] ),
    .S0(net622),
    .S1(net598),
    .X(_02838_));
 sky130_fd_sc_hd__mux2_1 _12533_ (.A0(_02835_),
    .A1(_02836_),
    .S(net481),
    .X(_02839_));
 sky130_fd_sc_hd__mux4_1 _12534_ (.A0(\core_pipeline.pipeline_registers.registers[8][28] ),
    .A1(\core_pipeline.pipeline_registers.registers[9][28] ),
    .A2(\core_pipeline.pipeline_registers.registers[10][28] ),
    .A3(\core_pipeline.pipeline_registers.registers[11][28] ),
    .S0(net622),
    .S1(net599),
    .X(_02840_));
 sky130_fd_sc_hd__mux4_1 _12535_ (.A0(\core_pipeline.pipeline_registers.registers[12][28] ),
    .A1(\core_pipeline.pipeline_registers.registers[13][28] ),
    .A2(\core_pipeline.pipeline_registers.registers[14][28] ),
    .A3(\core_pipeline.pipeline_registers.registers[15][28] ),
    .S0(net622),
    .S1(net599),
    .X(_02841_));
 sky130_fd_sc_hd__or2_1 _12536_ (.A(net478),
    .B(_02841_),
    .X(_02842_));
 sky130_fd_sc_hd__o21a_1 _12537_ (.A1(net580),
    .A2(_02840_),
    .B1(net574),
    .X(_02843_));
 sky130_fd_sc_hd__a221o_1 _12538_ (.A1(net470),
    .A2(_02839_),
    .B1(_02842_),
    .B2(_02843_),
    .C1(net568),
    .X(_02844_));
 sky130_fd_sc_hd__mux2_1 _12539_ (.A0(\core_pipeline.pipeline_registers.registers[30][28] ),
    .A1(\core_pipeline.pipeline_registers.registers[31][28] ),
    .S(net620),
    .X(_02845_));
 sky130_fd_sc_hd__and2_1 _12540_ (.A(net597),
    .B(_02845_),
    .X(_02846_));
 sky130_fd_sc_hd__mux2_1 _12541_ (.A0(\core_pipeline.pipeline_registers.registers[28][28] ),
    .A1(\core_pipeline.pipeline_registers.registers[29][28] ),
    .S(net620),
    .X(_02847_));
 sky130_fd_sc_hd__a21o_1 _12542_ (.A1(net484),
    .A2(_02847_),
    .B1(net478),
    .X(_02848_));
 sky130_fd_sc_hd__mux2_1 _12543_ (.A0(\core_pipeline.pipeline_registers.registers[26][28] ),
    .A1(\core_pipeline.pipeline_registers.registers[27][28] ),
    .S(net619),
    .X(_02849_));
 sky130_fd_sc_hd__and2_1 _12544_ (.A(net596),
    .B(_02849_),
    .X(_02850_));
 sky130_fd_sc_hd__mux2_1 _12545_ (.A0(\core_pipeline.pipeline_registers.registers[24][28] ),
    .A1(\core_pipeline.pipeline_registers.registers[25][28] ),
    .S(net623),
    .X(_02851_));
 sky130_fd_sc_hd__a21o_1 _12546_ (.A1(net485),
    .A2(_02851_),
    .B1(net580),
    .X(_02852_));
 sky130_fd_sc_hd__o221a_1 _12547_ (.A1(_02846_),
    .A2(_02848_),
    .B1(_02850_),
    .B2(_02852_),
    .C1(net574),
    .X(_02853_));
 sky130_fd_sc_hd__mux2_1 _12548_ (.A0(_02837_),
    .A1(_02838_),
    .S(net481),
    .X(_02854_));
 sky130_fd_sc_hd__a211o_1 _12549_ (.A1(net471),
    .A2(_02854_),
    .B1(_02853_),
    .C1(net466),
    .X(_02855_));
 sky130_fd_sc_hd__and3_1 _12550_ (.A(net145),
    .B(_02844_),
    .C(_02855_),
    .X(_02856_));
 sky130_fd_sc_hd__a21o_1 _12551_ (.A1(\core_pipeline.decode_to_execute_rs1_data[28] ),
    .A2(net135),
    .B1(_02856_),
    .X(_01949_));
 sky130_fd_sc_hd__mux4_1 _12552_ (.A0(\core_pipeline.pipeline_registers.registers[4][29] ),
    .A1(\core_pipeline.pipeline_registers.registers[5][29] ),
    .A2(\core_pipeline.pipeline_registers.registers[6][29] ),
    .A3(\core_pipeline.pipeline_registers.registers[7][29] ),
    .S0(net617),
    .S1(net595),
    .X(_02857_));
 sky130_fd_sc_hd__mux4_1 _12553_ (.A0(\core_pipeline.pipeline_registers.registers[0][29] ),
    .A1(\core_pipeline.pipeline_registers.registers[1][29] ),
    .A2(\core_pipeline.pipeline_registers.registers[2][29] ),
    .A3(\core_pipeline.pipeline_registers.registers[3][29] ),
    .S0(net617),
    .S1(net595),
    .X(_02858_));
 sky130_fd_sc_hd__mux4_1 _12554_ (.A0(\core_pipeline.pipeline_registers.registers[20][29] ),
    .A1(\core_pipeline.pipeline_registers.registers[21][29] ),
    .A2(\core_pipeline.pipeline_registers.registers[22][29] ),
    .A3(\core_pipeline.pipeline_registers.registers[23][29] ),
    .S0(net618),
    .S1(net595),
    .X(_02859_));
 sky130_fd_sc_hd__mux4_1 _12555_ (.A0(\core_pipeline.pipeline_registers.registers[16][29] ),
    .A1(\core_pipeline.pipeline_registers.registers[17][29] ),
    .A2(\core_pipeline.pipeline_registers.registers[18][29] ),
    .A3(\core_pipeline.pipeline_registers.registers[19][29] ),
    .S0(net618),
    .S1(net595),
    .X(_02860_));
 sky130_fd_sc_hd__mux2_1 _12556_ (.A0(_02857_),
    .A1(_02858_),
    .S(net480),
    .X(_02861_));
 sky130_fd_sc_hd__mux4_1 _12557_ (.A0(\core_pipeline.pipeline_registers.registers[8][29] ),
    .A1(\core_pipeline.pipeline_registers.registers[9][29] ),
    .A2(\core_pipeline.pipeline_registers.registers[10][29] ),
    .A3(\core_pipeline.pipeline_registers.registers[11][29] ),
    .S0(net618),
    .S1(net595),
    .X(_02862_));
 sky130_fd_sc_hd__mux4_1 _12558_ (.A0(\core_pipeline.pipeline_registers.registers[12][29] ),
    .A1(\core_pipeline.pipeline_registers.registers[13][29] ),
    .A2(\core_pipeline.pipeline_registers.registers[14][29] ),
    .A3(\core_pipeline.pipeline_registers.registers[15][29] ),
    .S0(net618),
    .S1(net595),
    .X(_02863_));
 sky130_fd_sc_hd__or2_1 _12559_ (.A(net480),
    .B(_02863_),
    .X(_02864_));
 sky130_fd_sc_hd__o21a_1 _12560_ (.A1(net579),
    .A2(_02862_),
    .B1(net573),
    .X(_02865_));
 sky130_fd_sc_hd__a221o_1 _12561_ (.A1(net471),
    .A2(_02861_),
    .B1(_02864_),
    .B2(_02865_),
    .C1(net568),
    .X(_02866_));
 sky130_fd_sc_hd__mux2_1 _12562_ (.A0(\core_pipeline.pipeline_registers.registers[30][29] ),
    .A1(\core_pipeline.pipeline_registers.registers[31][29] ),
    .S(net618),
    .X(_02867_));
 sky130_fd_sc_hd__and2_1 _12563_ (.A(net594),
    .B(_02867_),
    .X(_02868_));
 sky130_fd_sc_hd__mux2_1 _12564_ (.A0(\core_pipeline.pipeline_registers.registers[28][29] ),
    .A1(\core_pipeline.pipeline_registers.registers[29][29] ),
    .S(net618),
    .X(_02869_));
 sky130_fd_sc_hd__a21o_1 _12565_ (.A1(net484),
    .A2(_02869_),
    .B1(net477),
    .X(_02870_));
 sky130_fd_sc_hd__mux2_1 _12566_ (.A0(\core_pipeline.pipeline_registers.registers[26][29] ),
    .A1(\core_pipeline.pipeline_registers.registers[27][29] ),
    .S(net618),
    .X(_02871_));
 sky130_fd_sc_hd__and2_1 _12567_ (.A(net595),
    .B(_02871_),
    .X(_02872_));
 sky130_fd_sc_hd__mux2_1 _12568_ (.A0(\core_pipeline.pipeline_registers.registers[24][29] ),
    .A1(\core_pipeline.pipeline_registers.registers[25][29] ),
    .S(net618),
    .X(_02873_));
 sky130_fd_sc_hd__a21o_1 _12569_ (.A1(net484),
    .A2(_02873_),
    .B1(net579),
    .X(_02874_));
 sky130_fd_sc_hd__o221a_1 _12570_ (.A1(_02868_),
    .A2(_02870_),
    .B1(_02872_),
    .B2(_02874_),
    .C1(net573),
    .X(_02875_));
 sky130_fd_sc_hd__mux2_1 _12571_ (.A0(_02859_),
    .A1(_02860_),
    .S(net477),
    .X(_02876_));
 sky130_fd_sc_hd__a211o_1 _12572_ (.A1(net470),
    .A2(_02876_),
    .B1(_02875_),
    .C1(net466),
    .X(_02877_));
 sky130_fd_sc_hd__and3_1 _12573_ (.A(net145),
    .B(_02866_),
    .C(_02877_),
    .X(_02878_));
 sky130_fd_sc_hd__a21o_1 _12574_ (.A1(\core_pipeline.decode_to_execute_rs1_data[29] ),
    .A2(net131),
    .B1(_02878_),
    .X(_01950_));
 sky130_fd_sc_hd__mux4_1 _12575_ (.A0(\core_pipeline.pipeline_registers.registers[4][30] ),
    .A1(\core_pipeline.pipeline_registers.registers[5][30] ),
    .A2(\core_pipeline.pipeline_registers.registers[6][30] ),
    .A3(\core_pipeline.pipeline_registers.registers[7][30] ),
    .S0(net617),
    .S1(net594),
    .X(_02879_));
 sky130_fd_sc_hd__mux4_1 _12576_ (.A0(\core_pipeline.pipeline_registers.registers[0][30] ),
    .A1(\core_pipeline.pipeline_registers.registers[1][30] ),
    .A2(\core_pipeline.pipeline_registers.registers[2][30] ),
    .A3(\core_pipeline.pipeline_registers.registers[3][30] ),
    .S0(net617),
    .S1(net594),
    .X(_02880_));
 sky130_fd_sc_hd__mux4_1 _12577_ (.A0(\core_pipeline.pipeline_registers.registers[20][30] ),
    .A1(\core_pipeline.pipeline_registers.registers[21][30] ),
    .A2(\core_pipeline.pipeline_registers.registers[22][30] ),
    .A3(\core_pipeline.pipeline_registers.registers[23][30] ),
    .S0(net617),
    .S1(net594),
    .X(_02881_));
 sky130_fd_sc_hd__mux4_1 _12578_ (.A0(\core_pipeline.pipeline_registers.registers[16][30] ),
    .A1(\core_pipeline.pipeline_registers.registers[17][30] ),
    .A2(\core_pipeline.pipeline_registers.registers[18][30] ),
    .A3(\core_pipeline.pipeline_registers.registers[19][30] ),
    .S0(net617),
    .S1(net594),
    .X(_02882_));
 sky130_fd_sc_hd__mux2_1 _12579_ (.A0(_02879_),
    .A1(_02880_),
    .S(net477),
    .X(_02883_));
 sky130_fd_sc_hd__mux4_1 _12580_ (.A0(\core_pipeline.pipeline_registers.registers[8][30] ),
    .A1(\core_pipeline.pipeline_registers.registers[9][30] ),
    .A2(\core_pipeline.pipeline_registers.registers[10][30] ),
    .A3(\core_pipeline.pipeline_registers.registers[11][30] ),
    .S0(net615),
    .S1(net592),
    .X(_02884_));
 sky130_fd_sc_hd__mux4_1 _12581_ (.A0(\core_pipeline.pipeline_registers.registers[12][30] ),
    .A1(\core_pipeline.pipeline_registers.registers[13][30] ),
    .A2(\core_pipeline.pipeline_registers.registers[14][30] ),
    .A3(\core_pipeline.pipeline_registers.registers[15][30] ),
    .S0(net610),
    .S1(net588),
    .X(_02885_));
 sky130_fd_sc_hd__or2_1 _12582_ (.A(net473),
    .B(_02885_),
    .X(_02886_));
 sky130_fd_sc_hd__o21a_1 _12583_ (.A1(net579),
    .A2(_02884_),
    .B1(net573),
    .X(_02887_));
 sky130_fd_sc_hd__a221o_1 _12584_ (.A1(net470),
    .A2(_02883_),
    .B1(_02886_),
    .B2(_02887_),
    .C1(net568),
    .X(_02888_));
 sky130_fd_sc_hd__mux2_1 _12585_ (.A0(\core_pipeline.pipeline_registers.registers[30][30] ),
    .A1(\core_pipeline.pipeline_registers.registers[31][30] ),
    .S(net615),
    .X(_02889_));
 sky130_fd_sc_hd__and2_1 _12586_ (.A(net592),
    .B(_02889_),
    .X(_02890_));
 sky130_fd_sc_hd__mux2_1 _12587_ (.A0(\core_pipeline.pipeline_registers.registers[28][30] ),
    .A1(\core_pipeline.pipeline_registers.registers[29][30] ),
    .S(net615),
    .X(_02891_));
 sky130_fd_sc_hd__a21o_1 _12588_ (.A1(net484),
    .A2(_02891_),
    .B1(net481),
    .X(_02892_));
 sky130_fd_sc_hd__mux2_1 _12589_ (.A0(\core_pipeline.pipeline_registers.registers[26][30] ),
    .A1(\core_pipeline.pipeline_registers.registers[27][30] ),
    .S(net615),
    .X(_02893_));
 sky130_fd_sc_hd__and2_1 _12590_ (.A(net592),
    .B(_02893_),
    .X(_02894_));
 sky130_fd_sc_hd__mux2_1 _12591_ (.A0(\core_pipeline.pipeline_registers.registers[24][30] ),
    .A1(\core_pipeline.pipeline_registers.registers[25][30] ),
    .S(net615),
    .X(_02895_));
 sky130_fd_sc_hd__a21o_1 _12592_ (.A1(net484),
    .A2(_02895_),
    .B1(net579),
    .X(_02896_));
 sky130_fd_sc_hd__o221a_1 _12593_ (.A1(_02890_),
    .A2(_02892_),
    .B1(_02894_),
    .B2(_02896_),
    .C1(net573),
    .X(_02897_));
 sky130_fd_sc_hd__mux2_1 _12594_ (.A0(_02881_),
    .A1(_02882_),
    .S(net477),
    .X(_02898_));
 sky130_fd_sc_hd__a211o_1 _12595_ (.A1(net470),
    .A2(_02898_),
    .B1(_02897_),
    .C1(net466),
    .X(_02899_));
 sky130_fd_sc_hd__and3_1 _12596_ (.A(net144),
    .B(_02888_),
    .C(_02899_),
    .X(_02900_));
 sky130_fd_sc_hd__a21o_1 _12597_ (.A1(\core_pipeline.decode_to_execute_rs1_data[30] ),
    .A2(net125),
    .B1(_02900_),
    .X(_01951_));
 sky130_fd_sc_hd__mux4_1 _12598_ (.A0(\core_pipeline.pipeline_registers.registers[4][31] ),
    .A1(\core_pipeline.pipeline_registers.registers[5][31] ),
    .A2(\core_pipeline.pipeline_registers.registers[6][31] ),
    .A3(\core_pipeline.pipeline_registers.registers[7][31] ),
    .S0(net625),
    .S1(net598),
    .X(_02901_));
 sky130_fd_sc_hd__mux4_1 _12599_ (.A0(\core_pipeline.pipeline_registers.registers[0][31] ),
    .A1(\core_pipeline.pipeline_registers.registers[1][31] ),
    .A2(\core_pipeline.pipeline_registers.registers[2][31] ),
    .A3(\core_pipeline.pipeline_registers.registers[3][31] ),
    .S0(net624),
    .S1(net601),
    .X(_02902_));
 sky130_fd_sc_hd__mux4_1 _12600_ (.A0(\core_pipeline.pipeline_registers.registers[20][31] ),
    .A1(\core_pipeline.pipeline_registers.registers[21][31] ),
    .A2(\core_pipeline.pipeline_registers.registers[22][31] ),
    .A3(\core_pipeline.pipeline_registers.registers[23][31] ),
    .S0(net622),
    .S1(net599),
    .X(_02903_));
 sky130_fd_sc_hd__mux4_1 _12601_ (.A0(\core_pipeline.pipeline_registers.registers[16][31] ),
    .A1(\core_pipeline.pipeline_registers.registers[17][31] ),
    .A2(\core_pipeline.pipeline_registers.registers[18][31] ),
    .A3(\core_pipeline.pipeline_registers.registers[19][31] ),
    .S0(net622),
    .S1(net599),
    .X(_02904_));
 sky130_fd_sc_hd__mux2_1 _12602_ (.A0(_02901_),
    .A1(_02902_),
    .S(net479),
    .X(_02905_));
 sky130_fd_sc_hd__mux4_1 _12603_ (.A0(\core_pipeline.pipeline_registers.registers[8][31] ),
    .A1(\core_pipeline.pipeline_registers.registers[9][31] ),
    .A2(\core_pipeline.pipeline_registers.registers[10][31] ),
    .A3(\core_pipeline.pipeline_registers.registers[11][31] ),
    .S0(net622),
    .S1(net599),
    .X(_02906_));
 sky130_fd_sc_hd__mux4_1 _12604_ (.A0(\core_pipeline.pipeline_registers.registers[12][31] ),
    .A1(\core_pipeline.pipeline_registers.registers[13][31] ),
    .A2(\core_pipeline.pipeline_registers.registers[14][31] ),
    .A3(\core_pipeline.pipeline_registers.registers[15][31] ),
    .S0(net625),
    .S1(net599),
    .X(_02907_));
 sky130_fd_sc_hd__or2_1 _12605_ (.A(net479),
    .B(_02907_),
    .X(_02908_));
 sky130_fd_sc_hd__o21a_1 _12606_ (.A1(net580),
    .A2(_02906_),
    .B1(net574),
    .X(_02909_));
 sky130_fd_sc_hd__a221o_1 _12607_ (.A1(net471),
    .A2(_02905_),
    .B1(_02908_),
    .B2(_02909_),
    .C1(net568),
    .X(_02910_));
 sky130_fd_sc_hd__mux2_1 _12608_ (.A0(\core_pipeline.pipeline_registers.registers[30][31] ),
    .A1(\core_pipeline.pipeline_registers.registers[31][31] ),
    .S(net622),
    .X(_02911_));
 sky130_fd_sc_hd__and2_1 _12609_ (.A(net599),
    .B(_02911_),
    .X(_02912_));
 sky130_fd_sc_hd__mux2_1 _12610_ (.A0(\core_pipeline.pipeline_registers.registers[28][31] ),
    .A1(\core_pipeline.pipeline_registers.registers[29][31] ),
    .S(net622),
    .X(_02913_));
 sky130_fd_sc_hd__a21o_1 _12611_ (.A1(net485),
    .A2(_02913_),
    .B1(net479),
    .X(_02914_));
 sky130_fd_sc_hd__mux2_1 _12612_ (.A0(\core_pipeline.pipeline_registers.registers[26][31] ),
    .A1(\core_pipeline.pipeline_registers.registers[27][31] ),
    .S(net622),
    .X(_02915_));
 sky130_fd_sc_hd__and2_1 _12613_ (.A(net599),
    .B(_02915_),
    .X(_02916_));
 sky130_fd_sc_hd__mux2_1 _12614_ (.A0(\core_pipeline.pipeline_registers.registers[24][31] ),
    .A1(\core_pipeline.pipeline_registers.registers[25][31] ),
    .S(net621),
    .X(_02917_));
 sky130_fd_sc_hd__a21o_1 _12615_ (.A1(net485),
    .A2(_02917_),
    .B1(net580),
    .X(_02918_));
 sky130_fd_sc_hd__o221a_1 _12616_ (.A1(_02912_),
    .A2(_02914_),
    .B1(_02916_),
    .B2(_02918_),
    .C1(net574),
    .X(_02919_));
 sky130_fd_sc_hd__mux2_1 _12617_ (.A0(_02903_),
    .A1(_02904_),
    .S(net479),
    .X(_02920_));
 sky130_fd_sc_hd__a211o_1 _12618_ (.A1(net471),
    .A2(_02920_),
    .B1(_02919_),
    .C1(net466),
    .X(_02921_));
 sky130_fd_sc_hd__and3_1 _12619_ (.A(net146),
    .B(_02910_),
    .C(_02921_),
    .X(_02922_));
 sky130_fd_sc_hd__a21o_1 _12620_ (.A1(\core_pipeline.decode_to_execute_rs1_data[31] ),
    .A2(net135),
    .B1(_02922_),
    .X(_01952_));
 sky130_fd_sc_hd__nor2_4 _12621_ (.A(_03516_),
    .B(_00004_),
    .Y(_02923_));
 sky130_fd_sc_hd__or2_2 _12622_ (.A(_03516_),
    .B(_00004_),
    .X(_02924_));
 sky130_fd_sc_hd__nand2_1 _12623_ (.A(\core_pipeline.pipeline_fetch.pc[2] ),
    .B(net351),
    .Y(_02925_));
 sky130_fd_sc_hd__o211a_1 _12624_ (.A1(\core_busio.mem_address[2] ),
    .A2(net351),
    .B1(net445),
    .C1(_02925_),
    .X(_02926_));
 sky130_fd_sc_hd__a211o_1 _12625_ (.A1(\core_pipeline.csr_to_fetch_mret_vector[2] ),
    .A2(_03512_),
    .B1(_02926_),
    .C1(_03479_),
    .X(_02927_));
 sky130_fd_sc_hd__o21ai_1 _12626_ (.A1(\core_pipeline.csr_to_fetch_trap_vector[2] ),
    .A2(net400),
    .B1(_02927_),
    .Y(_02928_));
 sky130_fd_sc_hd__nand2_1 _12627_ (.A(net104),
    .B(_02928_),
    .Y(_02929_));
 sky130_fd_sc_hd__o211a_1 _12628_ (.A1(\core_pipeline.pipeline_fetch.pc[2] ),
    .A2(net104),
    .B1(_02929_),
    .C1(net638),
    .X(_01953_));
 sky130_fd_sc_hd__xor2_1 _12629_ (.A(\core_pipeline.pipeline_fetch.pc[3] ),
    .B(\core_pipeline.pipeline_fetch.pc[2] ),
    .X(_02930_));
 sky130_fd_sc_hd__mux2_1 _12630_ (.A0(\core_busio.mem_address[3] ),
    .A1(_02930_),
    .S(net351),
    .X(_02931_));
 sky130_fd_sc_hd__mux2_1 _12631_ (.A0(\core_pipeline.csr_to_fetch_mret_vector[3] ),
    .A1(_02931_),
    .S(net445),
    .X(_02932_));
 sky130_fd_sc_hd__mux2_1 _12632_ (.A0(\core_pipeline.csr_to_fetch_trap_vector[3] ),
    .A1(_02932_),
    .S(net400),
    .X(_02933_));
 sky130_fd_sc_hd__or2_1 _12633_ (.A(net105),
    .B(_02933_),
    .X(_02934_));
 sky130_fd_sc_hd__o211a_1 _12634_ (.A1(\core_pipeline.pipeline_fetch.pc[3] ),
    .A2(net104),
    .B1(_02934_),
    .C1(net638),
    .X(_01954_));
 sky130_fd_sc_hd__and3_1 _12635_ (.A(\core_pipeline.pipeline_fetch.pc[4] ),
    .B(\core_pipeline.pipeline_fetch.pc[3] ),
    .C(\core_pipeline.pipeline_fetch.pc[2] ),
    .X(_02935_));
 sky130_fd_sc_hd__a21oi_1 _12636_ (.A1(\core_pipeline.pipeline_fetch.pc[3] ),
    .A2(\core_pipeline.pipeline_fetch.pc[2] ),
    .B1(\core_pipeline.pipeline_fetch.pc[4] ),
    .Y(_02936_));
 sky130_fd_sc_hd__nor2_1 _12637_ (.A(_02935_),
    .B(_02936_),
    .Y(_02937_));
 sky130_fd_sc_hd__mux2_1 _12638_ (.A0(\core_busio.mem_address[4] ),
    .A1(_02937_),
    .S(net351),
    .X(_02938_));
 sky130_fd_sc_hd__mux2_1 _12639_ (.A0(\core_pipeline.csr_to_fetch_mret_vector[4] ),
    .A1(_02938_),
    .S(net445),
    .X(_02939_));
 sky130_fd_sc_hd__mux2_1 _12640_ (.A0(\core_pipeline.csr_to_fetch_trap_vector[4] ),
    .A1(_02939_),
    .S(net400),
    .X(_02940_));
 sky130_fd_sc_hd__or2_1 _12641_ (.A(net105),
    .B(_02940_),
    .X(_02941_));
 sky130_fd_sc_hd__o211a_1 _12642_ (.A1(\core_pipeline.pipeline_fetch.pc[4] ),
    .A2(net104),
    .B1(_02941_),
    .C1(net638),
    .X(_01955_));
 sky130_fd_sc_hd__and2_2 _12643_ (.A(\core_pipeline.pipeline_fetch.pc[5] ),
    .B(_02935_),
    .X(_02942_));
 sky130_fd_sc_hd__nor2_1 _12644_ (.A(\core_pipeline.pipeline_fetch.pc[5] ),
    .B(_02935_),
    .Y(_02943_));
 sky130_fd_sc_hd__nor2_1 _12645_ (.A(_02942_),
    .B(_02943_),
    .Y(_02944_));
 sky130_fd_sc_hd__mux2_1 _12646_ (.A0(\core_busio.mem_address[5] ),
    .A1(_02944_),
    .S(net351),
    .X(_02945_));
 sky130_fd_sc_hd__or3_1 _12647_ (.A(\core_pipeline.csr_to_fetch_mret_vector[5] ),
    .B(_03479_),
    .C(net445),
    .X(_02946_));
 sky130_fd_sc_hd__o221a_1 _12648_ (.A1(\core_pipeline.csr_to_fetch_trap_vector[5] ),
    .A2(net400),
    .B1(_03515_),
    .B2(_02945_),
    .C1(_02946_),
    .X(_02947_));
 sky130_fd_sc_hd__or2_1 _12649_ (.A(net105),
    .B(_02947_),
    .X(_02948_));
 sky130_fd_sc_hd__o211a_1 _12650_ (.A1(\core_pipeline.pipeline_fetch.pc[5] ),
    .A2(net104),
    .B1(_02948_),
    .C1(net638),
    .X(_01956_));
 sky130_fd_sc_hd__xor2_1 _12651_ (.A(\core_pipeline.pipeline_fetch.pc[6] ),
    .B(_02942_),
    .X(_02949_));
 sky130_fd_sc_hd__mux2_1 _12652_ (.A0(\core_busio.mem_address[6] ),
    .A1(_02949_),
    .S(net351),
    .X(_02950_));
 sky130_fd_sc_hd__mux2_1 _12653_ (.A0(\core_pipeline.csr_to_fetch_mret_vector[6] ),
    .A1(_02950_),
    .S(net445),
    .X(_02951_));
 sky130_fd_sc_hd__mux2_1 _12654_ (.A0(\core_pipeline.csr_to_fetch_trap_vector[6] ),
    .A1(_02951_),
    .S(net401),
    .X(_02952_));
 sky130_fd_sc_hd__or2_1 _12655_ (.A(net105),
    .B(_02952_),
    .X(_02953_));
 sky130_fd_sc_hd__o211a_1 _12656_ (.A1(\core_pipeline.pipeline_fetch.pc[6] ),
    .A2(net104),
    .B1(_02953_),
    .C1(net638),
    .X(_01957_));
 sky130_fd_sc_hd__and3_2 _12657_ (.A(\core_pipeline.pipeline_fetch.pc[7] ),
    .B(\core_pipeline.pipeline_fetch.pc[6] ),
    .C(_02942_),
    .X(_02954_));
 sky130_fd_sc_hd__a21oi_1 _12658_ (.A1(\core_pipeline.pipeline_fetch.pc[6] ),
    .A2(_02942_),
    .B1(\core_pipeline.pipeline_fetch.pc[7] ),
    .Y(_02955_));
 sky130_fd_sc_hd__nor2_1 _12659_ (.A(_02954_),
    .B(_02955_),
    .Y(_02956_));
 sky130_fd_sc_hd__mux2_1 _12660_ (.A0(\core_busio.mem_address[7] ),
    .A1(_02956_),
    .S(net351),
    .X(_02957_));
 sky130_fd_sc_hd__mux2_1 _12661_ (.A0(\core_pipeline.csr_to_fetch_mret_vector[7] ),
    .A1(_02957_),
    .S(net445),
    .X(_02958_));
 sky130_fd_sc_hd__mux2_1 _12662_ (.A0(\core_pipeline.csr_to_fetch_trap_vector[7] ),
    .A1(_02958_),
    .S(net401),
    .X(_02959_));
 sky130_fd_sc_hd__or2_1 _12663_ (.A(net105),
    .B(_02959_),
    .X(_02960_));
 sky130_fd_sc_hd__o211a_1 _12664_ (.A1(\core_pipeline.pipeline_fetch.pc[7] ),
    .A2(net104),
    .B1(_02960_),
    .C1(net638),
    .X(_01958_));
 sky130_fd_sc_hd__and2_2 _12665_ (.A(\core_pipeline.pipeline_fetch.pc[8] ),
    .B(_02954_),
    .X(_02961_));
 sky130_fd_sc_hd__nor2_1 _12666_ (.A(\core_pipeline.pipeline_fetch.pc[8] ),
    .B(_02954_),
    .Y(_02962_));
 sky130_fd_sc_hd__nor2_1 _12667_ (.A(_02961_),
    .B(_02962_),
    .Y(_02963_));
 sky130_fd_sc_hd__mux2_1 _12668_ (.A0(\core_busio.mem_address[8] ),
    .A1(_02963_),
    .S(net350),
    .X(_02964_));
 sky130_fd_sc_hd__mux2_1 _12669_ (.A0(\core_pipeline.csr_to_fetch_mret_vector[8] ),
    .A1(_02964_),
    .S(_03513_),
    .X(_02965_));
 sky130_fd_sc_hd__mux2_1 _12670_ (.A0(\core_pipeline.csr_to_fetch_trap_vector[8] ),
    .A1(_02965_),
    .S(net403),
    .X(_02966_));
 sky130_fd_sc_hd__or2_1 _12671_ (.A(net105),
    .B(_02966_),
    .X(_02967_));
 sky130_fd_sc_hd__o211a_1 _12672_ (.A1(\core_pipeline.pipeline_fetch.pc[8] ),
    .A2(net104),
    .B1(_02967_),
    .C1(net638),
    .X(_01959_));
 sky130_fd_sc_hd__xor2_1 _12673_ (.A(\core_pipeline.pipeline_fetch.pc[9] ),
    .B(_02961_),
    .X(_02968_));
 sky130_fd_sc_hd__mux2_1 _12674_ (.A0(\core_busio.mem_address[9] ),
    .A1(_02968_),
    .S(net350),
    .X(_02969_));
 sky130_fd_sc_hd__mux2_1 _12675_ (.A0(\core_pipeline.csr_to_fetch_mret_vector[9] ),
    .A1(_02969_),
    .S(net445),
    .X(_02970_));
 sky130_fd_sc_hd__mux2_1 _12676_ (.A0(\core_pipeline.csr_to_fetch_trap_vector[9] ),
    .A1(_02970_),
    .S(net402),
    .X(_02971_));
 sky130_fd_sc_hd__or2_1 _12677_ (.A(net106),
    .B(_02971_),
    .X(_02972_));
 sky130_fd_sc_hd__o211a_1 _12678_ (.A1(\core_pipeline.pipeline_fetch.pc[9] ),
    .A2(net103),
    .B1(_02972_),
    .C1(net636),
    .X(_01960_));
 sky130_fd_sc_hd__and3_2 _12679_ (.A(\core_pipeline.pipeline_fetch.pc[10] ),
    .B(\core_pipeline.pipeline_fetch.pc[9] ),
    .C(_02961_),
    .X(_02973_));
 sky130_fd_sc_hd__a21oi_1 _12680_ (.A1(\core_pipeline.pipeline_fetch.pc[9] ),
    .A2(_02961_),
    .B1(\core_pipeline.pipeline_fetch.pc[10] ),
    .Y(_02974_));
 sky130_fd_sc_hd__nor2_1 _12681_ (.A(_02973_),
    .B(_02974_),
    .Y(_02975_));
 sky130_fd_sc_hd__mux2_1 _12682_ (.A0(\core_busio.mem_address[10] ),
    .A1(_02975_),
    .S(net350),
    .X(_02976_));
 sky130_fd_sc_hd__mux2_1 _12683_ (.A0(\core_pipeline.csr_to_fetch_mret_vector[10] ),
    .A1(_02976_),
    .S(net445),
    .X(_02977_));
 sky130_fd_sc_hd__mux2_1 _12684_ (.A0(\core_pipeline.csr_to_fetch_trap_vector[10] ),
    .A1(_02977_),
    .S(net402),
    .X(_02978_));
 sky130_fd_sc_hd__or2_1 _12685_ (.A(net106),
    .B(_02978_),
    .X(_02979_));
 sky130_fd_sc_hd__o211a_1 _12686_ (.A1(\core_pipeline.pipeline_fetch.pc[10] ),
    .A2(net103),
    .B1(_02979_),
    .C1(net636),
    .X(_01961_));
 sky130_fd_sc_hd__and2_2 _12687_ (.A(\core_pipeline.pipeline_fetch.pc[11] ),
    .B(_02973_),
    .X(_02980_));
 sky130_fd_sc_hd__nor2_1 _12688_ (.A(\core_pipeline.pipeline_fetch.pc[11] ),
    .B(_02973_),
    .Y(_02981_));
 sky130_fd_sc_hd__nor2_1 _12689_ (.A(_02980_),
    .B(_02981_),
    .Y(_02982_));
 sky130_fd_sc_hd__mux2_1 _12690_ (.A0(\core_busio.mem_address[11] ),
    .A1(_02982_),
    .S(net350),
    .X(_02983_));
 sky130_fd_sc_hd__mux2_1 _12691_ (.A0(\core_pipeline.csr_to_fetch_mret_vector[11] ),
    .A1(_02983_),
    .S(_03513_),
    .X(_02984_));
 sky130_fd_sc_hd__mux2_1 _12692_ (.A0(\core_pipeline.csr_to_fetch_trap_vector[11] ),
    .A1(_02984_),
    .S(net402),
    .X(_02985_));
 sky130_fd_sc_hd__or2_1 _12693_ (.A(net106),
    .B(_02985_),
    .X(_02986_));
 sky130_fd_sc_hd__o211a_1 _12694_ (.A1(\core_pipeline.pipeline_fetch.pc[11] ),
    .A2(net103),
    .B1(_02986_),
    .C1(net636),
    .X(_01962_));
 sky130_fd_sc_hd__xor2_2 _12695_ (.A(\core_pipeline.pipeline_fetch.pc[12] ),
    .B(_02980_),
    .X(_02987_));
 sky130_fd_sc_hd__mux2_1 _12696_ (.A0(\core_busio.mem_address[12] ),
    .A1(_02987_),
    .S(net350),
    .X(_02988_));
 sky130_fd_sc_hd__mux2_1 _12697_ (.A0(\core_pipeline.csr_to_fetch_mret_vector[12] ),
    .A1(_02988_),
    .S(_03513_),
    .X(_02989_));
 sky130_fd_sc_hd__mux2_1 _12698_ (.A0(\core_pipeline.csr_to_fetch_trap_vector[12] ),
    .A1(_02989_),
    .S(net402),
    .X(_02990_));
 sky130_fd_sc_hd__or2_1 _12699_ (.A(net106),
    .B(_02990_),
    .X(_02991_));
 sky130_fd_sc_hd__o211a_1 _12700_ (.A1(\core_pipeline.pipeline_fetch.pc[12] ),
    .A2(net103),
    .B1(_02991_),
    .C1(net636),
    .X(_01963_));
 sky130_fd_sc_hd__and3_1 _12701_ (.A(\core_pipeline.pipeline_fetch.pc[13] ),
    .B(\core_pipeline.pipeline_fetch.pc[12] ),
    .C(_02980_),
    .X(_02992_));
 sky130_fd_sc_hd__a31o_1 _12702_ (.A1(\core_pipeline.pipeline_fetch.pc[12] ),
    .A2(\core_pipeline.pipeline_fetch.pc[11] ),
    .A3(_02973_),
    .B1(\core_pipeline.pipeline_fetch.pc[13] ),
    .X(_02993_));
 sky130_fd_sc_hd__and2b_1 _12703_ (.A_N(_02992_),
    .B(_02993_),
    .X(_02994_));
 sky130_fd_sc_hd__mux2_1 _12704_ (.A0(\core_busio.mem_address[13] ),
    .A1(_02994_),
    .S(net350),
    .X(_02995_));
 sky130_fd_sc_hd__mux2_1 _12705_ (.A0(\core_pipeline.csr_to_fetch_mret_vector[13] ),
    .A1(_02995_),
    .S(_03513_),
    .X(_02996_));
 sky130_fd_sc_hd__mux2_1 _12706_ (.A0(\core_pipeline.csr_to_fetch_trap_vector[13] ),
    .A1(_02996_),
    .S(net402),
    .X(_02997_));
 sky130_fd_sc_hd__or2_1 _12707_ (.A(net106),
    .B(_02997_),
    .X(_02998_));
 sky130_fd_sc_hd__o211a_1 _12708_ (.A1(\core_pipeline.pipeline_fetch.pc[13] ),
    .A2(net103),
    .B1(_02998_),
    .C1(net636),
    .X(_01964_));
 sky130_fd_sc_hd__and2_1 _12709_ (.A(\core_pipeline.pipeline_fetch.pc[14] ),
    .B(_02992_),
    .X(_02999_));
 sky130_fd_sc_hd__or2_1 _12710_ (.A(\core_pipeline.pipeline_fetch.pc[14] ),
    .B(_02992_),
    .X(_03000_));
 sky130_fd_sc_hd__and2b_1 _12711_ (.A_N(_02999_),
    .B(_03000_),
    .X(_03001_));
 sky130_fd_sc_hd__mux2_1 _12712_ (.A0(\core_busio.mem_address[14] ),
    .A1(_03001_),
    .S(net350),
    .X(_03002_));
 sky130_fd_sc_hd__mux2_1 _12713_ (.A0(\core_pipeline.csr_to_fetch_mret_vector[14] ),
    .A1(_03002_),
    .S(net445),
    .X(_03003_));
 sky130_fd_sc_hd__mux2_1 _12714_ (.A0(\core_pipeline.csr_to_fetch_trap_vector[14] ),
    .A1(_03003_),
    .S(net402),
    .X(_03004_));
 sky130_fd_sc_hd__or2_1 _12715_ (.A(net106),
    .B(_03004_),
    .X(_03005_));
 sky130_fd_sc_hd__o211a_1 _12716_ (.A1(\core_pipeline.pipeline_fetch.pc[14] ),
    .A2(net103),
    .B1(_03005_),
    .C1(net636),
    .X(_01965_));
 sky130_fd_sc_hd__xor2_1 _12717_ (.A(\core_pipeline.pipeline_fetch.pc[15] ),
    .B(_02999_),
    .X(_03006_));
 sky130_fd_sc_hd__mux2_1 _12718_ (.A0(\core_busio.mem_address[15] ),
    .A1(_03006_),
    .S(net350),
    .X(_03007_));
 sky130_fd_sc_hd__mux2_1 _12719_ (.A0(\core_pipeline.csr_to_fetch_mret_vector[15] ),
    .A1(_03007_),
    .S(net445),
    .X(_03008_));
 sky130_fd_sc_hd__mux2_1 _12720_ (.A0(\core_pipeline.csr_to_fetch_trap_vector[15] ),
    .A1(_03008_),
    .S(net402),
    .X(_03009_));
 sky130_fd_sc_hd__or2_1 _12721_ (.A(net106),
    .B(_03009_),
    .X(_03010_));
 sky130_fd_sc_hd__o211a_1 _12722_ (.A1(\core_pipeline.pipeline_fetch.pc[15] ),
    .A2(net103),
    .B1(_03010_),
    .C1(net636),
    .X(_01966_));
 sky130_fd_sc_hd__and3_2 _12723_ (.A(\core_pipeline.pipeline_fetch.pc[16] ),
    .B(\core_pipeline.pipeline_fetch.pc[15] ),
    .C(_02999_),
    .X(_03011_));
 sky130_fd_sc_hd__a21oi_1 _12724_ (.A1(\core_pipeline.pipeline_fetch.pc[15] ),
    .A2(_02999_),
    .B1(\core_pipeline.pipeline_fetch.pc[16] ),
    .Y(_03012_));
 sky130_fd_sc_hd__nor2_1 _12725_ (.A(_03011_),
    .B(_03012_),
    .Y(_03013_));
 sky130_fd_sc_hd__mux2_1 _12726_ (.A0(\core_busio.mem_address[16] ),
    .A1(_03013_),
    .S(net350),
    .X(_03014_));
 sky130_fd_sc_hd__mux2_1 _12727_ (.A0(\core_pipeline.csr_to_fetch_mret_vector[16] ),
    .A1(_03014_),
    .S(_03513_),
    .X(_03015_));
 sky130_fd_sc_hd__mux2_1 _12728_ (.A0(\core_pipeline.csr_to_fetch_trap_vector[16] ),
    .A1(_03015_),
    .S(net402),
    .X(_03016_));
 sky130_fd_sc_hd__or2_1 _12729_ (.A(net106),
    .B(_03016_),
    .X(_03017_));
 sky130_fd_sc_hd__o211a_1 _12730_ (.A1(\core_pipeline.pipeline_fetch.pc[16] ),
    .A2(net103),
    .B1(_03017_),
    .C1(net636),
    .X(_01967_));
 sky130_fd_sc_hd__and2_2 _12731_ (.A(\core_pipeline.pipeline_fetch.pc[17] ),
    .B(_03011_),
    .X(_03018_));
 sky130_fd_sc_hd__nor2_1 _12732_ (.A(\core_pipeline.pipeline_fetch.pc[17] ),
    .B(_03011_),
    .Y(_03019_));
 sky130_fd_sc_hd__nor2_1 _12733_ (.A(_03018_),
    .B(_03019_),
    .Y(_03020_));
 sky130_fd_sc_hd__mux2_1 _12734_ (.A0(\core_busio.mem_address[17] ),
    .A1(_03020_),
    .S(net350),
    .X(_03021_));
 sky130_fd_sc_hd__mux2_1 _12735_ (.A0(\core_pipeline.csr_to_fetch_mret_vector[17] ),
    .A1(_03021_),
    .S(net445),
    .X(_03022_));
 sky130_fd_sc_hd__mux2_1 _12736_ (.A0(\core_pipeline.csr_to_fetch_trap_vector[17] ),
    .A1(_03022_),
    .S(net403),
    .X(_03023_));
 sky130_fd_sc_hd__or2_1 _12737_ (.A(net106),
    .B(_03023_),
    .X(_03024_));
 sky130_fd_sc_hd__o211a_1 _12738_ (.A1(\core_pipeline.pipeline_fetch.pc[17] ),
    .A2(net103),
    .B1(_03024_),
    .C1(net636),
    .X(_01968_));
 sky130_fd_sc_hd__xor2_1 _12739_ (.A(\core_pipeline.pipeline_fetch.pc[18] ),
    .B(_03018_),
    .X(_03025_));
 sky130_fd_sc_hd__mux2_1 _12740_ (.A0(\core_busio.mem_address[18] ),
    .A1(_03025_),
    .S(net350),
    .X(_03026_));
 sky130_fd_sc_hd__mux2_1 _12741_ (.A0(\core_pipeline.csr_to_fetch_mret_vector[18] ),
    .A1(_03026_),
    .S(net445),
    .X(_03027_));
 sky130_fd_sc_hd__mux2_1 _12742_ (.A0(\core_pipeline.csr_to_fetch_trap_vector[18] ),
    .A1(_03027_),
    .S(net403),
    .X(_03028_));
 sky130_fd_sc_hd__or2_1 _12743_ (.A(net105),
    .B(_03028_),
    .X(_03029_));
 sky130_fd_sc_hd__o211a_1 _12744_ (.A1(\core_pipeline.pipeline_fetch.pc[18] ),
    .A2(net104),
    .B1(_03029_),
    .C1(net637),
    .X(_01969_));
 sky130_fd_sc_hd__and3_1 _12745_ (.A(\core_pipeline.pipeline_fetch.pc[19] ),
    .B(\core_pipeline.pipeline_fetch.pc[18] ),
    .C(_03018_),
    .X(_03030_));
 sky130_fd_sc_hd__a21oi_1 _12746_ (.A1(\core_pipeline.pipeline_fetch.pc[18] ),
    .A2(_03018_),
    .B1(\core_pipeline.pipeline_fetch.pc[19] ),
    .Y(_03031_));
 sky130_fd_sc_hd__nor2_1 _12747_ (.A(_03030_),
    .B(_03031_),
    .Y(_03032_));
 sky130_fd_sc_hd__mux2_1 _12748_ (.A0(\core_busio.mem_address[19] ),
    .A1(_03032_),
    .S(net350),
    .X(_03033_));
 sky130_fd_sc_hd__mux2_1 _12749_ (.A0(\core_pipeline.csr_to_fetch_mret_vector[19] ),
    .A1(_03033_),
    .S(net445),
    .X(_03034_));
 sky130_fd_sc_hd__mux2_1 _12750_ (.A0(\core_pipeline.csr_to_fetch_trap_vector[19] ),
    .A1(_03034_),
    .S(net403),
    .X(_03035_));
 sky130_fd_sc_hd__or2_1 _12751_ (.A(\core_pipeline.pipeline_fetch.pc[19] ),
    .B(net103),
    .X(_03036_));
 sky130_fd_sc_hd__o211a_1 _12752_ (.A1(net105),
    .A2(_03035_),
    .B1(_03036_),
    .C1(net637),
    .X(_01970_));
 sky130_fd_sc_hd__and2_2 _12753_ (.A(\core_pipeline.pipeline_fetch.pc[20] ),
    .B(_03030_),
    .X(_03037_));
 sky130_fd_sc_hd__or2_1 _12754_ (.A(\core_pipeline.pipeline_fetch.pc[20] ),
    .B(_03030_),
    .X(_03038_));
 sky130_fd_sc_hd__and2b_1 _12755_ (.A_N(_03037_),
    .B(_03038_),
    .X(_03039_));
 sky130_fd_sc_hd__mux2_1 _12756_ (.A0(\core_busio.mem_address[20] ),
    .A1(_03039_),
    .S(net351),
    .X(_03040_));
 sky130_fd_sc_hd__mux2_1 _12757_ (.A0(\core_pipeline.csr_to_fetch_mret_vector[20] ),
    .A1(_03040_),
    .S(net445),
    .X(_03041_));
 sky130_fd_sc_hd__mux2_1 _12758_ (.A0(\core_pipeline.csr_to_fetch_trap_vector[20] ),
    .A1(_03041_),
    .S(net403),
    .X(_03042_));
 sky130_fd_sc_hd__or2_1 _12759_ (.A(\core_pipeline.pipeline_fetch.pc[20] ),
    .B(net104),
    .X(_03043_));
 sky130_fd_sc_hd__o211a_1 _12760_ (.A1(net105),
    .A2(_03042_),
    .B1(_03043_),
    .C1(net637),
    .X(_01971_));
 sky130_fd_sc_hd__xor2_1 _12761_ (.A(\core_pipeline.pipeline_fetch.pc[21] ),
    .B(_03037_),
    .X(_03044_));
 sky130_fd_sc_hd__mux2_1 _12762_ (.A0(\core_busio.mem_address[21] ),
    .A1(_03044_),
    .S(net350),
    .X(_03045_));
 sky130_fd_sc_hd__mux2_1 _12763_ (.A0(\core_pipeline.csr_to_fetch_mret_vector[21] ),
    .A1(_03045_),
    .S(_03513_),
    .X(_03046_));
 sky130_fd_sc_hd__mux2_1 _12764_ (.A0(\core_pipeline.csr_to_fetch_trap_vector[21] ),
    .A1(_03046_),
    .S(net403),
    .X(_03047_));
 sky130_fd_sc_hd__or2_1 _12765_ (.A(\core_pipeline.pipeline_fetch.pc[21] ),
    .B(net103),
    .X(_03048_));
 sky130_fd_sc_hd__o211a_1 _12766_ (.A1(net106),
    .A2(_03047_),
    .B1(_03048_),
    .C1(net637),
    .X(_01972_));
 sky130_fd_sc_hd__and3_1 _12767_ (.A(\core_pipeline.pipeline_fetch.pc[22] ),
    .B(\core_pipeline.pipeline_fetch.pc[21] ),
    .C(_03037_),
    .X(_03049_));
 sky130_fd_sc_hd__a21oi_1 _12768_ (.A1(\core_pipeline.pipeline_fetch.pc[21] ),
    .A2(_03037_),
    .B1(\core_pipeline.pipeline_fetch.pc[22] ),
    .Y(_03050_));
 sky130_fd_sc_hd__nor2_1 _12769_ (.A(_03049_),
    .B(_03050_),
    .Y(_03051_));
 sky130_fd_sc_hd__or2_1 _12770_ (.A(_03511_),
    .B(_03051_),
    .X(_03052_));
 sky130_fd_sc_hd__or2_1 _12771_ (.A(\core_busio.mem_address[22] ),
    .B(net351),
    .X(_03053_));
 sky130_fd_sc_hd__a221o_1 _12772_ (.A1(\core_pipeline.csr_to_fetch_trap_vector[22] ),
    .A2(_03479_),
    .B1(_04385_),
    .B2(\core_pipeline.csr_to_fetch_mret_vector[22] ),
    .C1(net105),
    .X(_03054_));
 sky130_fd_sc_hd__a31o_1 _12773_ (.A1(_03514_),
    .A2(_03052_),
    .A3(_03053_),
    .B1(_03054_),
    .X(_03055_));
 sky130_fd_sc_hd__o211a_1 _12774_ (.A1(\core_pipeline.pipeline_fetch.pc[22] ),
    .A2(net103),
    .B1(_03055_),
    .C1(net637),
    .X(_01973_));
 sky130_fd_sc_hd__and2_1 _12775_ (.A(\core_pipeline.pipeline_fetch.pc[23] ),
    .B(_03049_),
    .X(_03056_));
 sky130_fd_sc_hd__or2_1 _12776_ (.A(\core_pipeline.pipeline_fetch.pc[23] ),
    .B(_03049_),
    .X(_03057_));
 sky130_fd_sc_hd__and2b_1 _12777_ (.A_N(_03056_),
    .B(_03057_),
    .X(_03058_));
 sky130_fd_sc_hd__or2_1 _12778_ (.A(_03511_),
    .B(_03058_),
    .X(_03059_));
 sky130_fd_sc_hd__or2_1 _12779_ (.A(\core_busio.mem_address[23] ),
    .B(net350),
    .X(_03060_));
 sky130_fd_sc_hd__a221o_2 _12780_ (.A1(\core_pipeline.csr_to_fetch_trap_vector[23] ),
    .A2(_03479_),
    .B1(_04385_),
    .B2(\core_pipeline.csr_to_fetch_mret_vector[23] ),
    .C1(net106),
    .X(_03061_));
 sky130_fd_sc_hd__a31o_1 _12781_ (.A1(_03514_),
    .A2(_03059_),
    .A3(_03060_),
    .B1(_03061_),
    .X(_03062_));
 sky130_fd_sc_hd__o211a_1 _12782_ (.A1(\core_pipeline.pipeline_fetch.pc[23] ),
    .A2(net103),
    .B1(_03062_),
    .C1(net636),
    .X(_01974_));
 sky130_fd_sc_hd__xor2_1 _12783_ (.A(\core_pipeline.pipeline_fetch.pc[24] ),
    .B(_03056_),
    .X(_03063_));
 sky130_fd_sc_hd__a21o_1 _12784_ (.A1(\core_pipeline.csr_to_fetch_trap_vector[24] ),
    .A2(_03479_),
    .B1(net106),
    .X(_03064_));
 sky130_fd_sc_hd__or2_1 _12785_ (.A(\core_pipeline.csr_to_fetch_mret_vector[24] ),
    .B(net445),
    .X(_03065_));
 sky130_fd_sc_hd__mux2_1 _12786_ (.A0(\core_busio.mem_address[24] ),
    .A1(_03063_),
    .S(net350),
    .X(_03066_));
 sky130_fd_sc_hd__o211a_1 _12787_ (.A1(_03512_),
    .A2(_03066_),
    .B1(_03065_),
    .C1(net403),
    .X(_03067_));
 sky130_fd_sc_hd__o221a_1 _12788_ (.A1(\core_pipeline.pipeline_fetch.pc[24] ),
    .A2(net103),
    .B1(_03064_),
    .B2(_03067_),
    .C1(net637),
    .X(_01975_));
 sky130_fd_sc_hd__and3_1 _12789_ (.A(\core_pipeline.pipeline_fetch.pc[25] ),
    .B(\core_pipeline.pipeline_fetch.pc[24] ),
    .C(_03056_),
    .X(_03068_));
 sky130_fd_sc_hd__a21oi_1 _12790_ (.A1(\core_pipeline.pipeline_fetch.pc[24] ),
    .A2(_03056_),
    .B1(\core_pipeline.pipeline_fetch.pc[25] ),
    .Y(_03069_));
 sky130_fd_sc_hd__o21ai_1 _12791_ (.A1(_03068_),
    .A2(_03069_),
    .B1(net350),
    .Y(_03070_));
 sky130_fd_sc_hd__or2_1 _12792_ (.A(\core_busio.mem_address[25] ),
    .B(net350),
    .X(_03071_));
 sky130_fd_sc_hd__a221o_2 _12793_ (.A1(\core_pipeline.csr_to_fetch_trap_vector[25] ),
    .A2(_03479_),
    .B1(_04385_),
    .B2(\core_pipeline.csr_to_fetch_mret_vector[25] ),
    .C1(net105),
    .X(_03072_));
 sky130_fd_sc_hd__a31o_1 _12794_ (.A1(_03514_),
    .A2(_03070_),
    .A3(_03071_),
    .B1(_03072_),
    .X(_03073_));
 sky130_fd_sc_hd__o211a_1 _12795_ (.A1(\core_pipeline.pipeline_fetch.pc[25] ),
    .A2(net103),
    .B1(_03073_),
    .C1(net636),
    .X(_01976_));
 sky130_fd_sc_hd__and2_2 _12796_ (.A(\core_pipeline.pipeline_fetch.pc[26] ),
    .B(_03068_),
    .X(_03074_));
 sky130_fd_sc_hd__or2_1 _12797_ (.A(\core_pipeline.pipeline_fetch.pc[26] ),
    .B(_03068_),
    .X(_03075_));
 sky130_fd_sc_hd__and2b_1 _12798_ (.A_N(_03074_),
    .B(_03075_),
    .X(_03076_));
 sky130_fd_sc_hd__or2_1 _12799_ (.A(_03511_),
    .B(_03076_),
    .X(_03077_));
 sky130_fd_sc_hd__or2_1 _12800_ (.A(\core_busio.mem_address[26] ),
    .B(net351),
    .X(_03078_));
 sky130_fd_sc_hd__a221o_2 _12801_ (.A1(\core_pipeline.csr_to_fetch_trap_vector[26] ),
    .A2(_03479_),
    .B1(_04385_),
    .B2(\core_pipeline.csr_to_fetch_mret_vector[26] ),
    .C1(net105),
    .X(_03079_));
 sky130_fd_sc_hd__a31o_1 _12802_ (.A1(_03514_),
    .A2(_03077_),
    .A3(_03078_),
    .B1(_03079_),
    .X(_03080_));
 sky130_fd_sc_hd__o211a_1 _12803_ (.A1(\core_pipeline.pipeline_fetch.pc[26] ),
    .A2(net103),
    .B1(_03080_),
    .C1(net636),
    .X(_01977_));
 sky130_fd_sc_hd__xor2_1 _12804_ (.A(\core_pipeline.pipeline_fetch.pc[27] ),
    .B(_03074_),
    .X(_03081_));
 sky130_fd_sc_hd__or2_1 _12805_ (.A(_03511_),
    .B(_03081_),
    .X(_03082_));
 sky130_fd_sc_hd__or2_1 _12806_ (.A(\core_busio.mem_address[27] ),
    .B(net351),
    .X(_03083_));
 sky130_fd_sc_hd__a221o_2 _12807_ (.A1(\core_pipeline.csr_to_fetch_trap_vector[27] ),
    .A2(_03479_),
    .B1(_04385_),
    .B2(\core_pipeline.csr_to_fetch_mret_vector[27] ),
    .C1(net105),
    .X(_03084_));
 sky130_fd_sc_hd__a31o_1 _12808_ (.A1(_03514_),
    .A2(_03082_),
    .A3(_03083_),
    .B1(_03084_),
    .X(_03085_));
 sky130_fd_sc_hd__o211a_1 _12809_ (.A1(\core_pipeline.pipeline_fetch.pc[27] ),
    .A2(net103),
    .B1(_03085_),
    .C1(net636),
    .X(_01978_));
 sky130_fd_sc_hd__and3_1 _12810_ (.A(\core_pipeline.pipeline_fetch.pc[28] ),
    .B(\core_pipeline.pipeline_fetch.pc[27] ),
    .C(_03074_),
    .X(_03086_));
 sky130_fd_sc_hd__a21oi_1 _12811_ (.A1(\core_pipeline.pipeline_fetch.pc[27] ),
    .A2(_03074_),
    .B1(\core_pipeline.pipeline_fetch.pc[28] ),
    .Y(_03087_));
 sky130_fd_sc_hd__nor2_1 _12812_ (.A(_03086_),
    .B(_03087_),
    .Y(_03088_));
 sky130_fd_sc_hd__or2_1 _12813_ (.A(_03511_),
    .B(_03088_),
    .X(_03089_));
 sky130_fd_sc_hd__or2_1 _12814_ (.A(\core_busio.mem_address[28] ),
    .B(net351),
    .X(_03090_));
 sky130_fd_sc_hd__a221o_1 _12815_ (.A1(\core_pipeline.csr_to_fetch_trap_vector[28] ),
    .A2(_03479_),
    .B1(_04385_),
    .B2(\core_pipeline.csr_to_fetch_mret_vector[28] ),
    .C1(net105),
    .X(_03091_));
 sky130_fd_sc_hd__a31o_1 _12816_ (.A1(_03514_),
    .A2(_03089_),
    .A3(_03090_),
    .B1(_03091_),
    .X(_03092_));
 sky130_fd_sc_hd__o211a_1 _12817_ (.A1(\core_pipeline.pipeline_fetch.pc[28] ),
    .A2(net104),
    .B1(_03092_),
    .C1(net638),
    .X(_01979_));
 sky130_fd_sc_hd__and2_2 _12818_ (.A(\core_pipeline.pipeline_fetch.pc[29] ),
    .B(_03086_),
    .X(_03093_));
 sky130_fd_sc_hd__nor2_1 _12819_ (.A(\core_pipeline.pipeline_fetch.pc[29] ),
    .B(_03086_),
    .Y(_03094_));
 sky130_fd_sc_hd__nor2_1 _12820_ (.A(_03093_),
    .B(_03094_),
    .Y(_03095_));
 sky130_fd_sc_hd__or2_1 _12821_ (.A(_03511_),
    .B(_03095_),
    .X(_03096_));
 sky130_fd_sc_hd__or2_1 _12822_ (.A(\core_busio.mem_address[29] ),
    .B(net351),
    .X(_03097_));
 sky130_fd_sc_hd__a221o_1 _12823_ (.A1(\core_pipeline.csr_to_fetch_trap_vector[29] ),
    .A2(_03479_),
    .B1(_04385_),
    .B2(\core_pipeline.csr_to_fetch_mret_vector[29] ),
    .C1(net105),
    .X(_03098_));
 sky130_fd_sc_hd__a31o_1 _12824_ (.A1(_03514_),
    .A2(_03096_),
    .A3(_03097_),
    .B1(_03098_),
    .X(_03099_));
 sky130_fd_sc_hd__o211a_1 _12825_ (.A1(\core_pipeline.pipeline_fetch.pc[29] ),
    .A2(net104),
    .B1(_03099_),
    .C1(net638),
    .X(_01980_));
 sky130_fd_sc_hd__nand2_1 _12826_ (.A(\core_pipeline.pipeline_fetch.pc[30] ),
    .B(_03093_),
    .Y(_03100_));
 sky130_fd_sc_hd__xor2_1 _12827_ (.A(\core_pipeline.pipeline_fetch.pc[30] ),
    .B(_03093_),
    .X(_03101_));
 sky130_fd_sc_hd__or2_1 _12828_ (.A(_03511_),
    .B(_03101_),
    .X(_03102_));
 sky130_fd_sc_hd__or2_1 _12829_ (.A(\core_busio.mem_address[30] ),
    .B(net351),
    .X(_03103_));
 sky130_fd_sc_hd__a221o_1 _12830_ (.A1(\core_pipeline.csr_to_fetch_trap_vector[30] ),
    .A2(_03479_),
    .B1(_04385_),
    .B2(\core_pipeline.csr_to_fetch_mret_vector[30] ),
    .C1(net105),
    .X(_03104_));
 sky130_fd_sc_hd__a31o_1 _12831_ (.A1(_03514_),
    .A2(_03102_),
    .A3(_03103_),
    .B1(_03104_),
    .X(_03105_));
 sky130_fd_sc_hd__o211a_1 _12832_ (.A1(\core_pipeline.pipeline_fetch.pc[30] ),
    .A2(net104),
    .B1(_03105_),
    .C1(net638),
    .X(_01981_));
 sky130_fd_sc_hd__xnor2_1 _12833_ (.A(\core_pipeline.pipeline_fetch.pc[31] ),
    .B(_03100_),
    .Y(_03106_));
 sky130_fd_sc_hd__or2_1 _12834_ (.A(\core_busio.mem_address[31] ),
    .B(net351),
    .X(_03107_));
 sky130_fd_sc_hd__o211a_1 _12835_ (.A1(_03511_),
    .A2(_03106_),
    .B1(_03107_),
    .C1(net445),
    .X(_03108_));
 sky130_fd_sc_hd__o21a_1 _12836_ (.A1(\core_pipeline.csr_to_fetch_mret_vector[31] ),
    .A2(_03479_),
    .B1(_03515_),
    .X(_03109_));
 sky130_fd_sc_hd__o221a_1 _12837_ (.A1(\core_pipeline.csr_to_fetch_trap_vector[31] ),
    .A2(net400),
    .B1(_03108_),
    .B2(_03109_),
    .C1(net104),
    .X(_03110_));
 sky130_fd_sc_hd__a211o_1 _12838_ (.A1(\core_pipeline.pipeline_fetch.pc[31] ),
    .A2(net105),
    .B1(_03110_),
    .C1(net35),
    .X(_01982_));
 sky130_fd_sc_hd__or3b_4 _12839_ (.A(\core_pipeline.memory_to_writeback_csr_address[0] ),
    .B(_03648_),
    .C_N(_05606_),
    .X(_03111_));
 sky130_fd_sc_hd__mux2_1 _12840_ (.A0(\core_pipeline.memory_to_writeback_alu_data[0] ),
    .A1(\core_pipeline.pipeline_csr.mtimecmp[0] ),
    .S(net166),
    .X(_01983_));
 sky130_fd_sc_hd__mux2_1 _12841_ (.A0(\core_pipeline.memory_to_writeback_alu_data[1] ),
    .A1(\core_pipeline.pipeline_csr.mtimecmp[1] ),
    .S(net166),
    .X(_01984_));
 sky130_fd_sc_hd__mux2_1 _12842_ (.A0(\core_pipeline.memory_to_writeback_alu_data[2] ),
    .A1(\core_pipeline.pipeline_csr.mtimecmp[2] ),
    .S(net166),
    .X(_01985_));
 sky130_fd_sc_hd__mux2_1 _12843_ (.A0(\core_pipeline.memory_to_writeback_alu_data[3] ),
    .A1(\core_pipeline.pipeline_csr.mtimecmp[3] ),
    .S(net166),
    .X(_01986_));
 sky130_fd_sc_hd__mux2_1 _12844_ (.A0(\core_pipeline.memory_to_writeback_alu_data[4] ),
    .A1(\core_pipeline.pipeline_csr.mtimecmp[4] ),
    .S(net166),
    .X(_01987_));
 sky130_fd_sc_hd__mux2_1 _12845_ (.A0(\core_pipeline.memory_to_writeback_alu_data[5] ),
    .A1(\core_pipeline.pipeline_csr.mtimecmp[5] ),
    .S(net166),
    .X(_01988_));
 sky130_fd_sc_hd__mux2_1 _12846_ (.A0(\core_pipeline.memory_to_writeback_alu_data[6] ),
    .A1(\core_pipeline.pipeline_csr.mtimecmp[6] ),
    .S(net166),
    .X(_01989_));
 sky130_fd_sc_hd__mux2_1 _12847_ (.A0(\core_pipeline.memory_to_writeback_alu_data[7] ),
    .A1(\core_pipeline.pipeline_csr.mtimecmp[7] ),
    .S(net166),
    .X(_01990_));
 sky130_fd_sc_hd__mux2_1 _12848_ (.A0(\core_pipeline.memory_to_writeback_alu_data[8] ),
    .A1(\core_pipeline.pipeline_csr.mtimecmp[8] ),
    .S(net165),
    .X(_01991_));
 sky130_fd_sc_hd__mux2_1 _12849_ (.A0(\core_pipeline.memory_to_writeback_alu_data[9] ),
    .A1(\core_pipeline.pipeline_csr.mtimecmp[9] ),
    .S(net165),
    .X(_01992_));
 sky130_fd_sc_hd__mux2_1 _12850_ (.A0(\core_pipeline.memory_to_writeback_alu_data[10] ),
    .A1(\core_pipeline.pipeline_csr.mtimecmp[10] ),
    .S(net165),
    .X(_01993_));
 sky130_fd_sc_hd__mux2_1 _12851_ (.A0(\core_pipeline.memory_to_writeback_alu_data[11] ),
    .A1(\core_pipeline.pipeline_csr.mtimecmp[11] ),
    .S(net165),
    .X(_01994_));
 sky130_fd_sc_hd__mux2_1 _12852_ (.A0(\core_pipeline.memory_to_writeback_alu_data[12] ),
    .A1(\core_pipeline.pipeline_csr.mtimecmp[12] ),
    .S(net165),
    .X(_01995_));
 sky130_fd_sc_hd__mux2_1 _12853_ (.A0(\core_pipeline.memory_to_writeback_alu_data[13] ),
    .A1(\core_pipeline.pipeline_csr.mtimecmp[13] ),
    .S(net165),
    .X(_01996_));
 sky130_fd_sc_hd__mux2_1 _12854_ (.A0(\core_pipeline.memory_to_writeback_alu_data[14] ),
    .A1(\core_pipeline.pipeline_csr.mtimecmp[14] ),
    .S(net165),
    .X(_01997_));
 sky130_fd_sc_hd__mux2_1 _12855_ (.A0(\core_pipeline.memory_to_writeback_alu_data[15] ),
    .A1(\core_pipeline.pipeline_csr.mtimecmp[15] ),
    .S(net165),
    .X(_01998_));
 sky130_fd_sc_hd__mux2_1 _12856_ (.A0(\core_pipeline.memory_to_writeback_alu_data[16] ),
    .A1(\core_pipeline.pipeline_csr.mtimecmp[16] ),
    .S(net165),
    .X(_01999_));
 sky130_fd_sc_hd__mux2_1 _12857_ (.A0(\core_pipeline.memory_to_writeback_alu_data[17] ),
    .A1(\core_pipeline.pipeline_csr.mtimecmp[17] ),
    .S(net165),
    .X(_02000_));
 sky130_fd_sc_hd__mux2_1 _12858_ (.A0(\core_pipeline.memory_to_writeback_alu_data[18] ),
    .A1(\core_pipeline.pipeline_csr.mtimecmp[18] ),
    .S(net166),
    .X(_02001_));
 sky130_fd_sc_hd__mux2_1 _12859_ (.A0(\core_pipeline.memory_to_writeback_alu_data[19] ),
    .A1(\core_pipeline.pipeline_csr.mtimecmp[19] ),
    .S(net165),
    .X(_02002_));
 sky130_fd_sc_hd__mux2_1 _12860_ (.A0(\core_pipeline.memory_to_writeback_alu_data[20] ),
    .A1(\core_pipeline.pipeline_csr.mtimecmp[20] ),
    .S(net165),
    .X(_02003_));
 sky130_fd_sc_hd__mux2_1 _12861_ (.A0(\core_pipeline.memory_to_writeback_alu_data[21] ),
    .A1(\core_pipeline.pipeline_csr.mtimecmp[21] ),
    .S(net166),
    .X(_02004_));
 sky130_fd_sc_hd__mux2_1 _12862_ (.A0(\core_pipeline.memory_to_writeback_alu_data[22] ),
    .A1(\core_pipeline.pipeline_csr.mtimecmp[22] ),
    .S(net165),
    .X(_02005_));
 sky130_fd_sc_hd__mux2_1 _12863_ (.A0(\core_pipeline.memory_to_writeback_alu_data[23] ),
    .A1(\core_pipeline.pipeline_csr.mtimecmp[23] ),
    .S(net165),
    .X(_02006_));
 sky130_fd_sc_hd__mux2_1 _12864_ (.A0(\core_pipeline.memory_to_writeback_alu_data[24] ),
    .A1(\core_pipeline.pipeline_csr.mtimecmp[24] ),
    .S(net165),
    .X(_02007_));
 sky130_fd_sc_hd__mux2_1 _12865_ (.A0(\core_pipeline.memory_to_writeback_alu_data[25] ),
    .A1(\core_pipeline.pipeline_csr.mtimecmp[25] ),
    .S(net165),
    .X(_02008_));
 sky130_fd_sc_hd__mux2_1 _12866_ (.A0(\core_pipeline.memory_to_writeback_alu_data[26] ),
    .A1(\core_pipeline.pipeline_csr.mtimecmp[26] ),
    .S(net165),
    .X(_02009_));
 sky130_fd_sc_hd__mux2_1 _12867_ (.A0(\core_pipeline.memory_to_writeback_alu_data[27] ),
    .A1(\core_pipeline.pipeline_csr.mtimecmp[27] ),
    .S(net166),
    .X(_02010_));
 sky130_fd_sc_hd__mux2_1 _12868_ (.A0(\core_pipeline.memory_to_writeback_alu_data[28] ),
    .A1(\core_pipeline.pipeline_csr.mtimecmp[28] ),
    .S(net166),
    .X(_02011_));
 sky130_fd_sc_hd__mux2_1 _12869_ (.A0(\core_pipeline.memory_to_writeback_alu_data[29] ),
    .A1(\core_pipeline.pipeline_csr.mtimecmp[29] ),
    .S(net166),
    .X(_02012_));
 sky130_fd_sc_hd__mux2_1 _12870_ (.A0(\core_pipeline.memory_to_writeback_alu_data[30] ),
    .A1(\core_pipeline.pipeline_csr.mtimecmp[30] ),
    .S(net166),
    .X(_02013_));
 sky130_fd_sc_hd__mux2_1 _12871_ (.A0(\core_pipeline.memory_to_writeback_alu_data[31] ),
    .A1(\core_pipeline.pipeline_csr.mtimecmp[31] ),
    .S(net166),
    .X(_02014_));
 sky130_fd_sc_hd__mux2_1 _12872_ (.A0(\core_pipeline.decode_to_execute_pc[2] ),
    .A1(\core_pipeline.fetch_to_decode_pc[2] ),
    .S(net147),
    .X(_02015_));
 sky130_fd_sc_hd__mux2_1 _12873_ (.A0(\core_pipeline.decode_to_execute_pc[3] ),
    .A1(\core_pipeline.fetch_to_decode_pc[3] ),
    .S(net157),
    .X(_02016_));
 sky130_fd_sc_hd__mux2_1 _12874_ (.A0(\core_pipeline.decode_to_execute_pc[4] ),
    .A1(\core_pipeline.fetch_to_decode_pc[4] ),
    .S(net152),
    .X(_02017_));
 sky130_fd_sc_hd__mux2_1 _12875_ (.A0(\core_pipeline.decode_to_execute_pc[5] ),
    .A1(\core_pipeline.fetch_to_decode_pc[5] ),
    .S(net152),
    .X(_02018_));
 sky130_fd_sc_hd__mux2_1 _12876_ (.A0(\core_pipeline.decode_to_execute_pc[6] ),
    .A1(\core_pipeline.fetch_to_decode_pc[6] ),
    .S(net152),
    .X(_02019_));
 sky130_fd_sc_hd__mux2_1 _12877_ (.A0(\core_pipeline.decode_to_execute_pc[7] ),
    .A1(\core_pipeline.fetch_to_decode_pc[7] ),
    .S(net158),
    .X(_02020_));
 sky130_fd_sc_hd__mux2_1 _12878_ (.A0(\core_pipeline.decode_to_execute_pc[8] ),
    .A1(\core_pipeline.fetch_to_decode_pc[8] ),
    .S(net150),
    .X(_02021_));
 sky130_fd_sc_hd__mux2_1 _12879_ (.A0(\core_pipeline.decode_to_execute_pc[9] ),
    .A1(\core_pipeline.fetch_to_decode_pc[9] ),
    .S(net153),
    .X(_02022_));
 sky130_fd_sc_hd__mux2_1 _12880_ (.A0(\core_pipeline.decode_to_execute_pc[10] ),
    .A1(\core_pipeline.fetch_to_decode_pc[10] ),
    .S(net154),
    .X(_02023_));
 sky130_fd_sc_hd__mux2_1 _12881_ (.A0(\core_pipeline.decode_to_execute_pc[11] ),
    .A1(\core_pipeline.fetch_to_decode_pc[11] ),
    .S(net156),
    .X(_02024_));
 sky130_fd_sc_hd__mux2_1 _12882_ (.A0(\core_pipeline.decode_to_execute_pc[12] ),
    .A1(\core_pipeline.fetch_to_decode_pc[12] ),
    .S(net156),
    .X(_02025_));
 sky130_fd_sc_hd__mux2_1 _12883_ (.A0(\core_pipeline.decode_to_execute_pc[13] ),
    .A1(\core_pipeline.fetch_to_decode_pc[13] ),
    .S(net153),
    .X(_02026_));
 sky130_fd_sc_hd__mux2_1 _12884_ (.A0(\core_pipeline.decode_to_execute_pc[14] ),
    .A1(\core_pipeline.fetch_to_decode_pc[14] ),
    .S(net154),
    .X(_02027_));
 sky130_fd_sc_hd__mux2_1 _12885_ (.A0(\core_pipeline.decode_to_execute_pc[15] ),
    .A1(\core_pipeline.fetch_to_decode_pc[15] ),
    .S(net156),
    .X(_02028_));
 sky130_fd_sc_hd__mux2_1 _12886_ (.A0(\core_pipeline.decode_to_execute_pc[16] ),
    .A1(\core_pipeline.fetch_to_decode_pc[16] ),
    .S(net153),
    .X(_02029_));
 sky130_fd_sc_hd__mux2_1 _12887_ (.A0(\core_pipeline.decode_to_execute_pc[17] ),
    .A1(\core_pipeline.fetch_to_decode_pc[17] ),
    .S(net161),
    .X(_02030_));
 sky130_fd_sc_hd__mux2_1 _12888_ (.A0(\core_pipeline.decode_to_execute_pc[18] ),
    .A1(\core_pipeline.fetch_to_decode_pc[18] ),
    .S(net161),
    .X(_02031_));
 sky130_fd_sc_hd__mux2_1 _12889_ (.A0(\core_pipeline.decode_to_execute_pc[19] ),
    .A1(\core_pipeline.fetch_to_decode_pc[19] ),
    .S(net161),
    .X(_02032_));
 sky130_fd_sc_hd__mux2_1 _12890_ (.A0(\core_pipeline.decode_to_execute_pc[20] ),
    .A1(\core_pipeline.fetch_to_decode_pc[20] ),
    .S(net160),
    .X(_02033_));
 sky130_fd_sc_hd__mux2_1 _12891_ (.A0(\core_pipeline.decode_to_execute_pc[21] ),
    .A1(\core_pipeline.fetch_to_decode_pc[21] ),
    .S(net157),
    .X(_02034_));
 sky130_fd_sc_hd__mux2_1 _12892_ (.A0(\core_pipeline.decode_to_execute_pc[22] ),
    .A1(\core_pipeline.fetch_to_decode_pc[22] ),
    .S(net160),
    .X(_02035_));
 sky130_fd_sc_hd__mux2_1 _12893_ (.A0(\core_pipeline.decode_to_execute_pc[23] ),
    .A1(\core_pipeline.fetch_to_decode_pc[23] ),
    .S(net155),
    .X(_02036_));
 sky130_fd_sc_hd__mux2_1 _12894_ (.A0(\core_pipeline.decode_to_execute_pc[24] ),
    .A1(\core_pipeline.fetch_to_decode_pc[24] ),
    .S(net155),
    .X(_02037_));
 sky130_fd_sc_hd__mux2_1 _12895_ (.A0(\core_pipeline.decode_to_execute_pc[25] ),
    .A1(\core_pipeline.fetch_to_decode_pc[25] ),
    .S(net155),
    .X(_02038_));
 sky130_fd_sc_hd__mux2_1 _12896_ (.A0(\core_pipeline.decode_to_execute_pc[26] ),
    .A1(\core_pipeline.fetch_to_decode_pc[26] ),
    .S(net160),
    .X(_02039_));
 sky130_fd_sc_hd__mux2_1 _12897_ (.A0(\core_pipeline.decode_to_execute_pc[27] ),
    .A1(\core_pipeline.fetch_to_decode_pc[27] ),
    .S(net158),
    .X(_02040_));
 sky130_fd_sc_hd__mux2_1 _12898_ (.A0(\core_pipeline.decode_to_execute_pc[28] ),
    .A1(\core_pipeline.fetch_to_decode_pc[28] ),
    .S(net157),
    .X(_02041_));
 sky130_fd_sc_hd__mux2_1 _12899_ (.A0(\core_pipeline.decode_to_execute_pc[29] ),
    .A1(\core_pipeline.fetch_to_decode_pc[29] ),
    .S(net151),
    .X(_02042_));
 sky130_fd_sc_hd__mux2_1 _12900_ (.A0(\core_pipeline.decode_to_execute_pc[30] ),
    .A1(\core_pipeline.fetch_to_decode_pc[30] ),
    .S(net152),
    .X(_02043_));
 sky130_fd_sc_hd__mux2_1 _12901_ (.A0(\core_pipeline.decode_to_execute_pc[31] ),
    .A1(\core_pipeline.fetch_to_decode_pc[31] ),
    .S(net157),
    .X(_02044_));
 sky130_fd_sc_hd__mux2_1 _12902_ (.A0(\core_pipeline.decode_to_execute_next_pc[0] ),
    .A1(\core_pipeline.fetch_to_decode_next_pc[0] ),
    .S(net149),
    .X(_02045_));
 sky130_fd_sc_hd__mux2_1 _12903_ (.A0(\core_pipeline.decode_to_execute_next_pc[1] ),
    .A1(\core_pipeline.fetch_to_decode_next_pc[1] ),
    .S(net147),
    .X(_02046_));
 sky130_fd_sc_hd__mux2_1 _12904_ (.A0(\core_pipeline.decode_to_execute_next_pc[2] ),
    .A1(\core_pipeline.fetch_to_decode_next_pc[2] ),
    .S(net147),
    .X(_02047_));
 sky130_fd_sc_hd__mux2_1 _12905_ (.A0(\core_pipeline.decode_to_execute_next_pc[3] ),
    .A1(\core_pipeline.fetch_to_decode_next_pc[3] ),
    .S(net157),
    .X(_02048_));
 sky130_fd_sc_hd__mux2_1 _12906_ (.A0(\core_pipeline.decode_to_execute_next_pc[4] ),
    .A1(\core_pipeline.fetch_to_decode_next_pc[4] ),
    .S(net149),
    .X(_02049_));
 sky130_fd_sc_hd__mux2_1 _12907_ (.A0(\core_pipeline.decode_to_execute_next_pc[5] ),
    .A1(\core_pipeline.fetch_to_decode_next_pc[5] ),
    .S(net157),
    .X(_02050_));
 sky130_fd_sc_hd__mux2_1 _12908_ (.A0(\core_pipeline.decode_to_execute_next_pc[6] ),
    .A1(\core_pipeline.fetch_to_decode_next_pc[6] ),
    .S(net151),
    .X(_02051_));
 sky130_fd_sc_hd__mux2_1 _12909_ (.A0(\core_pipeline.decode_to_execute_next_pc[7] ),
    .A1(\core_pipeline.fetch_to_decode_next_pc[7] ),
    .S(net158),
    .X(_02052_));
 sky130_fd_sc_hd__mux2_1 _12910_ (.A0(\core_pipeline.decode_to_execute_next_pc[8] ),
    .A1(\core_pipeline.fetch_to_decode_next_pc[8] ),
    .S(net151),
    .X(_02053_));
 sky130_fd_sc_hd__mux2_1 _12911_ (.A0(\core_pipeline.decode_to_execute_next_pc[9] ),
    .A1(\core_pipeline.fetch_to_decode_next_pc[9] ),
    .S(net154),
    .X(_02054_));
 sky130_fd_sc_hd__mux2_1 _12912_ (.A0(\core_pipeline.decode_to_execute_next_pc[10] ),
    .A1(\core_pipeline.fetch_to_decode_next_pc[10] ),
    .S(net154),
    .X(_02055_));
 sky130_fd_sc_hd__mux2_1 _12913_ (.A0(\core_pipeline.decode_to_execute_next_pc[11] ),
    .A1(\core_pipeline.fetch_to_decode_next_pc[11] ),
    .S(net154),
    .X(_02056_));
 sky130_fd_sc_hd__mux2_1 _12914_ (.A0(\core_pipeline.decode_to_execute_next_pc[12] ),
    .A1(\core_pipeline.fetch_to_decode_next_pc[12] ),
    .S(net153),
    .X(_02057_));
 sky130_fd_sc_hd__mux2_1 _12915_ (.A0(\core_pipeline.decode_to_execute_next_pc[13] ),
    .A1(\core_pipeline.fetch_to_decode_next_pc[13] ),
    .S(net154),
    .X(_02058_));
 sky130_fd_sc_hd__mux2_1 _12916_ (.A0(\core_pipeline.decode_to_execute_next_pc[14] ),
    .A1(\core_pipeline.fetch_to_decode_next_pc[14] ),
    .S(net161),
    .X(_02059_));
 sky130_fd_sc_hd__mux2_1 _12917_ (.A0(\core_pipeline.decode_to_execute_next_pc[15] ),
    .A1(\core_pipeline.fetch_to_decode_next_pc[15] ),
    .S(net153),
    .X(_02060_));
 sky130_fd_sc_hd__mux2_1 _12918_ (.A0(\core_pipeline.decode_to_execute_next_pc[16] ),
    .A1(\core_pipeline.fetch_to_decode_next_pc[16] ),
    .S(net154),
    .X(_02061_));
 sky130_fd_sc_hd__mux2_1 _12919_ (.A0(\core_pipeline.decode_to_execute_next_pc[17] ),
    .A1(\core_pipeline.fetch_to_decode_next_pc[17] ),
    .S(net161),
    .X(_02062_));
 sky130_fd_sc_hd__mux2_1 _12920_ (.A0(\core_pipeline.decode_to_execute_next_pc[18] ),
    .A1(\core_pipeline.fetch_to_decode_next_pc[18] ),
    .S(net161),
    .X(_02063_));
 sky130_fd_sc_hd__mux2_1 _12921_ (.A0(\core_pipeline.decode_to_execute_next_pc[19] ),
    .A1(\core_pipeline.fetch_to_decode_next_pc[19] ),
    .S(net161),
    .X(_02064_));
 sky130_fd_sc_hd__mux2_1 _12922_ (.A0(\core_pipeline.decode_to_execute_next_pc[20] ),
    .A1(\core_pipeline.fetch_to_decode_next_pc[20] ),
    .S(net160),
    .X(_02065_));
 sky130_fd_sc_hd__mux2_1 _12923_ (.A0(\core_pipeline.decode_to_execute_next_pc[21] ),
    .A1(\core_pipeline.fetch_to_decode_next_pc[21] ),
    .S(net160),
    .X(_02066_));
 sky130_fd_sc_hd__mux2_1 _12924_ (.A0(\core_pipeline.decode_to_execute_next_pc[22] ),
    .A1(\core_pipeline.fetch_to_decode_next_pc[22] ),
    .S(net160),
    .X(_02067_));
 sky130_fd_sc_hd__mux2_1 _12925_ (.A0(\core_pipeline.decode_to_execute_next_pc[23] ),
    .A1(\core_pipeline.fetch_to_decode_next_pc[23] ),
    .S(net160),
    .X(_02068_));
 sky130_fd_sc_hd__mux2_1 _12926_ (.A0(\core_pipeline.decode_to_execute_next_pc[24] ),
    .A1(\core_pipeline.fetch_to_decode_next_pc[24] ),
    .S(net155),
    .X(_02069_));
 sky130_fd_sc_hd__mux2_1 _12927_ (.A0(\core_pipeline.decode_to_execute_next_pc[25] ),
    .A1(\core_pipeline.fetch_to_decode_next_pc[25] ),
    .S(net155),
    .X(_02070_));
 sky130_fd_sc_hd__mux2_1 _12928_ (.A0(\core_pipeline.decode_to_execute_next_pc[26] ),
    .A1(\core_pipeline.fetch_to_decode_next_pc[26] ),
    .S(net161),
    .X(_02071_));
 sky130_fd_sc_hd__mux2_1 _12929_ (.A0(\core_pipeline.decode_to_execute_next_pc[27] ),
    .A1(\core_pipeline.fetch_to_decode_next_pc[27] ),
    .S(net160),
    .X(_02072_));
 sky130_fd_sc_hd__mux2_1 _12930_ (.A0(\core_pipeline.decode_to_execute_next_pc[28] ),
    .A1(\core_pipeline.fetch_to_decode_next_pc[28] ),
    .S(net158),
    .X(_02073_));
 sky130_fd_sc_hd__mux2_1 _12931_ (.A0(\core_pipeline.decode_to_execute_next_pc[29] ),
    .A1(\core_pipeline.fetch_to_decode_next_pc[29] ),
    .S(net158),
    .X(_02074_));
 sky130_fd_sc_hd__mux2_1 _12932_ (.A0(\core_pipeline.decode_to_execute_next_pc[30] ),
    .A1(\core_pipeline.fetch_to_decode_next_pc[30] ),
    .S(net157),
    .X(_02075_));
 sky130_fd_sc_hd__mux2_1 _12933_ (.A0(\core_pipeline.decode_to_execute_next_pc[31] ),
    .A1(\core_pipeline.fetch_to_decode_next_pc[31] ),
    .S(net158),
    .X(_02076_));
 sky130_fd_sc_hd__nand2_1 _12934_ (.A(\core_pipeline.execute_to_memory_valid ),
    .B(\core_pipeline.execute_to_memory_bypass_memory ),
    .Y(_03112_));
 sky130_fd_sc_hd__o21ai_1 _12935_ (.A1(net602),
    .A2(_04630_),
    .B1(_03112_),
    .Y(_03113_));
 sky130_fd_sc_hd__o211a_2 _12936_ (.A1(_03497_),
    .A2(_03112_),
    .B1(_03113_),
    .C1(_03499_),
    .X(_03114_));
 sky130_fd_sc_hd__mux2_1 _12937_ (.A0(_05840_),
    .A1(\core_pipeline.execute_to_memory_csr_data[0] ),
    .S(net499),
    .X(_03115_));
 sky130_fd_sc_hd__a22o_1 _12938_ (.A1(net573),
    .A2(_04468_),
    .B1(_04936_),
    .B2(net579),
    .X(_03116_));
 sky130_fd_sc_hd__o22ai_1 _12939_ (.A1(net626),
    .A2(_03913_),
    .B1(_03914_),
    .B2(net594),
    .Y(_03117_));
 sky130_fd_sc_hd__o2bb2a_1 _12940_ (.A1_N(net594),
    .A2_N(_03914_),
    .B1(_04468_),
    .B2(net575),
    .X(_03118_));
 sky130_fd_sc_hd__o221ai_2 _12941_ (.A1(net568),
    .A2(_03912_),
    .B1(_04936_),
    .B2(net579),
    .C1(_03118_),
    .Y(_03119_));
 sky130_fd_sc_hd__a221o_1 _12942_ (.A1(net568),
    .A2(_03912_),
    .B1(_03913_),
    .B2(net626),
    .C1(_03119_),
    .X(_03120_));
 sky130_fd_sc_hd__or3_2 _12943_ (.A(_03116_),
    .B(_03117_),
    .C(_03120_),
    .X(_03121_));
 sky130_fd_sc_hd__nor2_4 _12944_ (.A(net239),
    .B(_03121_),
    .Y(_03122_));
 sky130_fd_sc_hd__a22o_1 _12945_ (.A1(net240),
    .A2(_03115_),
    .B1(net117),
    .B2(_03922_),
    .X(_03123_));
 sky130_fd_sc_hd__nor2_4 _12946_ (.A(net132),
    .B(_04631_),
    .Y(_03124_));
 sky130_fd_sc_hd__a22o_1 _12947_ (.A1(\core_pipeline.decode_to_execute_rs1_bypass[0] ),
    .A2(net122),
    .B1(_03123_),
    .B2(net115),
    .X(_02077_));
 sky130_fd_sc_hd__mux2_2 _12948_ (.A0(_05845_),
    .A1(\core_pipeline.execute_to_memory_csr_data[1] ),
    .S(net499),
    .X(_03125_));
 sky130_fd_sc_hd__a22o_1 _12949_ (.A1(_03925_),
    .A2(net118),
    .B1(_03125_),
    .B2(net239),
    .X(_03126_));
 sky130_fd_sc_hd__a22o_1 _12950_ (.A1(\core_pipeline.decode_to_execute_rs1_bypass[1] ),
    .A2(net125),
    .B1(net116),
    .B2(_03126_),
    .X(_02078_));
 sky130_fd_sc_hd__mux2_2 _12951_ (.A0(_05849_),
    .A1(\core_pipeline.execute_to_memory_csr_data[2] ),
    .S(net499),
    .X(_03127_));
 sky130_fd_sc_hd__a22o_1 _12952_ (.A1(_03928_),
    .A2(net118),
    .B1(_03127_),
    .B2(net239),
    .X(_03128_));
 sky130_fd_sc_hd__a22o_1 _12953_ (.A1(\core_pipeline.decode_to_execute_rs1_bypass[2] ),
    .A2(net130),
    .B1(net116),
    .B2(_03128_),
    .X(_02079_));
 sky130_fd_sc_hd__mux2_2 _12954_ (.A0(_05853_),
    .A1(\core_pipeline.execute_to_memory_csr_data[3] ),
    .S(net499),
    .X(_03129_));
 sky130_fd_sc_hd__a22o_1 _12955_ (.A1(_03931_),
    .A2(net117),
    .B1(_03129_),
    .B2(net240),
    .X(_03130_));
 sky130_fd_sc_hd__a22o_1 _12956_ (.A1(\core_pipeline.decode_to_execute_rs1_bypass[3] ),
    .A2(net121),
    .B1(net115),
    .B2(_03130_),
    .X(_02080_));
 sky130_fd_sc_hd__mux2_2 _12957_ (.A0(_05857_),
    .A1(\core_pipeline.execute_to_memory_csr_data[4] ),
    .S(net499),
    .X(_03131_));
 sky130_fd_sc_hd__a22o_1 _12958_ (.A1(_03934_),
    .A2(net117),
    .B1(_03131_),
    .B2(net240),
    .X(_03132_));
 sky130_fd_sc_hd__a22o_1 _12959_ (.A1(\core_pipeline.decode_to_execute_rs1_bypass[4] ),
    .A2(net121),
    .B1(net115),
    .B2(_03132_),
    .X(_02081_));
 sky130_fd_sc_hd__mux2_2 _12960_ (.A0(_05861_),
    .A1(\core_pipeline.execute_to_memory_csr_data[5] ),
    .S(net499),
    .X(_03133_));
 sky130_fd_sc_hd__a22o_1 _12961_ (.A1(net339),
    .A2(net118),
    .B1(_03133_),
    .B2(net239),
    .X(_03134_));
 sky130_fd_sc_hd__a22o_1 _12962_ (.A1(\core_pipeline.decode_to_execute_rs1_bypass[5] ),
    .A2(net124),
    .B1(net116),
    .B2(_03134_),
    .X(_02082_));
 sky130_fd_sc_hd__mux2_4 _12963_ (.A0(_05865_),
    .A1(\core_pipeline.execute_to_memory_csr_data[6] ),
    .S(net499),
    .X(_03135_));
 sky130_fd_sc_hd__a22o_1 _12964_ (.A1(_03940_),
    .A2(net117),
    .B1(_03135_),
    .B2(net239),
    .X(_03136_));
 sky130_fd_sc_hd__a22o_1 _12965_ (.A1(\core_pipeline.decode_to_execute_rs1_bypass[6] ),
    .A2(net125),
    .B1(net115),
    .B2(_03136_),
    .X(_02083_));
 sky130_fd_sc_hd__mux2_2 _12966_ (.A0(_05869_),
    .A1(\core_pipeline.execute_to_memory_csr_data[7] ),
    .S(net499),
    .X(_03137_));
 sky130_fd_sc_hd__a22o_1 _12967_ (.A1(net334),
    .A2(net117),
    .B1(_03137_),
    .B2(net240),
    .X(_03138_));
 sky130_fd_sc_hd__a22o_1 _12968_ (.A1(\core_pipeline.decode_to_execute_rs1_bypass[7] ),
    .A2(net122),
    .B1(net115),
    .B2(_03138_),
    .X(_02084_));
 sky130_fd_sc_hd__mux2_4 _12969_ (.A0(_05873_),
    .A1(\core_pipeline.execute_to_memory_csr_data[8] ),
    .S(net498),
    .X(_03139_));
 sky130_fd_sc_hd__a22o_1 _12970_ (.A1(_03946_),
    .A2(net117),
    .B1(_03139_),
    .B2(net240),
    .X(_03140_));
 sky130_fd_sc_hd__a22o_1 _12971_ (.A1(\core_pipeline.decode_to_execute_rs1_bypass[8] ),
    .A2(net124),
    .B1(net115),
    .B2(_03140_),
    .X(_02085_));
 sky130_fd_sc_hd__mux2_8 _12972_ (.A0(_05877_),
    .A1(\core_pipeline.execute_to_memory_csr_data[9] ),
    .S(net498),
    .X(_03141_));
 sky130_fd_sc_hd__a22o_1 _12973_ (.A1(net330),
    .A2(net117),
    .B1(_03141_),
    .B2(net240),
    .X(_03142_));
 sky130_fd_sc_hd__a22o_1 _12974_ (.A1(\core_pipeline.decode_to_execute_rs1_bypass[9] ),
    .A2(net122),
    .B1(net115),
    .B2(_03142_),
    .X(_02086_));
 sky130_fd_sc_hd__mux2_4 _12975_ (.A0(_05881_),
    .A1(\core_pipeline.execute_to_memory_csr_data[10] ),
    .S(net498),
    .X(_03143_));
 sky130_fd_sc_hd__a22o_1 _12976_ (.A1(net328),
    .A2(net117),
    .B1(_03143_),
    .B2(net240),
    .X(_03144_));
 sky130_fd_sc_hd__a22o_1 _12977_ (.A1(\core_pipeline.decode_to_execute_rs1_bypass[10] ),
    .A2(net122),
    .B1(net115),
    .B2(_03144_),
    .X(_02087_));
 sky130_fd_sc_hd__mux2_4 _12978_ (.A0(_05885_),
    .A1(\core_pipeline.execute_to_memory_csr_data[11] ),
    .S(net498),
    .X(_03145_));
 sky130_fd_sc_hd__a22o_1 _12979_ (.A1(net326),
    .A2(net117),
    .B1(_03145_),
    .B2(net240),
    .X(_03146_));
 sky130_fd_sc_hd__a22o_1 _12980_ (.A1(\core_pipeline.decode_to_execute_rs1_bypass[11] ),
    .A2(net121),
    .B1(net115),
    .B2(_03146_),
    .X(_02088_));
 sky130_fd_sc_hd__mux2_8 _12981_ (.A0(_05889_),
    .A1(\core_pipeline.execute_to_memory_csr_data[12] ),
    .S(net498),
    .X(_03147_));
 sky130_fd_sc_hd__a22o_1 _12982_ (.A1(_03958_),
    .A2(net117),
    .B1(_03147_),
    .B2(net240),
    .X(_03148_));
 sky130_fd_sc_hd__a22o_1 _12983_ (.A1(\core_pipeline.decode_to_execute_rs1_bypass[12] ),
    .A2(net122),
    .B1(net115),
    .B2(_03148_),
    .X(_02089_));
 sky130_fd_sc_hd__mux2_8 _12984_ (.A0(_05893_),
    .A1(\core_pipeline.execute_to_memory_csr_data[13] ),
    .S(net498),
    .X(_03149_));
 sky130_fd_sc_hd__a22o_1 _12985_ (.A1(net322),
    .A2(net117),
    .B1(_03149_),
    .B2(net240),
    .X(_03150_));
 sky130_fd_sc_hd__a22o_1 _12986_ (.A1(\core_pipeline.decode_to_execute_rs1_bypass[13] ),
    .A2(net123),
    .B1(net115),
    .B2(_03150_),
    .X(_02090_));
 sky130_fd_sc_hd__mux2_8 _12987_ (.A0(_05897_),
    .A1(\core_pipeline.execute_to_memory_csr_data[14] ),
    .S(net498),
    .X(_03151_));
 sky130_fd_sc_hd__a22o_1 _12988_ (.A1(net320),
    .A2(net117),
    .B1(_03151_),
    .B2(net240),
    .X(_03152_));
 sky130_fd_sc_hd__a22o_1 _12989_ (.A1(\core_pipeline.decode_to_execute_rs1_bypass[14] ),
    .A2(net123),
    .B1(net115),
    .B2(_03152_),
    .X(_02091_));
 sky130_fd_sc_hd__mux2_4 _12990_ (.A0(_05901_),
    .A1(\core_pipeline.execute_to_memory_csr_data[15] ),
    .S(net498),
    .X(_03153_));
 sky130_fd_sc_hd__a22o_1 _12991_ (.A1(net318),
    .A2(net117),
    .B1(_03153_),
    .B2(net240),
    .X(_03154_));
 sky130_fd_sc_hd__a22o_1 _12992_ (.A1(\core_pipeline.decode_to_execute_rs1_bypass[15] ),
    .A2(net122),
    .B1(net115),
    .B2(_03154_),
    .X(_02092_));
 sky130_fd_sc_hd__mux2_8 _12993_ (.A0(_05905_),
    .A1(\core_pipeline.execute_to_memory_csr_data[16] ),
    .S(net498),
    .X(_03155_));
 sky130_fd_sc_hd__a22o_1 _12994_ (.A1(_03970_),
    .A2(net117),
    .B1(_03155_),
    .B2(net240),
    .X(_03156_));
 sky130_fd_sc_hd__a22o_1 _12995_ (.A1(\core_pipeline.decode_to_execute_rs1_bypass[16] ),
    .A2(net124),
    .B1(net115),
    .B2(_03156_),
    .X(_02093_));
 sky130_fd_sc_hd__mux2_8 _12996_ (.A0(_05909_),
    .A1(\core_pipeline.execute_to_memory_csr_data[17] ),
    .S(net499),
    .X(_03157_));
 sky130_fd_sc_hd__a22o_1 _12997_ (.A1(net314),
    .A2(net118),
    .B1(_03157_),
    .B2(net239),
    .X(_03158_));
 sky130_fd_sc_hd__a22o_1 _12998_ (.A1(\core_pipeline.decode_to_execute_rs1_bypass[17] ),
    .A2(net131),
    .B1(net116),
    .B2(_03158_),
    .X(_02094_));
 sky130_fd_sc_hd__mux2_4 _12999_ (.A0(_05913_),
    .A1(\core_pipeline.execute_to_memory_csr_data[18] ),
    .S(net498),
    .X(_03159_));
 sky130_fd_sc_hd__a22o_1 _13000_ (.A1(_03976_),
    .A2(net118),
    .B1(_03159_),
    .B2(net239),
    .X(_03160_));
 sky130_fd_sc_hd__a22o_1 _13001_ (.A1(\core_pipeline.decode_to_execute_rs1_bypass[18] ),
    .A2(net133),
    .B1(net116),
    .B2(_03160_),
    .X(_02095_));
 sky130_fd_sc_hd__mux2_8 _13002_ (.A0(_05917_),
    .A1(\core_pipeline.execute_to_memory_csr_data[19] ),
    .S(net498),
    .X(_03161_));
 sky130_fd_sc_hd__a22o_1 _13003_ (.A1(_03979_),
    .A2(net118),
    .B1(_03161_),
    .B2(net239),
    .X(_03162_));
 sky130_fd_sc_hd__a22o_1 _13004_ (.A1(\core_pipeline.decode_to_execute_rs1_bypass[19] ),
    .A2(net131),
    .B1(net116),
    .B2(_03162_),
    .X(_02096_));
 sky130_fd_sc_hd__mux2_4 _13005_ (.A0(_05921_),
    .A1(\core_pipeline.execute_to_memory_csr_data[20] ),
    .S(\core_pipeline.execute_to_memory_write_select[0] ),
    .X(_03163_));
 sky130_fd_sc_hd__a22o_1 _13006_ (.A1(net307),
    .A2(net118),
    .B1(_03163_),
    .B2(net239),
    .X(_03164_));
 sky130_fd_sc_hd__a22o_1 _13007_ (.A1(\core_pipeline.decode_to_execute_rs1_bypass[20] ),
    .A2(net131),
    .B1(net116),
    .B2(_03164_),
    .X(_02097_));
 sky130_fd_sc_hd__mux2_4 _13008_ (.A0(_05925_),
    .A1(\core_pipeline.execute_to_memory_csr_data[21] ),
    .S(net499),
    .X(_03165_));
 sky130_fd_sc_hd__a22o_1 _13009_ (.A1(_03985_),
    .A2(net118),
    .B1(_03165_),
    .B2(net239),
    .X(_03166_));
 sky130_fd_sc_hd__a22o_1 _13010_ (.A1(\core_pipeline.decode_to_execute_rs1_bypass[21] ),
    .A2(net133),
    .B1(net116),
    .B2(_03166_),
    .X(_02098_));
 sky130_fd_sc_hd__mux2_4 _13011_ (.A0(_05929_),
    .A1(\core_pipeline.execute_to_memory_csr_data[22] ),
    .S(net498),
    .X(_03167_));
 sky130_fd_sc_hd__a22o_1 _13012_ (.A1(_03988_),
    .A2(net118),
    .B1(_03167_),
    .B2(net239),
    .X(_03168_));
 sky130_fd_sc_hd__a22o_1 _13013_ (.A1(\core_pipeline.decode_to_execute_rs1_bypass[22] ),
    .A2(net130),
    .B1(net116),
    .B2(_03168_),
    .X(_02099_));
 sky130_fd_sc_hd__mux2_4 _13014_ (.A0(_05933_),
    .A1(\core_pipeline.execute_to_memory_csr_data[23] ),
    .S(net499),
    .X(_03169_));
 sky130_fd_sc_hd__a22o_1 _13015_ (.A1(net300),
    .A2(net118),
    .B1(_03169_),
    .B2(net239),
    .X(_03170_));
 sky130_fd_sc_hd__a22o_1 _13016_ (.A1(\core_pipeline.decode_to_execute_rs1_bypass[23] ),
    .A2(net124),
    .B1(net116),
    .B2(_03170_),
    .X(_02100_));
 sky130_fd_sc_hd__mux2_8 _13017_ (.A0(_05937_),
    .A1(\core_pipeline.execute_to_memory_csr_data[24] ),
    .S(net498),
    .X(_03171_));
 sky130_fd_sc_hd__a22o_1 _13018_ (.A1(net298),
    .A2(net117),
    .B1(_03171_),
    .B2(net240),
    .X(_03172_));
 sky130_fd_sc_hd__a22o_1 _13019_ (.A1(\core_pipeline.decode_to_execute_rs1_bypass[24] ),
    .A2(net124),
    .B1(net115),
    .B2(_03172_),
    .X(_02101_));
 sky130_fd_sc_hd__mux2_4 _13020_ (.A0(_05941_),
    .A1(\core_pipeline.execute_to_memory_csr_data[25] ),
    .S(net498),
    .X(_03173_));
 sky130_fd_sc_hd__a22o_1 _13021_ (.A1(net296),
    .A2(net117),
    .B1(_03173_),
    .B2(net240),
    .X(_03174_));
 sky130_fd_sc_hd__a22o_1 _13022_ (.A1(\core_pipeline.decode_to_execute_rs1_bypass[25] ),
    .A2(net124),
    .B1(net115),
    .B2(_03174_),
    .X(_02102_));
 sky130_fd_sc_hd__mux2_4 _13023_ (.A0(_05945_),
    .A1(\core_pipeline.execute_to_memory_csr_data[26] ),
    .S(net498),
    .X(_03175_));
 sky130_fd_sc_hd__a22o_1 _13024_ (.A1(net294),
    .A2(net117),
    .B1(_03175_),
    .B2(net240),
    .X(_03176_));
 sky130_fd_sc_hd__a22o_1 _13025_ (.A1(\core_pipeline.decode_to_execute_rs1_bypass[26] ),
    .A2(net122),
    .B1(net115),
    .B2(_03176_),
    .X(_02103_));
 sky130_fd_sc_hd__mux2_4 _13026_ (.A0(_05949_),
    .A1(\core_pipeline.execute_to_memory_csr_data[27] ),
    .S(net498),
    .X(_03177_));
 sky130_fd_sc_hd__a22o_1 _13027_ (.A1(_04003_),
    .A2(net118),
    .B1(_03177_),
    .B2(net239),
    .X(_03178_));
 sky130_fd_sc_hd__a22o_1 _13028_ (.A1(\core_pipeline.decode_to_execute_rs1_bypass[27] ),
    .A2(net133),
    .B1(net116),
    .B2(_03178_),
    .X(_02104_));
 sky130_fd_sc_hd__mux2_4 _13029_ (.A0(_05953_),
    .A1(\core_pipeline.execute_to_memory_csr_data[28] ),
    .S(net498),
    .X(_03179_));
 sky130_fd_sc_hd__a22o_1 _13030_ (.A1(_04006_),
    .A2(net118),
    .B1(_03179_),
    .B2(net239),
    .X(_03180_));
 sky130_fd_sc_hd__a22o_1 _13031_ (.A1(\core_pipeline.decode_to_execute_rs1_bypass[28] ),
    .A2(net131),
    .B1(net116),
    .B2(_03180_),
    .X(_02105_));
 sky130_fd_sc_hd__mux2_4 _13032_ (.A0(_05957_),
    .A1(\core_pipeline.execute_to_memory_csr_data[29] ),
    .S(net499),
    .X(_03181_));
 sky130_fd_sc_hd__a22o_1 _13033_ (.A1(net288),
    .A2(net118),
    .B1(_03181_),
    .B2(_03114_),
    .X(_03182_));
 sky130_fd_sc_hd__a22o_1 _13034_ (.A1(\core_pipeline.decode_to_execute_rs1_bypass[29] ),
    .A2(net130),
    .B1(net116),
    .B2(_03182_),
    .X(_02106_));
 sky130_fd_sc_hd__mux2_4 _13035_ (.A0(_05961_),
    .A1(\core_pipeline.execute_to_memory_csr_data[30] ),
    .S(net499),
    .X(_03183_));
 sky130_fd_sc_hd__a22o_1 _13036_ (.A1(_04012_),
    .A2(net118),
    .B1(_03183_),
    .B2(net239),
    .X(_03184_));
 sky130_fd_sc_hd__a22o_1 _13037_ (.A1(\core_pipeline.decode_to_execute_rs1_bypass[30] ),
    .A2(net125),
    .B1(net116),
    .B2(_03184_),
    .X(_02107_));
 sky130_fd_sc_hd__mux2_2 _13038_ (.A0(_05965_),
    .A1(\core_pipeline.execute_to_memory_csr_data[31] ),
    .S(net499),
    .X(_03185_));
 sky130_fd_sc_hd__a22o_1 _13039_ (.A1(_04015_),
    .A2(net118),
    .B1(_03185_),
    .B2(net239),
    .X(_03186_));
 sky130_fd_sc_hd__a22o_1 _13040_ (.A1(\core_pipeline.decode_to_execute_rs1_bypass[31] ),
    .A2(net133),
    .B1(net116),
    .B2(_03186_),
    .X(_02108_));
 sky130_fd_sc_hd__a21oi_4 _13041_ (.A1(net460),
    .A2(_04683_),
    .B1(net130),
    .Y(_03187_));
 sky130_fd_sc_hd__inv_2 _13042_ (.A(net114),
    .Y(_03188_));
 sky130_fd_sc_hd__o21ai_1 _13043_ (.A1(net513),
    .A2(_04684_),
    .B1(_03112_),
    .Y(_03189_));
 sky130_fd_sc_hd__o211a_2 _13044_ (.A1(_03492_),
    .A2(_03112_),
    .B1(_03189_),
    .C1(_03488_),
    .X(_03190_));
 sky130_fd_sc_hd__a22oi_1 _13045_ (.A1(net517),
    .A2(_04468_),
    .B1(_04936_),
    .B2(net524),
    .Y(_03191_));
 sky130_fd_sc_hd__o221a_1 _13046_ (.A1(net565),
    .A2(_03913_),
    .B1(_03914_),
    .B2(net542),
    .C1(_03191_),
    .X(_03192_));
 sky130_fd_sc_hd__a22oi_1 _13047_ (.A1(net512),
    .A2(_03912_),
    .B1(_03913_),
    .B2(net565),
    .Y(_03193_));
 sky130_fd_sc_hd__o2bb2a_1 _13048_ (.A1_N(net542),
    .A2_N(_03914_),
    .B1(_04468_),
    .B2(net517),
    .X(_03194_));
 sky130_fd_sc_hd__o221a_1 _13049_ (.A1(net512),
    .A2(_03912_),
    .B1(_04936_),
    .B2(net524),
    .C1(_03194_),
    .X(_03195_));
 sky130_fd_sc_hd__and3_1 _13050_ (.A(_03192_),
    .B(_03193_),
    .C(_03195_),
    .X(_03196_));
 sky130_fd_sc_hd__and2b_4 _13051_ (.A_N(net263),
    .B(_03196_),
    .X(_03197_));
 sky130_fd_sc_hd__a22o_1 _13052_ (.A1(_03115_),
    .A2(net264),
    .B1(net119),
    .B2(_03922_),
    .X(_03198_));
 sky130_fd_sc_hd__a22o_1 _13053_ (.A1(\core_pipeline.decode_to_execute_rs2_bypass[0] ),
    .A2(net122),
    .B1(net113),
    .B2(_03198_),
    .X(_02109_));
 sky130_fd_sc_hd__a22o_1 _13054_ (.A1(_03125_),
    .A2(net263),
    .B1(net120),
    .B2(_03925_),
    .X(_03199_));
 sky130_fd_sc_hd__a22o_1 _13055_ (.A1(\core_pipeline.decode_to_execute_rs2_bypass[1] ),
    .A2(net125),
    .B1(net114),
    .B2(_03199_),
    .X(_02110_));
 sky130_fd_sc_hd__a22o_1 _13056_ (.A1(_03127_),
    .A2(net263),
    .B1(net120),
    .B2(_03928_),
    .X(_03200_));
 sky130_fd_sc_hd__a22o_1 _13057_ (.A1(\core_pipeline.decode_to_execute_rs2_bypass[2] ),
    .A2(net130),
    .B1(net114),
    .B2(_03200_),
    .X(_02111_));
 sky130_fd_sc_hd__a22o_1 _13058_ (.A1(_03129_),
    .A2(net264),
    .B1(net119),
    .B2(_03931_),
    .X(_03201_));
 sky130_fd_sc_hd__a22o_1 _13059_ (.A1(\core_pipeline.decode_to_execute_rs2_bypass[3] ),
    .A2(net121),
    .B1(net113),
    .B2(_03201_),
    .X(_02112_));
 sky130_fd_sc_hd__a22o_1 _13060_ (.A1(_03131_),
    .A2(net264),
    .B1(net119),
    .B2(_03934_),
    .X(_03202_));
 sky130_fd_sc_hd__a22o_1 _13061_ (.A1(\core_pipeline.decode_to_execute_rs2_bypass[4] ),
    .A2(net121),
    .B1(net113),
    .B2(_03202_),
    .X(_02113_));
 sky130_fd_sc_hd__a22o_1 _13062_ (.A1(_03133_),
    .A2(net263),
    .B1(net120),
    .B2(net339),
    .X(_03203_));
 sky130_fd_sc_hd__a22o_1 _13063_ (.A1(\core_pipeline.decode_to_execute_rs2_bypass[5] ),
    .A2(net124),
    .B1(net114),
    .B2(_03203_),
    .X(_02114_));
 sky130_fd_sc_hd__a22o_1 _13064_ (.A1(_03135_),
    .A2(net263),
    .B1(net119),
    .B2(_03940_),
    .X(_03204_));
 sky130_fd_sc_hd__a22o_1 _13065_ (.A1(\core_pipeline.decode_to_execute_rs2_bypass[6] ),
    .A2(net125),
    .B1(net113),
    .B2(_03204_),
    .X(_02115_));
 sky130_fd_sc_hd__a22o_1 _13066_ (.A1(_03137_),
    .A2(net264),
    .B1(net119),
    .B2(net333),
    .X(_03205_));
 sky130_fd_sc_hd__a22o_1 _13067_ (.A1(\core_pipeline.decode_to_execute_rs2_bypass[7] ),
    .A2(net126),
    .B1(net113),
    .B2(_03205_),
    .X(_02116_));
 sky130_fd_sc_hd__a22o_1 _13068_ (.A1(_03139_),
    .A2(net264),
    .B1(net119),
    .B2(_03946_),
    .X(_03206_));
 sky130_fd_sc_hd__a22o_1 _13069_ (.A1(\core_pipeline.decode_to_execute_rs2_bypass[8] ),
    .A2(net124),
    .B1(net113),
    .B2(_03206_),
    .X(_02117_));
 sky130_fd_sc_hd__a22o_1 _13070_ (.A1(_03141_),
    .A2(net264),
    .B1(net119),
    .B2(net330),
    .X(_03207_));
 sky130_fd_sc_hd__a22o_1 _13071_ (.A1(\core_pipeline.decode_to_execute_rs2_bypass[9] ),
    .A2(net121),
    .B1(net113),
    .B2(_03207_),
    .X(_02118_));
 sky130_fd_sc_hd__a22o_1 _13072_ (.A1(_03143_),
    .A2(net264),
    .B1(net119),
    .B2(net328),
    .X(_03208_));
 sky130_fd_sc_hd__a22o_1 _13073_ (.A1(\core_pipeline.decode_to_execute_rs2_bypass[10] ),
    .A2(net122),
    .B1(net113),
    .B2(_03208_),
    .X(_02119_));
 sky130_fd_sc_hd__a22o_1 _13074_ (.A1(_03145_),
    .A2(net264),
    .B1(net119),
    .B2(net326),
    .X(_03209_));
 sky130_fd_sc_hd__a22o_1 _13075_ (.A1(\core_pipeline.decode_to_execute_rs2_bypass[11] ),
    .A2(net121),
    .B1(net113),
    .B2(_03209_),
    .X(_02120_));
 sky130_fd_sc_hd__a22o_1 _13076_ (.A1(_03147_),
    .A2(net264),
    .B1(net119),
    .B2(_03958_),
    .X(_03210_));
 sky130_fd_sc_hd__a22o_1 _13077_ (.A1(\core_pipeline.decode_to_execute_rs2_bypass[12] ),
    .A2(net121),
    .B1(net113),
    .B2(_03210_),
    .X(_02121_));
 sky130_fd_sc_hd__a22o_1 _13078_ (.A1(_03149_),
    .A2(net264),
    .B1(net119),
    .B2(net322),
    .X(_03211_));
 sky130_fd_sc_hd__a22o_1 _13079_ (.A1(\core_pipeline.decode_to_execute_rs2_bypass[13] ),
    .A2(net122),
    .B1(net113),
    .B2(_03211_),
    .X(_02122_));
 sky130_fd_sc_hd__a22o_1 _13080_ (.A1(_03151_),
    .A2(net264),
    .B1(net119),
    .B2(net320),
    .X(_03212_));
 sky130_fd_sc_hd__a22o_1 _13081_ (.A1(\core_pipeline.decode_to_execute_rs2_bypass[14] ),
    .A2(net121),
    .B1(net113),
    .B2(_03212_),
    .X(_02123_));
 sky130_fd_sc_hd__a22o_1 _13082_ (.A1(_03153_),
    .A2(net264),
    .B1(net119),
    .B2(net318),
    .X(_03213_));
 sky130_fd_sc_hd__a22o_1 _13083_ (.A1(\core_pipeline.decode_to_execute_rs2_bypass[15] ),
    .A2(net123),
    .B1(net113),
    .B2(_03213_),
    .X(_02124_));
 sky130_fd_sc_hd__a22o_1 _13084_ (.A1(_03155_),
    .A2(net264),
    .B1(net119),
    .B2(_03970_),
    .X(_03214_));
 sky130_fd_sc_hd__a22o_1 _13085_ (.A1(\core_pipeline.decode_to_execute_rs2_bypass[16] ),
    .A2(net124),
    .B1(net113),
    .B2(_03214_),
    .X(_02125_));
 sky130_fd_sc_hd__a22o_1 _13086_ (.A1(_03157_),
    .A2(net263),
    .B1(net120),
    .B2(net314),
    .X(_03215_));
 sky130_fd_sc_hd__a22o_1 _13087_ (.A1(\core_pipeline.decode_to_execute_rs2_bypass[17] ),
    .A2(net131),
    .B1(net114),
    .B2(_03215_),
    .X(_02126_));
 sky130_fd_sc_hd__a22o_1 _13088_ (.A1(_03159_),
    .A2(net263),
    .B1(net120),
    .B2(_03976_),
    .X(_03216_));
 sky130_fd_sc_hd__a22o_1 _13089_ (.A1(\core_pipeline.decode_to_execute_rs2_bypass[18] ),
    .A2(net132),
    .B1(net114),
    .B2(_03216_),
    .X(_02127_));
 sky130_fd_sc_hd__a22o_1 _13090_ (.A1(_03161_),
    .A2(net263),
    .B1(net120),
    .B2(_03979_),
    .X(_03217_));
 sky130_fd_sc_hd__a22o_1 _13091_ (.A1(\core_pipeline.decode_to_execute_rs2_bypass[19] ),
    .A2(net130),
    .B1(net114),
    .B2(_03217_),
    .X(_02128_));
 sky130_fd_sc_hd__a22o_1 _13092_ (.A1(_03163_),
    .A2(net263),
    .B1(net120),
    .B2(net307),
    .X(_03218_));
 sky130_fd_sc_hd__a22o_1 _13093_ (.A1(\core_pipeline.decode_to_execute_rs2_bypass[20] ),
    .A2(net131),
    .B1(net114),
    .B2(_03218_),
    .X(_02129_));
 sky130_fd_sc_hd__a22o_1 _13094_ (.A1(_03165_),
    .A2(net263),
    .B1(net120),
    .B2(_03985_),
    .X(_03219_));
 sky130_fd_sc_hd__a22o_1 _13095_ (.A1(\core_pipeline.decode_to_execute_rs2_bypass[21] ),
    .A2(net132),
    .B1(net114),
    .B2(_03219_),
    .X(_02130_));
 sky130_fd_sc_hd__a22o_1 _13096_ (.A1(_03167_),
    .A2(net263),
    .B1(net120),
    .B2(_03988_),
    .X(_03220_));
 sky130_fd_sc_hd__a22o_1 _13097_ (.A1(\core_pipeline.decode_to_execute_rs2_bypass[22] ),
    .A2(net130),
    .B1(net114),
    .B2(_03220_),
    .X(_02131_));
 sky130_fd_sc_hd__a22o_1 _13098_ (.A1(_03169_),
    .A2(net263),
    .B1(net120),
    .B2(net300),
    .X(_03221_));
 sky130_fd_sc_hd__a22o_1 _13099_ (.A1(\core_pipeline.decode_to_execute_rs2_bypass[23] ),
    .A2(net125),
    .B1(net114),
    .B2(_03221_),
    .X(_02132_));
 sky130_fd_sc_hd__a22o_1 _13100_ (.A1(_03171_),
    .A2(net264),
    .B1(net119),
    .B2(net298),
    .X(_03222_));
 sky130_fd_sc_hd__a22o_1 _13101_ (.A1(\core_pipeline.decode_to_execute_rs2_bypass[24] ),
    .A2(net124),
    .B1(net113),
    .B2(_03222_),
    .X(_02133_));
 sky130_fd_sc_hd__a22o_1 _13102_ (.A1(_03173_),
    .A2(net264),
    .B1(net119),
    .B2(net296),
    .X(_03223_));
 sky130_fd_sc_hd__a22o_1 _13103_ (.A1(\core_pipeline.decode_to_execute_rs2_bypass[25] ),
    .A2(net124),
    .B1(net113),
    .B2(_03223_),
    .X(_02134_));
 sky130_fd_sc_hd__a22o_1 _13104_ (.A1(_03175_),
    .A2(net264),
    .B1(net119),
    .B2(net294),
    .X(_03224_));
 sky130_fd_sc_hd__a22o_1 _13105_ (.A1(\core_pipeline.decode_to_execute_rs2_bypass[26] ),
    .A2(net122),
    .B1(net113),
    .B2(_03224_),
    .X(_02135_));
 sky130_fd_sc_hd__a22o_1 _13106_ (.A1(_03177_),
    .A2(net263),
    .B1(net120),
    .B2(_04003_),
    .X(_03225_));
 sky130_fd_sc_hd__a22o_1 _13107_ (.A1(\core_pipeline.decode_to_execute_rs2_bypass[27] ),
    .A2(net132),
    .B1(net114),
    .B2(_03225_),
    .X(_02136_));
 sky130_fd_sc_hd__a22o_1 _13108_ (.A1(_03179_),
    .A2(_03190_),
    .B1(net120),
    .B2(_04006_),
    .X(_03226_));
 sky130_fd_sc_hd__a22o_1 _13109_ (.A1(\core_pipeline.decode_to_execute_rs2_bypass[28] ),
    .A2(net130),
    .B1(net114),
    .B2(_03226_),
    .X(_02137_));
 sky130_fd_sc_hd__a22o_1 _13110_ (.A1(_03181_),
    .A2(net263),
    .B1(net120),
    .B2(net288),
    .X(_03227_));
 sky130_fd_sc_hd__a22o_1 _13111_ (.A1(\core_pipeline.decode_to_execute_rs2_bypass[29] ),
    .A2(net130),
    .B1(net114),
    .B2(_03227_),
    .X(_02138_));
 sky130_fd_sc_hd__a22o_1 _13112_ (.A1(_03183_),
    .A2(net263),
    .B1(net120),
    .B2(_04012_),
    .X(_03228_));
 sky130_fd_sc_hd__a22o_1 _13113_ (.A1(\core_pipeline.decode_to_execute_rs2_bypass[30] ),
    .A2(net125),
    .B1(net114),
    .B2(_03228_),
    .X(_02139_));
 sky130_fd_sc_hd__a22o_1 _13114_ (.A1(_03185_),
    .A2(net263),
    .B1(net120),
    .B2(_04015_),
    .X(_03229_));
 sky130_fd_sc_hd__a22o_1 _13115_ (.A1(\core_pipeline.decode_to_execute_rs2_bypass[31] ),
    .A2(net132),
    .B1(net114),
    .B2(_03229_),
    .X(_02140_));
 sky130_fd_sc_hd__and3b_1 _13116_ (.A_N(net239),
    .B(_03121_),
    .C(net116),
    .X(_03230_));
 sky130_fd_sc_hd__o21ba_1 _13117_ (.A1(net489),
    .A2(net147),
    .B1_N(_03230_),
    .X(_02141_));
 sky130_fd_sc_hd__o32a_1 _13118_ (.A1(_03188_),
    .A2(net263),
    .A3(_03196_),
    .B1(net147),
    .B2(net487),
    .X(_02142_));
 sky130_fd_sc_hd__mux2_1 _13119_ (.A0(\core_pipeline.fetch_to_decode_instruction[13] ),
    .A1(\core_pipeline.decode_to_execute_cmp_function[1] ),
    .S(net124),
    .X(_02143_));
 sky130_fd_sc_hd__mux2_1 _13120_ (.A0(\core_pipeline.fetch_to_decode_instruction[14] ),
    .A1(\core_pipeline.decode_to_execute_cmp_function[2] ),
    .S(net126),
    .X(_02144_));
 sky130_fd_sc_hd__o21a_1 _13121_ (.A1(\core_pipeline.decode_to_execute_jump ),
    .A2(net143),
    .B1(_04629_),
    .X(_02145_));
 sky130_fd_sc_hd__o22a_1 _13122_ (.A1(\core_pipeline.decode_to_execute_branch ),
    .A2(net143),
    .B1(_03445_),
    .B2(_04629_),
    .X(_02146_));
 sky130_fd_sc_hd__nor2_1 _13123_ (.A(net465),
    .B(net427),
    .Y(_03231_));
 sky130_fd_sc_hd__o2bb2a_1 _13124_ (.A1_N(_03328_),
    .A2_N(_04693_),
    .B1(_04709_),
    .B2(_03231_),
    .X(_03232_));
 sky130_fd_sc_hd__or3b_1 _13125_ (.A(_04682_),
    .B(net513),
    .C_N(\core_pipeline.decode_to_csr_read_address[7] ),
    .X(_03233_));
 sky130_fd_sc_hd__a211o_1 _13126_ (.A1(\core_pipeline.decode_to_csr_read_address[6] ),
    .A2(_03233_),
    .B1(_04686_),
    .C1(\core_pipeline.decode_to_csr_read_address[5] ),
    .X(_03234_));
 sky130_fd_sc_hd__or4b_1 _13127_ (.A(\core_pipeline.decode_to_csr_read_address[7] ),
    .B(\core_pipeline.decode_to_csr_read_address[6] ),
    .C(_04692_),
    .D_N(\core_pipeline.decode_to_csr_read_address[5] ),
    .X(_03235_));
 sky130_fd_sc_hd__o211a_1 _13128_ (.A1(net517),
    .A2(_03232_),
    .B1(_03234_),
    .C1(_03235_),
    .X(_03236_));
 sky130_fd_sc_hd__nor2_1 _13129_ (.A(net132),
    .B(_03236_),
    .Y(_03237_));
 sky130_fd_sc_hd__a211o_1 _13130_ (.A1(net427),
    .A2(_04694_),
    .B1(net277),
    .C1(net362),
    .X(_03238_));
 sky130_fd_sc_hd__nor3_1 _13131_ (.A(_03330_),
    .B(\core_pipeline.decode_to_csr_read_address[7] ),
    .C(_04685_),
    .Y(_03239_));
 sky130_fd_sc_hd__a2bb2o_1 _13132_ (.A1_N(\core_pipeline.decode_to_csr_read_address[9] ),
    .A2_N(\core_pipeline.decode_to_csr_read_address[8] ),
    .B1(_03238_),
    .B2(_03239_),
    .X(_03240_));
 sky130_fd_sc_hd__nor3_1 _13133_ (.A(\core_pipeline.decode_to_csr_read_address[5] ),
    .B(\core_pipeline.decode_to_csr_read_address[6] ),
    .C(_04702_),
    .Y(_03241_));
 sky130_fd_sc_hd__and3_1 _13134_ (.A(net146),
    .B(_03240_),
    .C(_03241_),
    .X(_03242_));
 sky130_fd_sc_hd__a211o_1 _13135_ (.A1(\core_pipeline.decode_to_execute_csr_readable ),
    .A2(net133),
    .B1(_03237_),
    .C1(_03242_),
    .X(_02147_));
 sky130_fd_sc_hd__a21o_1 _13136_ (.A1(\core_pipeline.decode_to_execute_csr_writeable ),
    .A2(net133),
    .B1(_03237_),
    .X(_02148_));
 sky130_fd_sc_hd__mux2_1 _13137_ (.A0(\core_pipeline.decode_to_execute_load ),
    .A1(_04626_),
    .S(net142),
    .X(_02149_));
 sky130_fd_sc_hd__mux2_1 _13138_ (.A0(\core_pipeline.decode_to_execute_store ),
    .A1(_04664_),
    .S(net142),
    .X(_02150_));
 sky130_fd_sc_hd__mux2_1 _13139_ (.A0(\core_pipeline.fetch_to_decode_instruction[12] ),
    .A1(\core_pipeline.decode_to_execute_cmp_function[0] ),
    .S(net125),
    .X(_02151_));
 sky130_fd_sc_hd__mux2_1 _13140_ (.A0(_03313_),
    .A1(\core_pipeline.decode_to_execute_load_signed ),
    .S(net127),
    .X(_02152_));
 sky130_fd_sc_hd__a2bb2o_1 _13141_ (.A1_N(_04716_),
    .A2_N(_04931_),
    .B1(\core_pipeline.decode_to_execute_mret ),
    .B2(net132),
    .X(_02153_));
 sky130_fd_sc_hd__a32o_1 _13142_ (.A1(_03632_),
    .A2(_04911_),
    .A3(_04922_),
    .B1(net132),
    .B2(\core_pipeline.decode_to_execute_wfi ),
    .X(_02154_));
 sky130_fd_sc_hd__mux2_1 _13143_ (.A0(net564),
    .A1(\core_pipeline.decode_to_execute_csr_address[0] ),
    .S(net134),
    .X(_02155_));
 sky130_fd_sc_hd__mux2_1 _13144_ (.A0(net541),
    .A1(\core_pipeline.decode_to_execute_csr_address[1] ),
    .S(net134),
    .X(_02156_));
 sky130_fd_sc_hd__mux2_1 _13145_ (.A0(net524),
    .A1(\core_pipeline.decode_to_execute_csr_address[2] ),
    .S(net134),
    .X(_02157_));
 sky130_fd_sc_hd__mux2_1 _13146_ (.A0(net517),
    .A1(\core_pipeline.decode_to_execute_csr_address[3] ),
    .S(net134),
    .X(_02158_));
 sky130_fd_sc_hd__mux2_1 _13147_ (.A0(net513),
    .A1(\core_pipeline.decode_to_execute_csr_address[4] ),
    .S(net134),
    .X(_02159_));
 sky130_fd_sc_hd__mux2_1 _13148_ (.A0(\core_pipeline.decode_to_csr_read_address[5] ),
    .A1(\core_pipeline.decode_to_execute_csr_address[5] ),
    .S(net134),
    .X(_02160_));
 sky130_fd_sc_hd__mux2_1 _13149_ (.A0(\core_pipeline.decode_to_csr_read_address[6] ),
    .A1(\core_pipeline.decode_to_execute_csr_address[6] ),
    .S(net135),
    .X(_02161_));
 sky130_fd_sc_hd__mux2_1 _13150_ (.A0(\core_pipeline.decode_to_csr_read_address[7] ),
    .A1(\core_pipeline.decode_to_execute_csr_address[7] ),
    .S(net134),
    .X(_02162_));
 sky130_fd_sc_hd__mux2_1 _13151_ (.A0(\core_pipeline.decode_to_csr_read_address[8] ),
    .A1(\core_pipeline.decode_to_execute_csr_address[8] ),
    .S(net134),
    .X(_02163_));
 sky130_fd_sc_hd__mux2_1 _13152_ (.A0(\core_pipeline.decode_to_csr_read_address[9] ),
    .A1(\core_pipeline.decode_to_execute_csr_address[9] ),
    .S(net134),
    .X(_02164_));
 sky130_fd_sc_hd__mux2_1 _13153_ (.A0(\core_pipeline.decode_to_csr_read_address[10] ),
    .A1(\core_pipeline.decode_to_execute_csr_address[10] ),
    .S(net134),
    .X(_02165_));
 sky130_fd_sc_hd__mux2_1 _13154_ (.A0(\core_pipeline.decode_to_csr_read_address[11] ),
    .A1(\core_pipeline.decode_to_execute_csr_address[11] ),
    .S(net134),
    .X(_02166_));
 sky130_fd_sc_hd__and3_4 _13155_ (.A(\core_pipeline.decode_to_execute_alu_function[2] ),
    .B(\core_pipeline.decode_to_execute_alu_function[1] ),
    .C(\core_pipeline.decode_to_execute_alu_function[0] ),
    .X(_03243_));
 sky130_fd_sc_hd__nand3_4 _13156_ (.A(\core_pipeline.decode_to_execute_alu_function[2] ),
    .B(\core_pipeline.decode_to_execute_alu_function[1] ),
    .C(\core_pipeline.decode_to_execute_alu_function[0] ),
    .Y(_03244_));
 sky130_fd_sc_hd__o221a_1 _13157_ (.A1(net631),
    .A2(_04495_),
    .B1(_04503_),
    .B2(_06052_),
    .C1(_03243_),
    .X(_03245_));
 sky130_fd_sc_hd__a21o_1 _13158_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_and_clr[0] ),
    .A2(net406),
    .B1(_03245_),
    .X(_02167_));
 sky130_fd_sc_hd__nand2_1 _13159_ (.A(net631),
    .B(_04502_),
    .Y(_03246_));
 sky130_fd_sc_hd__o21a_1 _13160_ (.A1(net631),
    .A2(_04502_),
    .B1(_03243_),
    .X(_03247_));
 sky130_fd_sc_hd__a32o_1 _13161_ (.A1(net379),
    .A2(_03246_),
    .A3(_03247_),
    .B1(net406),
    .B2(\core_pipeline.pipeline_execute.ex_alu.result_and_clr[1] ),
    .X(_02168_));
 sky130_fd_sc_hd__nand2_1 _13162_ (.A(net459),
    .B(_04511_),
    .Y(_03248_));
 sky130_fd_sc_hd__o211a_1 _13163_ (.A1(net459),
    .A2(_04511_),
    .B1(_03243_),
    .C1(net384),
    .X(_03249_));
 sky130_fd_sc_hd__a22o_1 _13164_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_and_clr[2] ),
    .A2(net406),
    .B1(_03248_),
    .B2(_03249_),
    .X(_02169_));
 sky130_fd_sc_hd__nand2_1 _13165_ (.A(net459),
    .B(_04517_),
    .Y(_03250_));
 sky130_fd_sc_hd__o211a_1 _13166_ (.A1(net459),
    .A2(_04517_),
    .B1(_03243_),
    .C1(net395),
    .X(_03251_));
 sky130_fd_sc_hd__a22o_1 _13167_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_and_clr[3] ),
    .A2(net406),
    .B1(_03250_),
    .B2(_03251_),
    .X(_02170_));
 sky130_fd_sc_hd__nand2_1 _13168_ (.A(net631),
    .B(_04522_),
    .Y(_03252_));
 sky130_fd_sc_hd__o211a_1 _13169_ (.A1(net631),
    .A2(_04522_),
    .B1(_03243_),
    .C1(net391),
    .X(_03253_));
 sky130_fd_sc_hd__a22o_1 _13170_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_and_clr[4] ),
    .A2(net406),
    .B1(_03252_),
    .B2(_03253_),
    .X(_02171_));
 sky130_fd_sc_hd__nor2_1 _13171_ (.A(net631),
    .B(_04530_),
    .Y(_03254_));
 sky130_fd_sc_hd__a211o_1 _13172_ (.A1(net631),
    .A2(_04530_),
    .B1(_05666_),
    .C1(net406),
    .X(_03255_));
 sky130_fd_sc_hd__a2bb2o_1 _13173_ (.A1_N(_03254_),
    .A2_N(_03255_),
    .B1(\core_pipeline.pipeline_execute.ex_alu.result_and_clr[5] ),
    .B2(net406),
    .X(_02172_));
 sky130_fd_sc_hd__a21oi_1 _13174_ (.A1(net632),
    .A2(_04538_),
    .B1(_05662_),
    .Y(_03256_));
 sky130_fd_sc_hd__o21a_1 _13175_ (.A1(net632),
    .A2(_04538_),
    .B1(_03243_),
    .X(_03257_));
 sky130_fd_sc_hd__a22o_1 _13176_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_and_clr[6] ),
    .A2(net406),
    .B1(_03256_),
    .B2(_03257_),
    .X(_02173_));
 sky130_fd_sc_hd__nor2_1 _13177_ (.A(_05657_),
    .B(net406),
    .Y(_03258_));
 sky130_fd_sc_hd__xnor2_1 _13178_ (.A(net632),
    .B(_04545_),
    .Y(_03259_));
 sky130_fd_sc_hd__a22o_1 _13179_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_and_clr[7] ),
    .A2(net406),
    .B1(_03258_),
    .B2(_03259_),
    .X(_02174_));
 sky130_fd_sc_hd__a21oi_1 _13180_ (.A1(net635),
    .A2(_04554_),
    .B1(_05633_),
    .Y(_03260_));
 sky130_fd_sc_hd__a21oi_1 _13181_ (.A1(net459),
    .A2(_04553_),
    .B1(net405),
    .Y(_03261_));
 sky130_fd_sc_hd__a22o_1 _13182_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_and_clr[8] ),
    .A2(net405),
    .B1(_03260_),
    .B2(_03261_),
    .X(_02175_));
 sky130_fd_sc_hd__nor2_1 _13183_ (.A(net635),
    .B(_04566_),
    .Y(_03262_));
 sky130_fd_sc_hd__a211o_1 _13184_ (.A1(net635),
    .A2(_04566_),
    .B1(_05636_),
    .C1(net405),
    .X(_03263_));
 sky130_fd_sc_hd__a2bb2o_1 _13185_ (.A1_N(_03262_),
    .A2_N(_03263_),
    .B1(\core_pipeline.pipeline_execute.ex_alu.result_and_clr[9] ),
    .B2(net405),
    .X(_02176_));
 sky130_fd_sc_hd__a21oi_1 _13186_ (.A1(net635),
    .A2(_04574_),
    .B1(_05651_),
    .Y(_03264_));
 sky130_fd_sc_hd__o21a_1 _13187_ (.A1(net635),
    .A2(_04574_),
    .B1(_03243_),
    .X(_03265_));
 sky130_fd_sc_hd__a22o_1 _13188_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_and_clr[10] ),
    .A2(net405),
    .B1(_03264_),
    .B2(_03265_),
    .X(_02177_));
 sky130_fd_sc_hd__nor2_1 _13189_ (.A(net635),
    .B(_04582_),
    .Y(_03266_));
 sky130_fd_sc_hd__a211o_1 _13190_ (.A1(net635),
    .A2(_04582_),
    .B1(_05639_),
    .C1(net405),
    .X(_03267_));
 sky130_fd_sc_hd__a2bb2o_1 _13191_ (.A1_N(_03266_),
    .A2_N(_03267_),
    .B1(\core_pipeline.pipeline_execute.ex_alu.result_and_clr[11] ),
    .B2(net405),
    .X(_02178_));
 sky130_fd_sc_hd__a21oi_1 _13192_ (.A1(_03423_),
    .A2(net371),
    .B1(net404),
    .Y(_03268_));
 sky130_fd_sc_hd__o211a_1 _13193_ (.A1(_03423_),
    .A2(net371),
    .B1(_05642_),
    .C1(_03268_),
    .X(_03269_));
 sky130_fd_sc_hd__a21o_1 _13194_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_and_clr[12] ),
    .A2(net404),
    .B1(_03269_),
    .X(_02179_));
 sky130_fd_sc_hd__nand2_1 _13195_ (.A(net459),
    .B(_04599_),
    .Y(_03270_));
 sky130_fd_sc_hd__o211a_1 _13196_ (.A1(_03423_),
    .A2(_04599_),
    .B1(_05623_),
    .C1(_03243_),
    .X(_03271_));
 sky130_fd_sc_hd__a22o_1 _13197_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_and_clr[13] ),
    .A2(net405),
    .B1(_03270_),
    .B2(_03271_),
    .X(_02180_));
 sky130_fd_sc_hd__and2_1 _13198_ (.A(\core_pipeline.pipeline_execute.ex_alu.result_and_clr[14] ),
    .B(net404),
    .X(_03272_));
 sky130_fd_sc_hd__or2_1 _13199_ (.A(net459),
    .B(_04608_),
    .X(_03273_));
 sky130_fd_sc_hd__a21oi_1 _13200_ (.A1(net459),
    .A2(_04608_),
    .B1(_05618_),
    .Y(_03274_));
 sky130_fd_sc_hd__a31o_1 _13201_ (.A1(_03243_),
    .A2(_03273_),
    .A3(_03274_),
    .B1(_03272_),
    .X(_02181_));
 sky130_fd_sc_hd__or2_1 _13202_ (.A(net634),
    .B(_04618_),
    .X(_03275_));
 sky130_fd_sc_hd__a21oi_1 _13203_ (.A1(net634),
    .A2(_04618_),
    .B1(net404),
    .Y(_03276_));
 sky130_fd_sc_hd__a32o_1 _13204_ (.A1(_05627_),
    .A2(_03275_),
    .A3(_03276_),
    .B1(net404),
    .B2(\core_pipeline.pipeline_execute.ex_alu.result_and_clr[15] ),
    .X(_02182_));
 sky130_fd_sc_hd__o21ba_1 _13205_ (.A1(net634),
    .A2(_05760_),
    .B1_N(_05758_),
    .X(_03277_));
 sky130_fd_sc_hd__a21oi_1 _13206_ (.A1(net634),
    .A2(_05760_),
    .B1(net404),
    .Y(_03278_));
 sky130_fd_sc_hd__a22o_1 _13207_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_and_clr[16] ),
    .A2(net404),
    .B1(_03277_),
    .B2(_03278_),
    .X(_02183_));
 sky130_fd_sc_hd__nor2_1 _13208_ (.A(net635),
    .B(_05748_),
    .Y(_03279_));
 sky130_fd_sc_hd__a211o_1 _13209_ (.A1(net634),
    .A2(_05748_),
    .B1(net405),
    .C1(_05745_),
    .X(_03280_));
 sky130_fd_sc_hd__a2bb2o_1 _13210_ (.A1_N(_03279_),
    .A2_N(_03280_),
    .B1(\core_pipeline.pipeline_execute.ex_alu.result_and_clr[17] ),
    .B2(net405),
    .X(_02184_));
 sky130_fd_sc_hd__a21oi_1 _13211_ (.A1(net634),
    .A2(_05781_),
    .B1(_05779_),
    .Y(_03281_));
 sky130_fd_sc_hd__o21a_1 _13212_ (.A1(net634),
    .A2(_05781_),
    .B1(_03243_),
    .X(_03282_));
 sky130_fd_sc_hd__a22o_1 _13213_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_and_clr[18] ),
    .A2(net404),
    .B1(_03281_),
    .B2(_03282_),
    .X(_02185_));
 sky130_fd_sc_hd__nor2_1 _13214_ (.A(_05786_),
    .B(net404),
    .Y(_03283_));
 sky130_fd_sc_hd__xnor2_1 _13215_ (.A(net634),
    .B(_05788_),
    .Y(_03284_));
 sky130_fd_sc_hd__a22o_1 _13216_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_and_clr[19] ),
    .A2(net405),
    .B1(_03283_),
    .B2(_03284_),
    .X(_02186_));
 sky130_fd_sc_hd__xnor2_1 _13217_ (.A(net459),
    .B(_05773_),
    .Y(_03285_));
 sky130_fd_sc_hd__nor2_1 _13218_ (.A(_05771_),
    .B(_03285_),
    .Y(_03286_));
 sky130_fd_sc_hd__mux2_1 _13219_ (.A0(\core_pipeline.pipeline_execute.ex_alu.result_and_clr[20] ),
    .A1(_03286_),
    .S(_03243_),
    .X(_02187_));
 sky130_fd_sc_hd__nor2_1 _13220_ (.A(net633),
    .B(_05765_),
    .Y(_03287_));
 sky130_fd_sc_hd__a211o_1 _13221_ (.A1(net633),
    .A2(_05765_),
    .B1(net404),
    .C1(_05763_),
    .X(_03288_));
 sky130_fd_sc_hd__a2bb2o_1 _13222_ (.A1_N(_03287_),
    .A2_N(_03288_),
    .B1(\core_pipeline.pipeline_execute.ex_alu.result_and_clr[21] ),
    .B2(net404),
    .X(_02188_));
 sky130_fd_sc_hd__nor2_1 _13223_ (.A(net633),
    .B(_05755_),
    .Y(_03289_));
 sky130_fd_sc_hd__a211o_1 _13224_ (.A1(net633),
    .A2(_05809_),
    .B1(net404),
    .C1(_03289_),
    .X(_03290_));
 sky130_fd_sc_hd__o21a_1 _13225_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_and_clr[22] ),
    .A2(_03243_),
    .B1(_03290_),
    .X(_02189_));
 sky130_fd_sc_hd__nor2_1 _13226_ (.A(net632),
    .B(_05740_),
    .Y(_03291_));
 sky130_fd_sc_hd__a211o_1 _13227_ (.A1(net632),
    .A2(_05740_),
    .B1(net406),
    .C1(_05738_),
    .X(_03292_));
 sky130_fd_sc_hd__a2bb2o_1 _13228_ (.A1_N(_03291_),
    .A2_N(_03292_),
    .B1(\core_pipeline.pipeline_execute.ex_alu.result_and_clr[23] ),
    .B2(net406),
    .X(_02190_));
 sky130_fd_sc_hd__nor2_1 _13229_ (.A(net635),
    .B(_05719_),
    .Y(_03293_));
 sky130_fd_sc_hd__a211o_1 _13230_ (.A1(net635),
    .A2(_05796_),
    .B1(net405),
    .C1(_03293_),
    .X(_03294_));
 sky130_fd_sc_hd__o21a_1 _13231_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_and_clr[24] ),
    .A2(_03243_),
    .B1(_03294_),
    .X(_02191_));
 sky130_fd_sc_hd__or2_1 _13232_ (.A(net634),
    .B(_05731_),
    .X(_03295_));
 sky130_fd_sc_hd__nand2_1 _13233_ (.A(net634),
    .B(_05731_),
    .Y(_03296_));
 sky130_fd_sc_hd__a31o_1 _13234_ (.A1(_05729_),
    .A2(_03295_),
    .A3(_03296_),
    .B1(net404),
    .X(_03297_));
 sky130_fd_sc_hd__o21a_1 _13235_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_and_clr[25] ),
    .A2(_03243_),
    .B1(_03297_),
    .X(_02192_));
 sky130_fd_sc_hd__nor2_1 _13236_ (.A(net633),
    .B(_05712_),
    .Y(_03298_));
 sky130_fd_sc_hd__a211o_1 _13237_ (.A1(net633),
    .A2(_05712_),
    .B1(net404),
    .C1(_05710_),
    .X(_03299_));
 sky130_fd_sc_hd__a2bb2o_1 _13238_ (.A1_N(_03298_),
    .A2_N(_03299_),
    .B1(\core_pipeline.pipeline_execute.ex_alu.result_and_clr[26] ),
    .B2(net404),
    .X(_02193_));
 sky130_fd_sc_hd__o21a_1 _13239_ (.A1(_03423_),
    .A2(net360),
    .B1(_05722_),
    .X(_03300_));
 sky130_fd_sc_hd__a21oi_1 _13240_ (.A1(net459),
    .A2(net360),
    .B1(net405),
    .Y(_03301_));
 sky130_fd_sc_hd__a22o_1 _13241_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_and_clr[27] ),
    .A2(net405),
    .B1(_03300_),
    .B2(_03301_),
    .X(_02194_));
 sky130_fd_sc_hd__nor2_1 _13242_ (.A(net632),
    .B(_05699_),
    .Y(_03302_));
 sky130_fd_sc_hd__a211o_1 _13243_ (.A1(net632),
    .A2(_05699_),
    .B1(net406),
    .C1(_05697_),
    .X(_03303_));
 sky130_fd_sc_hd__a2bb2o_1 _13244_ (.A1_N(_03302_),
    .A2_N(_03303_),
    .B1(\core_pipeline.pipeline_execute.ex_alu.result_and_clr[28] ),
    .B2(net406),
    .X(_02195_));
 sky130_fd_sc_hd__o21a_1 _13245_ (.A1(net459),
    .A2(_05704_),
    .B1(_05702_),
    .X(_03304_));
 sky130_fd_sc_hd__a21oi_1 _13246_ (.A1(net459),
    .A2(_05704_),
    .B1(net404),
    .Y(_03305_));
 sky130_fd_sc_hd__a22o_1 _13247_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_and_clr[29] ),
    .A2(net404),
    .B1(_03304_),
    .B2(_03305_),
    .X(_02196_));
 sky130_fd_sc_hd__a21oi_1 _13248_ (.A1(net632),
    .A2(_05687_),
    .B1(_05691_),
    .Y(_03306_));
 sky130_fd_sc_hd__o21a_1 _13249_ (.A1(net632),
    .A2(_05687_),
    .B1(_03243_),
    .X(_03307_));
 sky130_fd_sc_hd__a22o_1 _13250_ (.A1(\core_pipeline.pipeline_execute.ex_alu.result_and_clr[30] ),
    .A2(net406),
    .B1(_03306_),
    .B2(_03307_),
    .X(_02197_));
 sky130_fd_sc_hd__or2_1 _13251_ (.A(net631),
    .B(_05614_),
    .X(_03308_));
 sky130_fd_sc_hd__nor2_1 _13252_ (.A(_05612_),
    .B(net406),
    .Y(_03309_));
 sky130_fd_sc_hd__a32o_1 _13253_ (.A1(_06094_),
    .A2(_03308_),
    .A3(_03309_),
    .B1(net406),
    .B2(\core_pipeline.pipeline_execute.ex_alu.result_and_clr[31] ),
    .X(_02198_));
 sky130_fd_sc_hd__mux2_1 _13254_ (.A0(\core_pipeline.pipeline_fetch.pc[2] ),
    .A1(\core_pipeline.fetch_to_decode_pc[2] ),
    .S(net109),
    .X(_02199_));
 sky130_fd_sc_hd__mux2_1 _13255_ (.A0(\core_pipeline.pipeline_fetch.pc[3] ),
    .A1(\core_pipeline.fetch_to_decode_pc[3] ),
    .S(net109),
    .X(_02200_));
 sky130_fd_sc_hd__mux2_1 _13256_ (.A0(\core_pipeline.pipeline_fetch.pc[4] ),
    .A1(\core_pipeline.fetch_to_decode_pc[4] ),
    .S(net108),
    .X(_02201_));
 sky130_fd_sc_hd__mux2_1 _13257_ (.A0(\core_pipeline.pipeline_fetch.pc[5] ),
    .A1(\core_pipeline.fetch_to_decode_pc[5] ),
    .S(net108),
    .X(_02202_));
 sky130_fd_sc_hd__mux2_1 _13258_ (.A0(\core_pipeline.pipeline_fetch.pc[6] ),
    .A1(\core_pipeline.fetch_to_decode_pc[6] ),
    .S(net108),
    .X(_02203_));
 sky130_fd_sc_hd__mux2_1 _13259_ (.A0(\core_pipeline.pipeline_fetch.pc[7] ),
    .A1(\core_pipeline.fetch_to_decode_pc[7] ),
    .S(net109),
    .X(_02204_));
 sky130_fd_sc_hd__mux2_1 _13260_ (.A0(\core_pipeline.pipeline_fetch.pc[8] ),
    .A1(\core_pipeline.fetch_to_decode_pc[8] ),
    .S(net110),
    .X(_02205_));
 sky130_fd_sc_hd__mux2_1 _13261_ (.A0(\core_pipeline.pipeline_fetch.pc[9] ),
    .A1(\core_pipeline.fetch_to_decode_pc[9] ),
    .S(net112),
    .X(_02206_));
 sky130_fd_sc_hd__mux2_1 _13262_ (.A0(\core_pipeline.pipeline_fetch.pc[10] ),
    .A1(\core_pipeline.fetch_to_decode_pc[10] ),
    .S(net110),
    .X(_02207_));
 sky130_fd_sc_hd__mux2_1 _13263_ (.A0(\core_pipeline.pipeline_fetch.pc[11] ),
    .A1(\core_pipeline.fetch_to_decode_pc[11] ),
    .S(net110),
    .X(_02208_));
 sky130_fd_sc_hd__mux2_1 _13264_ (.A0(\core_pipeline.pipeline_fetch.pc[12] ),
    .A1(\core_pipeline.fetch_to_decode_pc[12] ),
    .S(net110),
    .X(_02209_));
 sky130_fd_sc_hd__mux2_1 _13265_ (.A0(\core_pipeline.pipeline_fetch.pc[13] ),
    .A1(\core_pipeline.fetch_to_decode_pc[13] ),
    .S(net110),
    .X(_02210_));
 sky130_fd_sc_hd__mux2_1 _13266_ (.A0(\core_pipeline.pipeline_fetch.pc[14] ),
    .A1(\core_pipeline.fetch_to_decode_pc[14] ),
    .S(net110),
    .X(_02211_));
 sky130_fd_sc_hd__mux2_1 _13267_ (.A0(\core_pipeline.pipeline_fetch.pc[15] ),
    .A1(\core_pipeline.fetch_to_decode_pc[15] ),
    .S(net110),
    .X(_02212_));
 sky130_fd_sc_hd__mux2_1 _13268_ (.A0(\core_pipeline.pipeline_fetch.pc[16] ),
    .A1(\core_pipeline.fetch_to_decode_pc[16] ),
    .S(net112),
    .X(_02213_));
 sky130_fd_sc_hd__mux2_1 _13269_ (.A0(\core_pipeline.pipeline_fetch.pc[17] ),
    .A1(\core_pipeline.fetch_to_decode_pc[17] ),
    .S(net111),
    .X(_02214_));
 sky130_fd_sc_hd__mux2_1 _13270_ (.A0(\core_pipeline.pipeline_fetch.pc[18] ),
    .A1(\core_pipeline.fetch_to_decode_pc[18] ),
    .S(net111),
    .X(_02215_));
 sky130_fd_sc_hd__mux2_1 _13271_ (.A0(\core_pipeline.pipeline_fetch.pc[19] ),
    .A1(\core_pipeline.fetch_to_decode_pc[19] ),
    .S(net112),
    .X(_02216_));
 sky130_fd_sc_hd__mux2_1 _13272_ (.A0(\core_pipeline.pipeline_fetch.pc[20] ),
    .A1(\core_pipeline.fetch_to_decode_pc[20] ),
    .S(net112),
    .X(_02217_));
 sky130_fd_sc_hd__mux2_1 _13273_ (.A0(\core_pipeline.pipeline_fetch.pc[21] ),
    .A1(\core_pipeline.fetch_to_decode_pc[21] ),
    .S(net111),
    .X(_02218_));
 sky130_fd_sc_hd__mux2_1 _13274_ (.A0(\core_pipeline.pipeline_fetch.pc[22] ),
    .A1(\core_pipeline.fetch_to_decode_pc[22] ),
    .S(net111),
    .X(_02219_));
 sky130_fd_sc_hd__mux2_1 _13275_ (.A0(\core_pipeline.pipeline_fetch.pc[23] ),
    .A1(\core_pipeline.fetch_to_decode_pc[23] ),
    .S(net111),
    .X(_02220_));
 sky130_fd_sc_hd__mux2_1 _13276_ (.A0(\core_pipeline.pipeline_fetch.pc[24] ),
    .A1(\core_pipeline.fetch_to_decode_pc[24] ),
    .S(net110),
    .X(_02221_));
 sky130_fd_sc_hd__mux2_1 _13277_ (.A0(\core_pipeline.pipeline_fetch.pc[25] ),
    .A1(\core_pipeline.fetch_to_decode_pc[25] ),
    .S(net110),
    .X(_02222_));
 sky130_fd_sc_hd__mux2_1 _13278_ (.A0(\core_pipeline.pipeline_fetch.pc[26] ),
    .A1(\core_pipeline.fetch_to_decode_pc[26] ),
    .S(net111),
    .X(_02223_));
 sky130_fd_sc_hd__mux2_1 _13279_ (.A0(\core_pipeline.pipeline_fetch.pc[27] ),
    .A1(\core_pipeline.fetch_to_decode_pc[27] ),
    .S(net111),
    .X(_02224_));
 sky130_fd_sc_hd__mux2_1 _13280_ (.A0(\core_pipeline.pipeline_fetch.pc[28] ),
    .A1(\core_pipeline.fetch_to_decode_pc[28] ),
    .S(net111),
    .X(_02225_));
 sky130_fd_sc_hd__mux2_1 _13281_ (.A0(\core_pipeline.pipeline_fetch.pc[29] ),
    .A1(\core_pipeline.fetch_to_decode_pc[29] ),
    .S(net108),
    .X(_02226_));
 sky130_fd_sc_hd__mux2_1 _13282_ (.A0(\core_pipeline.pipeline_fetch.pc[30] ),
    .A1(\core_pipeline.fetch_to_decode_pc[30] ),
    .S(net108),
    .X(_02227_));
 sky130_fd_sc_hd__mux2_1 _13283_ (.A0(\core_pipeline.pipeline_fetch.pc[31] ),
    .A1(\core_pipeline.fetch_to_decode_pc[31] ),
    .S(net109),
    .X(_02228_));
 sky130_fd_sc_hd__mux2_1 _13284_ (.A0(\core_pipeline.pipeline_fetch.pc[0] ),
    .A1(\core_pipeline.fetch_to_decode_next_pc[0] ),
    .S(net107),
    .X(_02229_));
 sky130_fd_sc_hd__mux2_1 _13285_ (.A0(\core_pipeline.pipeline_fetch.pc[1] ),
    .A1(\core_pipeline.fetch_to_decode_next_pc[1] ),
    .S(net109),
    .X(_02230_));
 sky130_fd_sc_hd__mux2_1 _13286_ (.A0(_03312_),
    .A1(\core_pipeline.fetch_to_decode_next_pc[2] ),
    .S(net109),
    .X(_02231_));
 sky130_fd_sc_hd__mux2_1 _13287_ (.A0(_02930_),
    .A1(\core_pipeline.fetch_to_decode_next_pc[3] ),
    .S(net109),
    .X(_02232_));
 sky130_fd_sc_hd__mux2_1 _13288_ (.A0(_02937_),
    .A1(\core_pipeline.fetch_to_decode_next_pc[4] ),
    .S(net112),
    .X(_02233_));
 sky130_fd_sc_hd__mux2_1 _13289_ (.A0(_02944_),
    .A1(\core_pipeline.fetch_to_decode_next_pc[5] ),
    .S(net109),
    .X(_02234_));
 sky130_fd_sc_hd__mux2_1 _13290_ (.A0(_02949_),
    .A1(\core_pipeline.fetch_to_decode_next_pc[6] ),
    .S(net109),
    .X(_02235_));
 sky130_fd_sc_hd__mux2_1 _13291_ (.A0(_02956_),
    .A1(\core_pipeline.fetch_to_decode_next_pc[7] ),
    .S(net109),
    .X(_02236_));
 sky130_fd_sc_hd__mux2_1 _13292_ (.A0(_02963_),
    .A1(\core_pipeline.fetch_to_decode_next_pc[8] ),
    .S(net111),
    .X(_02237_));
 sky130_fd_sc_hd__mux2_1 _13293_ (.A0(_02968_),
    .A1(\core_pipeline.fetch_to_decode_next_pc[9] ),
    .S(net110),
    .X(_02238_));
 sky130_fd_sc_hd__mux2_1 _13294_ (.A0(_02975_),
    .A1(\core_pipeline.fetch_to_decode_next_pc[10] ),
    .S(net110),
    .X(_02239_));
 sky130_fd_sc_hd__mux2_1 _13295_ (.A0(_02982_),
    .A1(\core_pipeline.fetch_to_decode_next_pc[11] ),
    .S(net110),
    .X(_02240_));
 sky130_fd_sc_hd__mux2_1 _13296_ (.A0(_02987_),
    .A1(\core_pipeline.fetch_to_decode_next_pc[12] ),
    .S(net110),
    .X(_02241_));
 sky130_fd_sc_hd__mux2_1 _13297_ (.A0(_02994_),
    .A1(\core_pipeline.fetch_to_decode_next_pc[13] ),
    .S(net110),
    .X(_02242_));
 sky130_fd_sc_hd__mux2_1 _13298_ (.A0(_03001_),
    .A1(\core_pipeline.fetch_to_decode_next_pc[14] ),
    .S(net111),
    .X(_02243_));
 sky130_fd_sc_hd__mux2_1 _13299_ (.A0(_03006_),
    .A1(\core_pipeline.fetch_to_decode_next_pc[15] ),
    .S(net110),
    .X(_02244_));
 sky130_fd_sc_hd__mux2_1 _13300_ (.A0(_03013_),
    .A1(\core_pipeline.fetch_to_decode_next_pc[16] ),
    .S(net110),
    .X(_02245_));
 sky130_fd_sc_hd__mux2_1 _13301_ (.A0(_03020_),
    .A1(\core_pipeline.fetch_to_decode_next_pc[17] ),
    .S(net111),
    .X(_02246_));
 sky130_fd_sc_hd__mux2_1 _13302_ (.A0(_03025_),
    .A1(\core_pipeline.fetch_to_decode_next_pc[18] ),
    .S(net111),
    .X(_02247_));
 sky130_fd_sc_hd__mux2_1 _13303_ (.A0(\core_pipeline.fetch_to_decode_next_pc[19] ),
    .A1(_03032_),
    .S(_03506_),
    .X(_02248_));
 sky130_fd_sc_hd__mux2_1 _13304_ (.A0(\core_pipeline.fetch_to_decode_next_pc[20] ),
    .A1(_03039_),
    .S(_03506_),
    .X(_02249_));
 sky130_fd_sc_hd__mux2_1 _13305_ (.A0(\core_pipeline.fetch_to_decode_next_pc[21] ),
    .A1(_03044_),
    .S(_03506_),
    .X(_02250_));
 sky130_fd_sc_hd__mux2_1 _13306_ (.A0(\core_pipeline.fetch_to_decode_next_pc[22] ),
    .A1(_03051_),
    .S(_03506_),
    .X(_02251_));
 sky130_fd_sc_hd__mux2_1 _13307_ (.A0(\core_pipeline.fetch_to_decode_next_pc[23] ),
    .A1(_03058_),
    .S(_03506_),
    .X(_02252_));
 sky130_fd_sc_hd__mux2_1 _13308_ (.A0(\core_pipeline.fetch_to_decode_next_pc[24] ),
    .A1(_03063_),
    .S(_03506_),
    .X(_02253_));
 sky130_fd_sc_hd__or3_1 _13309_ (.A(net111),
    .B(_03068_),
    .C(_03069_),
    .X(_03310_));
 sky130_fd_sc_hd__a21bo_1 _13310_ (.A1(\core_pipeline.fetch_to_decode_next_pc[25] ),
    .A2(net111),
    .B1_N(_03310_),
    .X(_02254_));
 sky130_fd_sc_hd__mux2_1 _13311_ (.A0(\core_pipeline.fetch_to_decode_next_pc[26] ),
    .A1(_03076_),
    .S(_03506_),
    .X(_02255_));
 sky130_fd_sc_hd__mux2_1 _13312_ (.A0(\core_pipeline.fetch_to_decode_next_pc[27] ),
    .A1(_03081_),
    .S(_03506_),
    .X(_02256_));
 sky130_fd_sc_hd__mux2_1 _13313_ (.A0(\core_pipeline.fetch_to_decode_next_pc[28] ),
    .A1(_03088_),
    .S(_03506_),
    .X(_02257_));
 sky130_fd_sc_hd__mux2_1 _13314_ (.A0(\core_pipeline.fetch_to_decode_next_pc[29] ),
    .A1(_03095_),
    .S(_03506_),
    .X(_02258_));
 sky130_fd_sc_hd__mux2_1 _13315_ (.A0(\core_pipeline.fetch_to_decode_next_pc[30] ),
    .A1(_03101_),
    .S(_03506_),
    .X(_02259_));
 sky130_fd_sc_hd__mux2_1 _13316_ (.A0(\core_pipeline.fetch_to_decode_next_pc[31] ),
    .A1(_03106_),
    .S(_03506_),
    .X(_02260_));
 sky130_fd_sc_hd__a22o_1 _13317_ (.A1(\core_pipeline.memory_to_writeback_ecause[0] ),
    .A2(net458),
    .B1(_05827_),
    .B2(\core_pipeline.execute_to_memory_ecause[0] ),
    .X(_02261_));
 sky130_fd_sc_hd__or4_4 _13318_ (.A(\core_pipeline.memory_to_writeback_rd_address[2] ),
    .B(\core_pipeline.memory_to_writeback_rd_address[3] ),
    .C(_03912_),
    .D(_04934_),
    .X(_03311_));
 sky130_fd_sc_hd__mux2_1 _13319_ (.A0(net349),
    .A1(\core_pipeline.pipeline_registers.registers[18][0] ),
    .S(net163),
    .X(_02262_));
 sky130_fd_sc_hd__mux2_1 _13320_ (.A0(net347),
    .A1(\core_pipeline.pipeline_registers.registers[18][1] ),
    .S(net164),
    .X(_02263_));
 sky130_fd_sc_hd__mux2_1 _13321_ (.A0(net345),
    .A1(\core_pipeline.pipeline_registers.registers[18][2] ),
    .S(net164),
    .X(_02264_));
 sky130_fd_sc_hd__mux2_1 _13322_ (.A0(net343),
    .A1(\core_pipeline.pipeline_registers.registers[18][3] ),
    .S(net163),
    .X(_02265_));
 sky130_fd_sc_hd__mux2_1 _13323_ (.A0(net340),
    .A1(\core_pipeline.pipeline_registers.registers[18][4] ),
    .S(net163),
    .X(_02266_));
 sky130_fd_sc_hd__mux2_1 _13324_ (.A0(net339),
    .A1(\core_pipeline.pipeline_registers.registers[18][5] ),
    .S(net164),
    .X(_02267_));
 sky130_fd_sc_hd__mux2_1 _13325_ (.A0(net336),
    .A1(\core_pipeline.pipeline_registers.registers[18][6] ),
    .S(net164),
    .X(_02268_));
 sky130_fd_sc_hd__mux2_1 _13326_ (.A0(net333),
    .A1(\core_pipeline.pipeline_registers.registers[18][7] ),
    .S(net163),
    .X(_02269_));
 sky130_fd_sc_hd__mux2_1 _13327_ (.A0(net331),
    .A1(\core_pipeline.pipeline_registers.registers[18][8] ),
    .S(net163),
    .X(_02270_));
 sky130_fd_sc_hd__mux2_1 _13328_ (.A0(net330),
    .A1(\core_pipeline.pipeline_registers.registers[18][9] ),
    .S(net163),
    .X(_02271_));
 sky130_fd_sc_hd__mux2_1 _13329_ (.A0(net327),
    .A1(\core_pipeline.pipeline_registers.registers[18][10] ),
    .S(net163),
    .X(_02272_));
 sky130_fd_sc_hd__mux2_1 _13330_ (.A0(net325),
    .A1(\core_pipeline.pipeline_registers.registers[18][11] ),
    .S(net163),
    .X(_02273_));
 sky130_fd_sc_hd__mux2_1 _13331_ (.A0(net323),
    .A1(\core_pipeline.pipeline_registers.registers[18][12] ),
    .S(net163),
    .X(_02274_));
 sky130_fd_sc_hd__mux2_1 _13332_ (.A0(net321),
    .A1(\core_pipeline.pipeline_registers.registers[18][13] ),
    .S(net163),
    .X(_02275_));
 sky130_fd_sc_hd__mux2_1 _13333_ (.A0(net319),
    .A1(\core_pipeline.pipeline_registers.registers[18][14] ),
    .S(net163),
    .X(_02276_));
 sky130_fd_sc_hd__mux2_1 _13334_ (.A0(net317),
    .A1(\core_pipeline.pipeline_registers.registers[18][15] ),
    .S(net163),
    .X(_02277_));
 sky130_fd_sc_hd__mux2_1 _13335_ (.A0(net316),
    .A1(\core_pipeline.pipeline_registers.registers[18][16] ),
    .S(net163),
    .X(_02278_));
 sky130_fd_sc_hd__mux2_1 _13336_ (.A0(net313),
    .A1(\core_pipeline.pipeline_registers.registers[18][17] ),
    .S(net164),
    .X(_02279_));
 sky130_fd_sc_hd__mux2_1 _13337_ (.A0(net310),
    .A1(\core_pipeline.pipeline_registers.registers[18][18] ),
    .S(net164),
    .X(_02280_));
 sky130_fd_sc_hd__mux2_1 _13338_ (.A0(net309),
    .A1(\core_pipeline.pipeline_registers.registers[18][19] ),
    .S(net164),
    .X(_02281_));
 sky130_fd_sc_hd__mux2_1 _13339_ (.A0(net306),
    .A1(\core_pipeline.pipeline_registers.registers[18][20] ),
    .S(net164),
    .X(_02282_));
 sky130_fd_sc_hd__mux2_1 _13340_ (.A0(net304),
    .A1(\core_pipeline.pipeline_registers.registers[18][21] ),
    .S(net164),
    .X(_02283_));
 sky130_fd_sc_hd__mux2_1 _13341_ (.A0(net302),
    .A1(\core_pipeline.pipeline_registers.registers[18][22] ),
    .S(net163),
    .X(_02284_));
 sky130_fd_sc_hd__mux2_1 _13342_ (.A0(net299),
    .A1(\core_pipeline.pipeline_registers.registers[18][23] ),
    .S(net164),
    .X(_02285_));
 sky130_fd_sc_hd__mux2_1 _13343_ (.A0(net298),
    .A1(\core_pipeline.pipeline_registers.registers[18][24] ),
    .S(net163),
    .X(_02286_));
 sky130_fd_sc_hd__mux2_1 _13344_ (.A0(net296),
    .A1(\core_pipeline.pipeline_registers.registers[18][25] ),
    .S(net163),
    .X(_02287_));
 sky130_fd_sc_hd__mux2_1 _13345_ (.A0(net293),
    .A1(\core_pipeline.pipeline_registers.registers[18][26] ),
    .S(net163),
    .X(_02288_));
 sky130_fd_sc_hd__mux2_1 _13346_ (.A0(net291),
    .A1(\core_pipeline.pipeline_registers.registers[18][27] ),
    .S(net164),
    .X(_02289_));
 sky130_fd_sc_hd__mux2_1 _13347_ (.A0(net290),
    .A1(\core_pipeline.pipeline_registers.registers[18][28] ),
    .S(net164),
    .X(_02290_));
 sky130_fd_sc_hd__mux2_1 _13348_ (.A0(net287),
    .A1(\core_pipeline.pipeline_registers.registers[18][29] ),
    .S(net164),
    .X(_02291_));
 sky130_fd_sc_hd__mux2_1 _13349_ (.A0(net285),
    .A1(\core_pipeline.pipeline_registers.registers[18][30] ),
    .S(net164),
    .X(_02292_));
 sky130_fd_sc_hd__mux2_1 _13350_ (.A0(net282),
    .A1(\core_pipeline.pipeline_registers.registers[18][31] ),
    .S(net164),
    .X(_02293_));
 sky130_fd_sc_hd__clkbuf_2 _13351_ (.A(\core_pipeline.pipeline_registers.registers[0][0] ),
    .X(_01079_));
 sky130_fd_sc_hd__clkbuf_2 _13352_ (.A(\core_pipeline.pipeline_registers.registers[0][1] ),
    .X(_01080_));
 sky130_fd_sc_hd__clkbuf_2 _13353_ (.A(\core_pipeline.pipeline_registers.registers[0][2] ),
    .X(_01081_));
 sky130_fd_sc_hd__clkbuf_2 _13354_ (.A(\core_pipeline.pipeline_registers.registers[0][3] ),
    .X(_01082_));
 sky130_fd_sc_hd__clkbuf_2 _13355_ (.A(\core_pipeline.pipeline_registers.registers[0][4] ),
    .X(_01083_));
 sky130_fd_sc_hd__clkbuf_2 _13356_ (.A(\core_pipeline.pipeline_registers.registers[0][5] ),
    .X(_01084_));
 sky130_fd_sc_hd__clkbuf_2 _13357_ (.A(\core_pipeline.pipeline_registers.registers[0][6] ),
    .X(_01085_));
 sky130_fd_sc_hd__clkbuf_2 _13358_ (.A(\core_pipeline.pipeline_registers.registers[0][7] ),
    .X(_01086_));
 sky130_fd_sc_hd__clkbuf_2 _13359_ (.A(\core_pipeline.pipeline_registers.registers[0][8] ),
    .X(_01087_));
 sky130_fd_sc_hd__clkbuf_2 _13360_ (.A(\core_pipeline.pipeline_registers.registers[0][9] ),
    .X(_01088_));
 sky130_fd_sc_hd__clkbuf_2 _13361_ (.A(\core_pipeline.pipeline_registers.registers[0][10] ),
    .X(_01089_));
 sky130_fd_sc_hd__clkbuf_2 _13362_ (.A(\core_pipeline.pipeline_registers.registers[0][11] ),
    .X(_01090_));
 sky130_fd_sc_hd__clkbuf_2 _13363_ (.A(\core_pipeline.pipeline_registers.registers[0][12] ),
    .X(_01091_));
 sky130_fd_sc_hd__clkbuf_2 _13364_ (.A(\core_pipeline.pipeline_registers.registers[0][13] ),
    .X(_01092_));
 sky130_fd_sc_hd__clkbuf_2 _13365_ (.A(\core_pipeline.pipeline_registers.registers[0][14] ),
    .X(_01093_));
 sky130_fd_sc_hd__clkbuf_2 _13366_ (.A(\core_pipeline.pipeline_registers.registers[0][15] ),
    .X(_01094_));
 sky130_fd_sc_hd__clkbuf_2 _13367_ (.A(\core_pipeline.pipeline_registers.registers[0][16] ),
    .X(_01095_));
 sky130_fd_sc_hd__clkbuf_2 _13368_ (.A(\core_pipeline.pipeline_registers.registers[0][17] ),
    .X(_01096_));
 sky130_fd_sc_hd__clkbuf_2 _13369_ (.A(\core_pipeline.pipeline_registers.registers[0][18] ),
    .X(_01097_));
 sky130_fd_sc_hd__clkbuf_2 _13370_ (.A(\core_pipeline.pipeline_registers.registers[0][19] ),
    .X(_01098_));
 sky130_fd_sc_hd__clkbuf_2 _13371_ (.A(\core_pipeline.pipeline_registers.registers[0][20] ),
    .X(_01099_));
 sky130_fd_sc_hd__clkbuf_2 _13372_ (.A(\core_pipeline.pipeline_registers.registers[0][21] ),
    .X(_01100_));
 sky130_fd_sc_hd__clkbuf_2 _13373_ (.A(\core_pipeline.pipeline_registers.registers[0][22] ),
    .X(_01101_));
 sky130_fd_sc_hd__clkbuf_2 _13374_ (.A(\core_pipeline.pipeline_registers.registers[0][23] ),
    .X(_01102_));
 sky130_fd_sc_hd__clkbuf_2 _13375_ (.A(\core_pipeline.pipeline_registers.registers[0][24] ),
    .X(_01103_));
 sky130_fd_sc_hd__clkbuf_2 _13376_ (.A(\core_pipeline.pipeline_registers.registers[0][25] ),
    .X(_01104_));
 sky130_fd_sc_hd__clkbuf_2 _13377_ (.A(\core_pipeline.pipeline_registers.registers[0][26] ),
    .X(_01105_));
 sky130_fd_sc_hd__clkbuf_2 _13378_ (.A(\core_pipeline.pipeline_registers.registers[0][27] ),
    .X(_01106_));
 sky130_fd_sc_hd__clkbuf_2 _13379_ (.A(\core_pipeline.pipeline_registers.registers[0][28] ),
    .X(_01107_));
 sky130_fd_sc_hd__clkbuf_2 _13380_ (.A(\core_pipeline.pipeline_registers.registers[0][29] ),
    .X(_01108_));
 sky130_fd_sc_hd__clkbuf_2 _13381_ (.A(\core_pipeline.pipeline_registers.registers[0][30] ),
    .X(_01109_));
 sky130_fd_sc_hd__clkbuf_2 _13382_ (.A(\core_pipeline.pipeline_registers.registers[0][31] ),
    .X(_01110_));
 sky130_fd_sc_hd__dfxtp_1 _13383_ (.CLK(clknet_leaf_250_clk),
    .D(_00041_),
    .Q(\core_pipeline.pipeline_registers.registers[19][0] ));
 sky130_fd_sc_hd__dfxtp_1 _13384_ (.CLK(clknet_leaf_161_clk),
    .D(_00042_),
    .Q(\core_pipeline.pipeline_registers.registers[19][1] ));
 sky130_fd_sc_hd__dfxtp_1 _13385_ (.CLK(clknet_leaf_197_clk),
    .D(_00043_),
    .Q(\core_pipeline.pipeline_registers.registers[19][2] ));
 sky130_fd_sc_hd__dfxtp_1 _13386_ (.CLK(clknet_leaf_235_clk),
    .D(_00044_),
    .Q(\core_pipeline.pipeline_registers.registers[19][3] ));
 sky130_fd_sc_hd__dfxtp_1 _13387_ (.CLK(clknet_leaf_5_clk),
    .D(_00045_),
    .Q(\core_pipeline.pipeline_registers.registers[19][4] ));
 sky130_fd_sc_hd__dfxtp_1 _13388_ (.CLK(clknet_leaf_198_clk),
    .D(_00046_),
    .Q(\core_pipeline.pipeline_registers.registers[19][5] ));
 sky130_fd_sc_hd__dfxtp_1 _13389_ (.CLK(clknet_leaf_206_clk),
    .D(_00047_),
    .Q(\core_pipeline.pipeline_registers.registers[19][6] ));
 sky130_fd_sc_hd__dfxtp_1 _13390_ (.CLK(clknet_leaf_232_clk),
    .D(_00048_),
    .Q(\core_pipeline.pipeline_registers.registers[19][7] ));
 sky130_fd_sc_hd__dfxtp_1 _13391_ (.CLK(clknet_leaf_242_clk),
    .D(_00049_),
    .Q(\core_pipeline.pipeline_registers.registers[19][8] ));
 sky130_fd_sc_hd__dfxtp_1 _13392_ (.CLK(clknet_leaf_6_clk),
    .D(_00050_),
    .Q(\core_pipeline.pipeline_registers.registers[19][9] ));
 sky130_fd_sc_hd__dfxtp_1 _13393_ (.CLK(clknet_leaf_10_clk),
    .D(_00051_),
    .Q(\core_pipeline.pipeline_registers.registers[19][10] ));
 sky130_fd_sc_hd__dfxtp_1 _13394_ (.CLK(clknet_leaf_5_clk),
    .D(_00052_),
    .Q(\core_pipeline.pipeline_registers.registers[19][11] ));
 sky130_fd_sc_hd__dfxtp_1 _13395_ (.CLK(clknet_leaf_25_clk),
    .D(_00053_),
    .Q(\core_pipeline.pipeline_registers.registers[19][12] ));
 sky130_fd_sc_hd__dfxtp_1 _13396_ (.CLK(clknet_leaf_9_clk),
    .D(_00054_),
    .Q(\core_pipeline.pipeline_registers.registers[19][13] ));
 sky130_fd_sc_hd__dfxtp_1 _13397_ (.CLK(clknet_leaf_4_clk),
    .D(_00055_),
    .Q(\core_pipeline.pipeline_registers.registers[19][14] ));
 sky130_fd_sc_hd__dfxtp_1 _13398_ (.CLK(clknet_leaf_20_clk),
    .D(_00056_),
    .Q(\core_pipeline.pipeline_registers.registers[19][15] ));
 sky130_fd_sc_hd__dfxtp_1 _13399_ (.CLK(clknet_leaf_245_clk),
    .D(_00057_),
    .Q(\core_pipeline.pipeline_registers.registers[19][16] ));
 sky130_fd_sc_hd__dfxtp_1 _13400_ (.CLK(clknet_leaf_213_clk),
    .D(_00058_),
    .Q(\core_pipeline.pipeline_registers.registers[19][17] ));
 sky130_fd_sc_hd__dfxtp_1 _13401_ (.CLK(clknet_leaf_179_clk),
    .D(_00059_),
    .Q(\core_pipeline.pipeline_registers.registers[19][18] ));
 sky130_fd_sc_hd__dfxtp_1 _13402_ (.CLK(clknet_leaf_195_clk),
    .D(_00060_),
    .Q(\core_pipeline.pipeline_registers.registers[19][19] ));
 sky130_fd_sc_hd__dfxtp_1 _13403_ (.CLK(clknet_leaf_183_clk),
    .D(_00061_),
    .Q(\core_pipeline.pipeline_registers.registers[19][20] ));
 sky130_fd_sc_hd__dfxtp_1 _13404_ (.CLK(clknet_leaf_168_clk),
    .D(_00062_),
    .Q(\core_pipeline.pipeline_registers.registers[19][21] ));
 sky130_fd_sc_hd__dfxtp_1 _13405_ (.CLK(clknet_leaf_211_clk),
    .D(_00063_),
    .Q(\core_pipeline.pipeline_registers.registers[19][22] ));
 sky130_fd_sc_hd__dfxtp_1 _13406_ (.CLK(clknet_leaf_209_clk),
    .D(_00064_),
    .Q(\core_pipeline.pipeline_registers.registers[19][23] ));
 sky130_fd_sc_hd__dfxtp_1 _13407_ (.CLK(clknet_leaf_224_clk),
    .D(_00065_),
    .Q(\core_pipeline.pipeline_registers.registers[19][24] ));
 sky130_fd_sc_hd__dfxtp_1 _13408_ (.CLK(clknet_leaf_10_clk),
    .D(_00066_),
    .Q(\core_pipeline.pipeline_registers.registers[19][25] ));
 sky130_fd_sc_hd__dfxtp_1 _13409_ (.CLK(clknet_leaf_18_clk),
    .D(_00067_),
    .Q(\core_pipeline.pipeline_registers.registers[19][26] ));
 sky130_fd_sc_hd__dfxtp_1 _13410_ (.CLK(clknet_leaf_166_clk),
    .D(_00068_),
    .Q(\core_pipeline.pipeline_registers.registers[19][27] ));
 sky130_fd_sc_hd__dfxtp_1 _13411_ (.CLK(clknet_leaf_182_clk),
    .D(_00069_),
    .Q(\core_pipeline.pipeline_registers.registers[19][28] ));
 sky130_fd_sc_hd__dfxtp_1 _13412_ (.CLK(clknet_leaf_210_clk),
    .D(_00070_),
    .Q(\core_pipeline.pipeline_registers.registers[19][29] ));
 sky130_fd_sc_hd__dfxtp_1 _13413_ (.CLK(clknet_leaf_210_clk),
    .D(_00071_),
    .Q(\core_pipeline.pipeline_registers.registers[19][30] ));
 sky130_fd_sc_hd__dfxtp_1 _13414_ (.CLK(clknet_leaf_176_clk),
    .D(_00072_),
    .Q(\core_pipeline.pipeline_registers.registers[19][31] ));
 sky130_fd_sc_hd__dfxtp_1 _13415_ (.CLK(clknet_leaf_148_clk),
    .D(_00073_),
    .Q(\core_pipeline.csr_to_fetch_trap_vector[2] ));
 sky130_fd_sc_hd__dfxtp_1 _13416_ (.CLK(clknet_leaf_147_clk),
    .D(_00074_),
    .Q(\core_pipeline.csr_to_fetch_trap_vector[3] ));
 sky130_fd_sc_hd__dfxtp_2 _13417_ (.CLK(clknet_leaf_148_clk),
    .D(_00075_),
    .Q(\core_pipeline.csr_to_fetch_trap_vector[4] ));
 sky130_fd_sc_hd__dfxtp_1 _13418_ (.CLK(clknet_leaf_145_clk),
    .D(_00076_),
    .Q(\core_pipeline.csr_to_fetch_trap_vector[5] ));
 sky130_fd_sc_hd__dfxtp_2 _13419_ (.CLK(clknet_leaf_144_clk),
    .D(_00077_),
    .Q(\core_pipeline.csr_to_fetch_trap_vector[6] ));
 sky130_fd_sc_hd__dfxtp_1 _13420_ (.CLK(clknet_leaf_145_clk),
    .D(_00078_),
    .Q(\core_pipeline.csr_to_fetch_trap_vector[7] ));
 sky130_fd_sc_hd__dfxtp_1 _13421_ (.CLK(clknet_leaf_100_clk),
    .D(_00079_),
    .Q(\core_pipeline.csr_to_fetch_trap_vector[8] ));
 sky130_fd_sc_hd__dfxtp_2 _13422_ (.CLK(clknet_leaf_114_clk),
    .D(_00080_),
    .Q(\core_pipeline.csr_to_fetch_trap_vector[9] ));
 sky130_fd_sc_hd__dfxtp_2 _13423_ (.CLK(clknet_leaf_114_clk),
    .D(_00081_),
    .Q(\core_pipeline.csr_to_fetch_trap_vector[10] ));
 sky130_fd_sc_hd__dfxtp_4 _13424_ (.CLK(clknet_leaf_114_clk),
    .D(_00082_),
    .Q(\core_pipeline.csr_to_fetch_trap_vector[11] ));
 sky130_fd_sc_hd__dfxtp_1 _13425_ (.CLK(clknet_leaf_111_clk),
    .D(_00083_),
    .Q(\core_pipeline.csr_to_fetch_trap_vector[12] ));
 sky130_fd_sc_hd__dfxtp_1 _13426_ (.CLK(clknet_leaf_113_clk),
    .D(_00084_),
    .Q(\core_pipeline.csr_to_fetch_trap_vector[13] ));
 sky130_fd_sc_hd__dfxtp_2 _13427_ (.CLK(clknet_leaf_113_clk),
    .D(_00085_),
    .Q(\core_pipeline.csr_to_fetch_trap_vector[14] ));
 sky130_fd_sc_hd__dfxtp_2 _13428_ (.CLK(clknet_leaf_113_clk),
    .D(_00086_),
    .Q(\core_pipeline.csr_to_fetch_trap_vector[15] ));
 sky130_fd_sc_hd__dfxtp_2 _13429_ (.CLK(clknet_leaf_113_clk),
    .D(_00087_),
    .Q(\core_pipeline.csr_to_fetch_trap_vector[16] ));
 sky130_fd_sc_hd__dfxtp_2 _13430_ (.CLK(clknet_leaf_113_clk),
    .D(_00088_),
    .Q(\core_pipeline.csr_to_fetch_trap_vector[17] ));
 sky130_fd_sc_hd__dfxtp_2 _13431_ (.CLK(clknet_leaf_121_clk),
    .D(_00089_),
    .Q(\core_pipeline.csr_to_fetch_trap_vector[18] ));
 sky130_fd_sc_hd__dfxtp_2 _13432_ (.CLK(clknet_leaf_120_clk),
    .D(_00090_),
    .Q(\core_pipeline.csr_to_fetch_trap_vector[19] ));
 sky130_fd_sc_hd__dfxtp_1 _13433_ (.CLK(clknet_leaf_120_clk),
    .D(_00091_),
    .Q(\core_pipeline.csr_to_fetch_trap_vector[20] ));
 sky130_fd_sc_hd__dfxtp_1 _13434_ (.CLK(clknet_leaf_119_clk),
    .D(_00092_),
    .Q(\core_pipeline.csr_to_fetch_trap_vector[21] ));
 sky130_fd_sc_hd__dfxtp_1 _13435_ (.CLK(clknet_leaf_130_clk),
    .D(_00093_),
    .Q(\core_pipeline.csr_to_fetch_trap_vector[22] ));
 sky130_fd_sc_hd__dfxtp_1 _13436_ (.CLK(clknet_leaf_130_clk),
    .D(_00094_),
    .Q(\core_pipeline.csr_to_fetch_trap_vector[23] ));
 sky130_fd_sc_hd__dfxtp_1 _13437_ (.CLK(clknet_leaf_130_clk),
    .D(_00095_),
    .Q(\core_pipeline.csr_to_fetch_trap_vector[24] ));
 sky130_fd_sc_hd__dfxtp_1 _13438_ (.CLK(clknet_leaf_130_clk),
    .D(_00096_),
    .Q(\core_pipeline.csr_to_fetch_trap_vector[25] ));
 sky130_fd_sc_hd__dfxtp_1 _13439_ (.CLK(clknet_leaf_100_clk),
    .D(_00097_),
    .Q(\core_pipeline.csr_to_fetch_trap_vector[26] ));
 sky130_fd_sc_hd__dfxtp_1 _13440_ (.CLK(clknet_leaf_130_clk),
    .D(_00098_),
    .Q(\core_pipeline.csr_to_fetch_trap_vector[27] ));
 sky130_fd_sc_hd__dfxtp_1 _13441_ (.CLK(clknet_leaf_145_clk),
    .D(_00099_),
    .Q(\core_pipeline.csr_to_fetch_trap_vector[28] ));
 sky130_fd_sc_hd__dfxtp_2 _13442_ (.CLK(clknet_leaf_145_clk),
    .D(_00100_),
    .Q(\core_pipeline.csr_to_fetch_trap_vector[29] ));
 sky130_fd_sc_hd__dfxtp_1 _13443_ (.CLK(clknet_leaf_146_clk),
    .D(_00101_),
    .Q(\core_pipeline.csr_to_fetch_trap_vector[30] ));
 sky130_fd_sc_hd__dfxtp_2 _13444_ (.CLK(clknet_leaf_146_clk),
    .D(_00102_),
    .Q(\core_pipeline.csr_to_fetch_trap_vector[31] ));
 sky130_fd_sc_hd__dfxtp_2 _13445_ (.CLK(clknet_leaf_140_clk),
    .D(_00103_),
    .Q(\core_pipeline.pipeline_csr.cycle[0] ));
 sky130_fd_sc_hd__dfxtp_2 _13446_ (.CLK(clknet_leaf_140_clk),
    .D(_00104_),
    .Q(\core_pipeline.pipeline_csr.cycle[1] ));
 sky130_fd_sc_hd__dfxtp_1 _13447_ (.CLK(clknet_leaf_142_clk),
    .D(_00105_),
    .Q(\core_pipeline.pipeline_csr.cycle[2] ));
 sky130_fd_sc_hd__dfxtp_2 _13448_ (.CLK(clknet_leaf_142_clk),
    .D(_00106_),
    .Q(\core_pipeline.pipeline_csr.cycle[3] ));
 sky130_fd_sc_hd__dfxtp_2 _13449_ (.CLK(clknet_leaf_143_clk),
    .D(_00107_),
    .Q(\core_pipeline.pipeline_csr.cycle[4] ));
 sky130_fd_sc_hd__dfxtp_2 _13450_ (.CLK(clknet_leaf_143_clk),
    .D(_00108_),
    .Q(\core_pipeline.pipeline_csr.cycle[5] ));
 sky130_fd_sc_hd__dfxtp_2 _13451_ (.CLK(clknet_leaf_144_clk),
    .D(_00109_),
    .Q(\core_pipeline.pipeline_csr.cycle[6] ));
 sky130_fd_sc_hd__dfxtp_2 _13452_ (.CLK(clknet_leaf_100_clk),
    .D(_00110_),
    .Q(\core_pipeline.pipeline_csr.cycle[7] ));
 sky130_fd_sc_hd__dfxtp_1 _13453_ (.CLK(clknet_leaf_118_clk),
    .D(_00111_),
    .Q(\core_pipeline.pipeline_csr.cycle[8] ));
 sky130_fd_sc_hd__dfxtp_1 _13454_ (.CLK(clknet_leaf_118_clk),
    .D(_00112_),
    .Q(\core_pipeline.pipeline_csr.cycle[9] ));
 sky130_fd_sc_hd__dfxtp_1 _13455_ (.CLK(clknet_leaf_118_clk),
    .D(_00113_),
    .Q(\core_pipeline.pipeline_csr.cycle[10] ));
 sky130_fd_sc_hd__dfxtp_2 _13456_ (.CLK(clknet_leaf_114_clk),
    .D(_00114_),
    .Q(\core_pipeline.pipeline_csr.cycle[11] ));
 sky130_fd_sc_hd__dfxtp_1 _13457_ (.CLK(clknet_leaf_113_clk),
    .D(_00115_),
    .Q(\core_pipeline.pipeline_csr.cycle[12] ));
 sky130_fd_sc_hd__dfxtp_2 _13458_ (.CLK(clknet_leaf_113_clk),
    .D(_00116_),
    .Q(\core_pipeline.pipeline_csr.cycle[13] ));
 sky130_fd_sc_hd__dfxtp_2 _13459_ (.CLK(clknet_leaf_113_clk),
    .D(_00117_),
    .Q(\core_pipeline.pipeline_csr.cycle[14] ));
 sky130_fd_sc_hd__dfxtp_1 _13460_ (.CLK(clknet_leaf_121_clk),
    .D(_00118_),
    .Q(\core_pipeline.pipeline_csr.cycle[15] ));
 sky130_fd_sc_hd__dfxtp_2 _13461_ (.CLK(clknet_leaf_122_clk),
    .D(_00119_),
    .Q(\core_pipeline.pipeline_csr.cycle[16] ));
 sky130_fd_sc_hd__dfxtp_2 _13462_ (.CLK(clknet_leaf_123_clk),
    .D(_00120_),
    .Q(\core_pipeline.pipeline_csr.cycle[17] ));
 sky130_fd_sc_hd__dfxtp_2 _13463_ (.CLK(clknet_leaf_123_clk),
    .D(_00121_),
    .Q(\core_pipeline.pipeline_csr.cycle[18] ));
 sky130_fd_sc_hd__dfxtp_1 _13464_ (.CLK(clknet_leaf_123_clk),
    .D(_00122_),
    .Q(\core_pipeline.pipeline_csr.cycle[19] ));
 sky130_fd_sc_hd__dfxtp_2 _13465_ (.CLK(clknet_leaf_123_clk),
    .D(_00123_),
    .Q(\core_pipeline.pipeline_csr.cycle[20] ));
 sky130_fd_sc_hd__dfxtp_2 _13466_ (.CLK(clknet_leaf_120_clk),
    .D(_00124_),
    .Q(\core_pipeline.pipeline_csr.cycle[21] ));
 sky130_fd_sc_hd__dfxtp_1 _13467_ (.CLK(clknet_leaf_129_clk),
    .D(_00125_),
    .Q(\core_pipeline.pipeline_csr.cycle[22] ));
 sky130_fd_sc_hd__dfxtp_1 _13468_ (.CLK(clknet_leaf_129_clk),
    .D(_00126_),
    .Q(\core_pipeline.pipeline_csr.cycle[23] ));
 sky130_fd_sc_hd__dfxtp_4 _13469_ (.CLK(clknet_leaf_129_clk),
    .D(_00127_),
    .Q(\core_pipeline.pipeline_csr.cycle[24] ));
 sky130_fd_sc_hd__dfxtp_2 _13470_ (.CLK(clknet_leaf_130_clk),
    .D(_00128_),
    .Q(\core_pipeline.pipeline_csr.cycle[25] ));
 sky130_fd_sc_hd__dfxtp_2 _13471_ (.CLK(clknet_leaf_134_clk),
    .D(_00129_),
    .Q(\core_pipeline.pipeline_csr.cycle[26] ));
 sky130_fd_sc_hd__dfxtp_1 _13472_ (.CLK(clknet_leaf_134_clk),
    .D(_00130_),
    .Q(\core_pipeline.pipeline_csr.cycle[27] ));
 sky130_fd_sc_hd__dfxtp_2 _13473_ (.CLK(clknet_leaf_133_clk),
    .D(_00131_),
    .Q(\core_pipeline.pipeline_csr.cycle[28] ));
 sky130_fd_sc_hd__dfxtp_2 _13474_ (.CLK(clknet_leaf_133_clk),
    .D(_00132_),
    .Q(\core_pipeline.pipeline_csr.cycle[29] ));
 sky130_fd_sc_hd__dfxtp_2 _13475_ (.CLK(clknet_leaf_133_clk),
    .D(_00133_),
    .Q(\core_pipeline.pipeline_csr.cycle[30] ));
 sky130_fd_sc_hd__dfxtp_2 _13476_ (.CLK(clknet_leaf_137_clk),
    .D(_00134_),
    .Q(\core_pipeline.pipeline_csr.cycle[31] ));
 sky130_fd_sc_hd__dfxtp_2 _13477_ (.CLK(clknet_leaf_139_clk),
    .D(_00135_),
    .Q(\core_pipeline.pipeline_csr.cycle[32] ));
 sky130_fd_sc_hd__dfxtp_4 _13478_ (.CLK(clknet_leaf_139_clk),
    .D(_00136_),
    .Q(\core_pipeline.pipeline_csr.cycle[33] ));
 sky130_fd_sc_hd__dfxtp_4 _13479_ (.CLK(clknet_leaf_137_clk),
    .D(_00137_),
    .Q(\core_pipeline.pipeline_csr.cycle[34] ));
 sky130_fd_sc_hd__dfxtp_2 _13480_ (.CLK(clknet_leaf_140_clk),
    .D(_00138_),
    .Q(\core_pipeline.pipeline_csr.cycle[35] ));
 sky130_fd_sc_hd__dfxtp_2 _13481_ (.CLK(clknet_leaf_143_clk),
    .D(_00139_),
    .Q(\core_pipeline.pipeline_csr.cycle[36] ));
 sky130_fd_sc_hd__dfxtp_2 _13482_ (.CLK(clknet_leaf_143_clk),
    .D(_00140_),
    .Q(\core_pipeline.pipeline_csr.cycle[37] ));
 sky130_fd_sc_hd__dfxtp_2 _13483_ (.CLK(clknet_leaf_132_clk),
    .D(_00141_),
    .Q(\core_pipeline.pipeline_csr.cycle[38] ));
 sky130_fd_sc_hd__dfxtp_2 _13484_ (.CLK(clknet_leaf_131_clk),
    .D(_00142_),
    .Q(\core_pipeline.pipeline_csr.cycle[39] ));
 sky130_fd_sc_hd__dfxtp_2 _13485_ (.CLK(clknet_leaf_130_clk),
    .D(_00143_),
    .Q(\core_pipeline.pipeline_csr.cycle[40] ));
 sky130_fd_sc_hd__dfxtp_2 _13486_ (.CLK(clknet_leaf_119_clk),
    .D(_00144_),
    .Q(\core_pipeline.pipeline_csr.cycle[41] ));
 sky130_fd_sc_hd__dfxtp_2 _13487_ (.CLK(clknet_leaf_118_clk),
    .D(_00145_),
    .Q(\core_pipeline.pipeline_csr.cycle[42] ));
 sky130_fd_sc_hd__dfxtp_4 _13488_ (.CLK(clknet_leaf_119_clk),
    .D(_00146_),
    .Q(\core_pipeline.pipeline_csr.cycle[43] ));
 sky130_fd_sc_hd__dfxtp_4 _13489_ (.CLK(clknet_leaf_121_clk),
    .D(_00147_),
    .Q(\core_pipeline.pipeline_csr.cycle[44] ));
 sky130_fd_sc_hd__dfxtp_2 _13490_ (.CLK(clknet_leaf_121_clk),
    .D(_00148_),
    .Q(\core_pipeline.pipeline_csr.cycle[45] ));
 sky130_fd_sc_hd__dfxtp_2 _13491_ (.CLK(clknet_leaf_121_clk),
    .D(_00149_),
    .Q(\core_pipeline.pipeline_csr.cycle[46] ));
 sky130_fd_sc_hd__dfxtp_2 _13492_ (.CLK(clknet_leaf_120_clk),
    .D(_00150_),
    .Q(\core_pipeline.pipeline_csr.cycle[47] ));
 sky130_fd_sc_hd__dfxtp_2 _13493_ (.CLK(clknet_leaf_123_clk),
    .D(_00151_),
    .Q(\core_pipeline.pipeline_csr.cycle[48] ));
 sky130_fd_sc_hd__dfxtp_2 _13494_ (.CLK(clknet_leaf_125_clk),
    .D(_00152_),
    .Q(\core_pipeline.pipeline_csr.cycle[49] ));
 sky130_fd_sc_hd__dfxtp_2 _13495_ (.CLK(clknet_leaf_125_clk),
    .D(_00153_),
    .Q(\core_pipeline.pipeline_csr.cycle[50] ));
 sky130_fd_sc_hd__dfxtp_1 _13496_ (.CLK(clknet_leaf_125_clk),
    .D(_00154_),
    .Q(\core_pipeline.pipeline_csr.cycle[51] ));
 sky130_fd_sc_hd__dfxtp_2 _13497_ (.CLK(clknet_leaf_125_clk),
    .D(_00155_),
    .Q(\core_pipeline.pipeline_csr.cycle[52] ));
 sky130_fd_sc_hd__dfxtp_2 _13498_ (.CLK(clknet_leaf_127_clk),
    .D(_00156_),
    .Q(\core_pipeline.pipeline_csr.cycle[53] ));
 sky130_fd_sc_hd__dfxtp_2 _13499_ (.CLK(clknet_leaf_127_clk),
    .D(_00157_),
    .Q(\core_pipeline.pipeline_csr.cycle[54] ));
 sky130_fd_sc_hd__dfxtp_1 _13500_ (.CLK(clknet_leaf_127_clk),
    .D(_00158_),
    .Q(\core_pipeline.pipeline_csr.cycle[55] ));
 sky130_fd_sc_hd__dfxtp_2 _13501_ (.CLK(clknet_leaf_127_clk),
    .D(_00159_),
    .Q(\core_pipeline.pipeline_csr.cycle[56] ));
 sky130_fd_sc_hd__dfxtp_2 _13502_ (.CLK(clknet_leaf_128_clk),
    .D(_00160_),
    .Q(\core_pipeline.pipeline_csr.cycle[57] ));
 sky130_fd_sc_hd__dfxtp_2 _13503_ (.CLK(clknet_leaf_134_clk),
    .D(_00161_),
    .Q(\core_pipeline.pipeline_csr.cycle[58] ));
 sky130_fd_sc_hd__dfxtp_2 _13504_ (.CLK(clknet_leaf_134_clk),
    .D(_00162_),
    .Q(\core_pipeline.pipeline_csr.cycle[59] ));
 sky130_fd_sc_hd__dfxtp_1 _13505_ (.CLK(clknet_leaf_134_clk),
    .D(_00163_),
    .Q(\core_pipeline.pipeline_csr.cycle[60] ));
 sky130_fd_sc_hd__dfxtp_2 _13506_ (.CLK(clknet_leaf_135_clk),
    .D(_00164_),
    .Q(\core_pipeline.pipeline_csr.cycle[61] ));
 sky130_fd_sc_hd__dfxtp_2 _13507_ (.CLK(clknet_leaf_136_clk),
    .D(_00165_),
    .Q(\core_pipeline.pipeline_csr.cycle[62] ));
 sky130_fd_sc_hd__dfxtp_1 _13508_ (.CLK(clknet_leaf_136_clk),
    .D(_00166_),
    .Q(\core_pipeline.pipeline_csr.cycle[63] ));
 sky130_fd_sc_hd__dfxtp_1 _13509_ (.CLK(clknet_leaf_149_clk),
    .D(_00167_),
    .Q(\core_pipeline.pipeline_csr.instret[0] ));
 sky130_fd_sc_hd__dfxtp_1 _13510_ (.CLK(clknet_leaf_142_clk),
    .D(_00168_),
    .Q(\core_pipeline.pipeline_csr.instret[1] ));
 sky130_fd_sc_hd__dfxtp_2 _13511_ (.CLK(clknet_leaf_142_clk),
    .D(_00169_),
    .Q(\core_pipeline.pipeline_csr.instret[2] ));
 sky130_fd_sc_hd__dfxtp_1 _13512_ (.CLK(clknet_leaf_142_clk),
    .D(_00170_),
    .Q(\core_pipeline.pipeline_csr.instret[3] ));
 sky130_fd_sc_hd__dfxtp_1 _13513_ (.CLK(clknet_leaf_146_clk),
    .D(_00171_),
    .Q(\core_pipeline.pipeline_csr.instret[4] ));
 sky130_fd_sc_hd__dfxtp_1 _13514_ (.CLK(clknet_leaf_144_clk),
    .D(_00172_),
    .Q(\core_pipeline.pipeline_csr.instret[5] ));
 sky130_fd_sc_hd__dfxtp_1 _13515_ (.CLK(clknet_leaf_144_clk),
    .D(_00173_),
    .Q(\core_pipeline.pipeline_csr.instret[6] ));
 sky130_fd_sc_hd__dfxtp_1 _13516_ (.CLK(clknet_leaf_144_clk),
    .D(_00174_),
    .Q(\core_pipeline.pipeline_csr.instret[7] ));
 sky130_fd_sc_hd__dfxtp_1 _13517_ (.CLK(clknet_leaf_131_clk),
    .D(_00175_),
    .Q(\core_pipeline.pipeline_csr.instret[8] ));
 sky130_fd_sc_hd__dfxtp_2 _13518_ (.CLK(clknet_leaf_117_clk),
    .D(_00176_),
    .Q(\core_pipeline.pipeline_csr.instret[9] ));
 sky130_fd_sc_hd__dfxtp_1 _13519_ (.CLK(clknet_leaf_117_clk),
    .D(_00177_),
    .Q(\core_pipeline.pipeline_csr.instret[10] ));
 sky130_fd_sc_hd__dfxtp_1 _13520_ (.CLK(clknet_leaf_114_clk),
    .D(_00178_),
    .Q(\core_pipeline.pipeline_csr.instret[11] ));
 sky130_fd_sc_hd__dfxtp_1 _13521_ (.CLK(clknet_leaf_113_clk),
    .D(_00179_),
    .Q(\core_pipeline.pipeline_csr.instret[12] ));
 sky130_fd_sc_hd__dfxtp_1 _13522_ (.CLK(clknet_leaf_113_clk),
    .D(_00180_),
    .Q(\core_pipeline.pipeline_csr.instret[13] ));
 sky130_fd_sc_hd__dfxtp_1 _13523_ (.CLK(clknet_leaf_113_clk),
    .D(_00181_),
    .Q(\core_pipeline.pipeline_csr.instret[14] ));
 sky130_fd_sc_hd__dfxtp_1 _13524_ (.CLK(clknet_leaf_122_clk),
    .D(_00182_),
    .Q(\core_pipeline.pipeline_csr.instret[15] ));
 sky130_fd_sc_hd__dfxtp_1 _13525_ (.CLK(clknet_leaf_122_clk),
    .D(_00183_),
    .Q(\core_pipeline.pipeline_csr.instret[16] ));
 sky130_fd_sc_hd__dfxtp_1 _13526_ (.CLK(clknet_leaf_122_clk),
    .D(_00184_),
    .Q(\core_pipeline.pipeline_csr.instret[17] ));
 sky130_fd_sc_hd__dfxtp_1 _13527_ (.CLK(clknet_leaf_124_clk),
    .D(_00185_),
    .Q(\core_pipeline.pipeline_csr.instret[18] ));
 sky130_fd_sc_hd__dfxtp_2 _13528_ (.CLK(clknet_leaf_125_clk),
    .D(_00186_),
    .Q(\core_pipeline.pipeline_csr.instret[19] ));
 sky130_fd_sc_hd__dfxtp_1 _13529_ (.CLK(clknet_leaf_125_clk),
    .D(_00187_),
    .Q(\core_pipeline.pipeline_csr.instret[20] ));
 sky130_fd_sc_hd__dfxtp_1 _13530_ (.CLK(clknet_leaf_126_clk),
    .D(_00188_),
    .Q(\core_pipeline.pipeline_csr.instret[21] ));
 sky130_fd_sc_hd__dfxtp_1 _13531_ (.CLK(clknet_leaf_127_clk),
    .D(_00189_),
    .Q(\core_pipeline.pipeline_csr.instret[22] ));
 sky130_fd_sc_hd__dfxtp_1 _13532_ (.CLK(clknet_leaf_127_clk),
    .D(_00190_),
    .Q(\core_pipeline.pipeline_csr.instret[23] ));
 sky130_fd_sc_hd__dfxtp_1 _13533_ (.CLK(clknet_leaf_128_clk),
    .D(_00191_),
    .Q(\core_pipeline.pipeline_csr.instret[24] ));
 sky130_fd_sc_hd__dfxtp_1 _13534_ (.CLK(clknet_leaf_128_clk),
    .D(_00192_),
    .Q(\core_pipeline.pipeline_csr.instret[25] ));
 sky130_fd_sc_hd__dfxtp_1 _13535_ (.CLK(clknet_leaf_134_clk),
    .D(_00193_),
    .Q(\core_pipeline.pipeline_csr.instret[26] ));
 sky130_fd_sc_hd__dfxtp_1 _13536_ (.CLK(clknet_leaf_128_clk),
    .D(_00194_),
    .Q(\core_pipeline.pipeline_csr.instret[27] ));
 sky130_fd_sc_hd__dfxtp_1 _13537_ (.CLK(clknet_leaf_134_clk),
    .D(_00195_),
    .Q(\core_pipeline.pipeline_csr.instret[28] ));
 sky130_fd_sc_hd__dfxtp_1 _13538_ (.CLK(clknet_leaf_136_clk),
    .D(_00196_),
    .Q(\core_pipeline.pipeline_csr.instret[29] ));
 sky130_fd_sc_hd__dfxtp_2 _13539_ (.CLK(clknet_leaf_136_clk),
    .D(_00197_),
    .Q(\core_pipeline.pipeline_csr.instret[30] ));
 sky130_fd_sc_hd__dfxtp_1 _13540_ (.CLK(clknet_leaf_137_clk),
    .D(_00198_),
    .Q(\core_pipeline.pipeline_csr.instret[31] ));
 sky130_fd_sc_hd__dfxtp_2 _13541_ (.CLK(clknet_leaf_139_clk),
    .D(_00199_),
    .Q(\core_pipeline.pipeline_csr.instret[32] ));
 sky130_fd_sc_hd__dfxtp_2 _13542_ (.CLK(clknet_leaf_139_clk),
    .D(_00200_),
    .Q(\core_pipeline.pipeline_csr.instret[33] ));
 sky130_fd_sc_hd__dfxtp_1 _13543_ (.CLK(clknet_leaf_137_clk),
    .D(_00201_),
    .Q(\core_pipeline.pipeline_csr.instret[34] ));
 sky130_fd_sc_hd__dfxtp_2 _13544_ (.CLK(clknet_leaf_143_clk),
    .D(_00202_),
    .Q(\core_pipeline.pipeline_csr.instret[35] ));
 sky130_fd_sc_hd__dfxtp_1 _13545_ (.CLK(clknet_leaf_143_clk),
    .D(_00203_),
    .Q(\core_pipeline.pipeline_csr.instret[36] ));
 sky130_fd_sc_hd__dfxtp_1 _13546_ (.CLK(clknet_leaf_143_clk),
    .D(_00204_),
    .Q(\core_pipeline.pipeline_csr.instret[37] ));
 sky130_fd_sc_hd__dfxtp_1 _13547_ (.CLK(clknet_leaf_144_clk),
    .D(_00205_),
    .Q(\core_pipeline.pipeline_csr.instret[38] ));
 sky130_fd_sc_hd__dfxtp_1 _13548_ (.CLK(clknet_leaf_131_clk),
    .D(_00206_),
    .Q(\core_pipeline.pipeline_csr.instret[39] ));
 sky130_fd_sc_hd__dfxtp_1 _13549_ (.CLK(clknet_leaf_131_clk),
    .D(_00207_),
    .Q(\core_pipeline.pipeline_csr.instret[40] ));
 sky130_fd_sc_hd__dfxtp_1 _13550_ (.CLK(clknet_leaf_119_clk),
    .D(_00208_),
    .Q(\core_pipeline.pipeline_csr.instret[41] ));
 sky130_fd_sc_hd__dfxtp_1 _13551_ (.CLK(clknet_leaf_119_clk),
    .D(_00209_),
    .Q(\core_pipeline.pipeline_csr.instret[42] ));
 sky130_fd_sc_hd__dfxtp_1 _13552_ (.CLK(clknet_leaf_119_clk),
    .D(_00210_),
    .Q(\core_pipeline.pipeline_csr.instret[43] ));
 sky130_fd_sc_hd__dfxtp_1 _13553_ (.CLK(clknet_leaf_122_clk),
    .D(_00211_),
    .Q(\core_pipeline.pipeline_csr.instret[44] ));
 sky130_fd_sc_hd__dfxtp_1 _13554_ (.CLK(clknet_leaf_122_clk),
    .D(_00212_),
    .Q(\core_pipeline.pipeline_csr.instret[45] ));
 sky130_fd_sc_hd__dfxtp_2 _13555_ (.CLK(clknet_leaf_122_clk),
    .D(_00213_),
    .Q(\core_pipeline.pipeline_csr.instret[46] ));
 sky130_fd_sc_hd__dfxtp_1 _13556_ (.CLK(clknet_leaf_122_clk),
    .D(_00214_),
    .Q(\core_pipeline.pipeline_csr.instret[47] ));
 sky130_fd_sc_hd__dfxtp_1 _13557_ (.CLK(clknet_leaf_124_clk),
    .D(_00215_),
    .Q(\core_pipeline.pipeline_csr.instret[48] ));
 sky130_fd_sc_hd__dfxtp_2 _13558_ (.CLK(clknet_leaf_124_clk),
    .D(_00216_),
    .Q(\core_pipeline.pipeline_csr.instret[49] ));
 sky130_fd_sc_hd__dfxtp_1 _13559_ (.CLK(clknet_leaf_124_clk),
    .D(_00217_),
    .Q(\core_pipeline.pipeline_csr.instret[50] ));
 sky130_fd_sc_hd__dfxtp_1 _13560_ (.CLK(clknet_leaf_125_clk),
    .D(_00218_),
    .Q(\core_pipeline.pipeline_csr.instret[51] ));
 sky130_fd_sc_hd__dfxtp_2 _13561_ (.CLK(clknet_leaf_125_clk),
    .D(_00219_),
    .Q(\core_pipeline.pipeline_csr.instret[52] ));
 sky130_fd_sc_hd__dfxtp_1 _13562_ (.CLK(clknet_leaf_125_clk),
    .D(_00220_),
    .Q(\core_pipeline.pipeline_csr.instret[53] ));
 sky130_fd_sc_hd__dfxtp_2 _13563_ (.CLK(clknet_leaf_127_clk),
    .D(_00221_),
    .Q(\core_pipeline.pipeline_csr.instret[54] ));
 sky130_fd_sc_hd__dfxtp_1 _13564_ (.CLK(clknet_leaf_127_clk),
    .D(_00222_),
    .Q(\core_pipeline.pipeline_csr.instret[55] ));
 sky130_fd_sc_hd__dfxtp_1 _13565_ (.CLK(clknet_leaf_127_clk),
    .D(_00223_),
    .Q(\core_pipeline.pipeline_csr.instret[56] ));
 sky130_fd_sc_hd__dfxtp_2 _13566_ (.CLK(clknet_leaf_128_clk),
    .D(_00224_),
    .Q(\core_pipeline.pipeline_csr.instret[57] ));
 sky130_fd_sc_hd__dfxtp_2 _13567_ (.CLK(clknet_leaf_128_clk),
    .D(_00225_),
    .Q(\core_pipeline.pipeline_csr.instret[58] ));
 sky130_fd_sc_hd__dfxtp_1 _13568_ (.CLK(clknet_leaf_135_clk),
    .D(_00226_),
    .Q(\core_pipeline.pipeline_csr.instret[59] ));
 sky130_fd_sc_hd__dfxtp_2 _13569_ (.CLK(clknet_leaf_135_clk),
    .D(_00227_),
    .Q(\core_pipeline.pipeline_csr.instret[60] ));
 sky130_fd_sc_hd__dfxtp_1 _13570_ (.CLK(clknet_leaf_136_clk),
    .D(_00228_),
    .Q(\core_pipeline.pipeline_csr.instret[61] ));
 sky130_fd_sc_hd__dfxtp_1 _13571_ (.CLK(clknet_leaf_136_clk),
    .D(_00229_),
    .Q(\core_pipeline.pipeline_csr.instret[62] ));
 sky130_fd_sc_hd__dfxtp_1 _13572_ (.CLK(clknet_leaf_136_clk),
    .D(_00230_),
    .Q(\core_pipeline.pipeline_csr.instret[63] ));
 sky130_fd_sc_hd__dfxtp_1 _13573_ (.CLK(clknet_leaf_148_clk),
    .D(_00231_),
    .Q(\core_pipeline.pipeline_csr.pie ));
 sky130_fd_sc_hd__dfxtp_4 _13574_ (.CLK(clknet_leaf_148_clk),
    .D(_00232_),
    .Q(\core_pipeline.pipeline_csr.ie ));
 sky130_fd_sc_hd__dfxtp_2 _13575_ (.CLK(clknet_leaf_145_clk),
    .D(_00233_),
    .Q(\core_pipeline.pipeline_csr.meie ));
 sky130_fd_sc_hd__dfxtp_1 _13576_ (.CLK(clknet_leaf_148_clk),
    .D(_00234_),
    .Q(\core_pipeline.pipeline_csr.msie ));
 sky130_fd_sc_hd__dfxtp_1 _13577_ (.CLK(clknet_leaf_142_clk),
    .D(_00235_),
    .Q(\core_pipeline.pipeline_csr.msip ));
 sky130_fd_sc_hd__dfxtp_1 _13578_ (.CLK(clknet_leaf_145_clk),
    .D(_00003_),
    .Q(\core_pipeline.pipeline_csr.mtip ));
 sky130_fd_sc_hd__dfxtp_1 _13579_ (.CLK(clknet_leaf_145_clk),
    .D(_00236_),
    .Q(\core_pipeline.pipeline_csr.mtie ));
 sky130_fd_sc_hd__dfxtp_1 _13580_ (.CLK(clknet_leaf_93_clk),
    .D(_00005_),
    .Q(\core_pipeline.csr_to_fetch_mret_vector[0] ));
 sky130_fd_sc_hd__dfxtp_2 _13581_ (.CLK(clknet_leaf_153_clk),
    .D(_00016_),
    .Q(\core_pipeline.csr_to_fetch_mret_vector[1] ));
 sky130_fd_sc_hd__dfxtp_1 _13582_ (.CLK(clknet_leaf_150_clk),
    .D(_00027_),
    .Q(\core_pipeline.csr_to_fetch_mret_vector[2] ));
 sky130_fd_sc_hd__dfxtp_1 _13583_ (.CLK(clknet_leaf_151_clk),
    .D(_00030_),
    .Q(\core_pipeline.csr_to_fetch_mret_vector[3] ));
 sky130_fd_sc_hd__dfxtp_2 _13584_ (.CLK(clknet_leaf_93_clk),
    .D(_00031_),
    .Q(\core_pipeline.csr_to_fetch_mret_vector[4] ));
 sky130_fd_sc_hd__dfxtp_1 _13585_ (.CLK(clknet_leaf_147_clk),
    .D(_00032_),
    .Q(\core_pipeline.csr_to_fetch_mret_vector[5] ));
 sky130_fd_sc_hd__dfxtp_2 _13586_ (.CLK(clknet_leaf_95_clk),
    .D(_00033_),
    .Q(\core_pipeline.csr_to_fetch_mret_vector[6] ));
 sky130_fd_sc_hd__dfxtp_1 _13587_ (.CLK(clknet_leaf_98_clk),
    .D(_00034_),
    .Q(\core_pipeline.csr_to_fetch_mret_vector[7] ));
 sky130_fd_sc_hd__dfxtp_2 _13588_ (.CLK(clknet_leaf_103_clk),
    .D(_00035_),
    .Q(\core_pipeline.csr_to_fetch_mret_vector[8] ));
 sky130_fd_sc_hd__dfxtp_2 _13589_ (.CLK(clknet_leaf_107_clk),
    .D(_00036_),
    .Q(\core_pipeline.csr_to_fetch_mret_vector[9] ));
 sky130_fd_sc_hd__dfxtp_2 _13590_ (.CLK(clknet_leaf_107_clk),
    .D(_00006_),
    .Q(\core_pipeline.csr_to_fetch_mret_vector[10] ));
 sky130_fd_sc_hd__dfxtp_4 _13591_ (.CLK(clknet_leaf_107_clk),
    .D(_00007_),
    .Q(\core_pipeline.csr_to_fetch_mret_vector[11] ));
 sky130_fd_sc_hd__dfxtp_1 _13592_ (.CLK(clknet_leaf_107_clk),
    .D(_00008_),
    .Q(\core_pipeline.csr_to_fetch_mret_vector[12] ));
 sky130_fd_sc_hd__dfxtp_2 _13593_ (.CLK(clknet_leaf_108_clk),
    .D(_00009_),
    .Q(\core_pipeline.csr_to_fetch_mret_vector[13] ));
 sky130_fd_sc_hd__dfxtp_2 _13594_ (.CLK(clknet_leaf_108_clk),
    .D(_00010_),
    .Q(\core_pipeline.csr_to_fetch_mret_vector[14] ));
 sky130_fd_sc_hd__dfxtp_2 _13595_ (.CLK(clknet_leaf_108_clk),
    .D(_00011_),
    .Q(\core_pipeline.csr_to_fetch_mret_vector[15] ));
 sky130_fd_sc_hd__dfxtp_2 _13596_ (.CLK(clknet_leaf_108_clk),
    .D(_00012_),
    .Q(\core_pipeline.csr_to_fetch_mret_vector[16] ));
 sky130_fd_sc_hd__dfxtp_2 _13597_ (.CLK(clknet_leaf_111_clk),
    .D(_00013_),
    .Q(\core_pipeline.csr_to_fetch_mret_vector[17] ));
 sky130_fd_sc_hd__dfxtp_2 _13598_ (.CLK(clknet_leaf_111_clk),
    .D(_00014_),
    .Q(\core_pipeline.csr_to_fetch_mret_vector[18] ));
 sky130_fd_sc_hd__dfxtp_2 _13599_ (.CLK(clknet_leaf_110_clk),
    .D(_00015_),
    .Q(\core_pipeline.csr_to_fetch_mret_vector[19] ));
 sky130_fd_sc_hd__dfxtp_2 _13600_ (.CLK(clknet_leaf_115_clk),
    .D(_00017_),
    .Q(\core_pipeline.csr_to_fetch_mret_vector[20] ));
 sky130_fd_sc_hd__dfxtp_2 _13601_ (.CLK(clknet_leaf_116_clk),
    .D(_00018_),
    .Q(\core_pipeline.csr_to_fetch_mret_vector[21] ));
 sky130_fd_sc_hd__dfxtp_2 _13602_ (.CLK(clknet_leaf_117_clk),
    .D(_00019_),
    .Q(\core_pipeline.csr_to_fetch_mret_vector[22] ));
 sky130_fd_sc_hd__dfxtp_2 _13603_ (.CLK(clknet_leaf_117_clk),
    .D(_00020_),
    .Q(\core_pipeline.csr_to_fetch_mret_vector[23] ));
 sky130_fd_sc_hd__dfxtp_2 _13604_ (.CLK(clknet_leaf_103_clk),
    .D(_00021_),
    .Q(\core_pipeline.csr_to_fetch_mret_vector[24] ));
 sky130_fd_sc_hd__dfxtp_2 _13605_ (.CLK(clknet_leaf_100_clk),
    .D(_00022_),
    .Q(\core_pipeline.csr_to_fetch_mret_vector[25] ));
 sky130_fd_sc_hd__dfxtp_1 _13606_ (.CLK(clknet_leaf_99_clk),
    .D(_00023_),
    .Q(\core_pipeline.csr_to_fetch_mret_vector[26] ));
 sky130_fd_sc_hd__dfxtp_1 _13607_ (.CLK(clknet_leaf_100_clk),
    .D(_00024_),
    .Q(\core_pipeline.csr_to_fetch_mret_vector[27] ));
 sky130_fd_sc_hd__dfxtp_2 _13608_ (.CLK(clknet_leaf_100_clk),
    .D(_00025_),
    .Q(\core_pipeline.csr_to_fetch_mret_vector[28] ));
 sky130_fd_sc_hd__dfxtp_2 _13609_ (.CLK(clknet_leaf_98_clk),
    .D(_00026_),
    .Q(\core_pipeline.csr_to_fetch_mret_vector[29] ));
 sky130_fd_sc_hd__dfxtp_2 _13610_ (.CLK(clknet_leaf_146_clk),
    .D(_00028_),
    .Q(\core_pipeline.csr_to_fetch_mret_vector[30] ));
 sky130_fd_sc_hd__dfxtp_1 _13611_ (.CLK(clknet_leaf_146_clk),
    .D(_00029_),
    .Q(\core_pipeline.csr_to_fetch_mret_vector[31] ));
 sky130_fd_sc_hd__dfxtp_1 _13612_ (.CLK(clknet_leaf_148_clk),
    .D(_00237_),
    .Q(\core_pipeline.pipeline_csr.mscratch[0] ));
 sky130_fd_sc_hd__dfxtp_1 _13613_ (.CLK(clknet_leaf_140_clk),
    .D(_00238_),
    .Q(\core_pipeline.pipeline_csr.mscratch[1] ));
 sky130_fd_sc_hd__dfxtp_1 _13614_ (.CLK(clknet_leaf_140_clk),
    .D(_00239_),
    .Q(\core_pipeline.pipeline_csr.mscratch[2] ));
 sky130_fd_sc_hd__dfxtp_1 _13615_ (.CLK(clknet_leaf_148_clk),
    .D(_00240_),
    .Q(\core_pipeline.pipeline_csr.mscratch[3] ));
 sky130_fd_sc_hd__dfxtp_1 _13616_ (.CLK(clknet_leaf_142_clk),
    .D(_00241_),
    .Q(\core_pipeline.pipeline_csr.mscratch[4] ));
 sky130_fd_sc_hd__dfxtp_1 _13617_ (.CLK(clknet_leaf_144_clk),
    .D(_00242_),
    .Q(\core_pipeline.pipeline_csr.mscratch[5] ));
 sky130_fd_sc_hd__dfxtp_1 _13618_ (.CLK(clknet_leaf_144_clk),
    .D(_00243_),
    .Q(\core_pipeline.pipeline_csr.mscratch[6] ));
 sky130_fd_sc_hd__dfxtp_1 _13619_ (.CLK(clknet_leaf_145_clk),
    .D(_00244_),
    .Q(\core_pipeline.pipeline_csr.mscratch[7] ));
 sky130_fd_sc_hd__dfxtp_1 _13620_ (.CLK(clknet_leaf_118_clk),
    .D(_00245_),
    .Q(\core_pipeline.pipeline_csr.mscratch[8] ));
 sky130_fd_sc_hd__dfxtp_1 _13621_ (.CLK(clknet_leaf_117_clk),
    .D(_00246_),
    .Q(\core_pipeline.pipeline_csr.mscratch[9] ));
 sky130_fd_sc_hd__dfxtp_1 _13622_ (.CLK(clknet_leaf_117_clk),
    .D(_00247_),
    .Q(\core_pipeline.pipeline_csr.mscratch[10] ));
 sky130_fd_sc_hd__dfxtp_1 _13623_ (.CLK(clknet_leaf_100_clk),
    .D(_00248_),
    .Q(\core_pipeline.pipeline_csr.mscratch[11] ));
 sky130_fd_sc_hd__dfxtp_1 _13624_ (.CLK(clknet_leaf_113_clk),
    .D(_00249_),
    .Q(\core_pipeline.pipeline_csr.mscratch[12] ));
 sky130_fd_sc_hd__dfxtp_1 _13625_ (.CLK(clknet_leaf_114_clk),
    .D(_00250_),
    .Q(\core_pipeline.pipeline_csr.mscratch[13] ));
 sky130_fd_sc_hd__dfxtp_1 _13626_ (.CLK(clknet_leaf_121_clk),
    .D(_00251_),
    .Q(\core_pipeline.pipeline_csr.mscratch[14] ));
 sky130_fd_sc_hd__dfxtp_1 _13627_ (.CLK(clknet_leaf_122_clk),
    .D(_00252_),
    .Q(\core_pipeline.pipeline_csr.mscratch[15] ));
 sky130_fd_sc_hd__dfxtp_1 _13628_ (.CLK(clknet_leaf_113_clk),
    .D(_00253_),
    .Q(\core_pipeline.pipeline_csr.mscratch[16] ));
 sky130_fd_sc_hd__dfxtp_1 _13629_ (.CLK(clknet_leaf_124_clk),
    .D(_00254_),
    .Q(\core_pipeline.pipeline_csr.mscratch[17] ));
 sky130_fd_sc_hd__dfxtp_1 _13630_ (.CLK(clknet_leaf_124_clk),
    .D(_00255_),
    .Q(\core_pipeline.pipeline_csr.mscratch[18] ));
 sky130_fd_sc_hd__dfxtp_1 _13631_ (.CLK(clknet_leaf_120_clk),
    .D(_00256_),
    .Q(\core_pipeline.pipeline_csr.mscratch[19] ));
 sky130_fd_sc_hd__dfxtp_1 _13632_ (.CLK(clknet_leaf_125_clk),
    .D(_00257_),
    .Q(\core_pipeline.pipeline_csr.mscratch[20] ));
 sky130_fd_sc_hd__dfxtp_1 _13633_ (.CLK(clknet_leaf_126_clk),
    .D(_00258_),
    .Q(\core_pipeline.pipeline_csr.mscratch[21] ));
 sky130_fd_sc_hd__dfxtp_1 _13634_ (.CLK(clknet_leaf_129_clk),
    .D(_00259_),
    .Q(\core_pipeline.pipeline_csr.mscratch[22] ));
 sky130_fd_sc_hd__dfxtp_1 _13635_ (.CLK(clknet_leaf_129_clk),
    .D(_00260_),
    .Q(\core_pipeline.pipeline_csr.mscratch[23] ));
 sky130_fd_sc_hd__dfxtp_1 _13636_ (.CLK(clknet_leaf_129_clk),
    .D(_00261_),
    .Q(\core_pipeline.pipeline_csr.mscratch[24] ));
 sky130_fd_sc_hd__dfxtp_1 _13637_ (.CLK(clknet_leaf_128_clk),
    .D(_00262_),
    .Q(\core_pipeline.pipeline_csr.mscratch[25] ));
 sky130_fd_sc_hd__dfxtp_1 _13638_ (.CLK(clknet_leaf_131_clk),
    .D(_00263_),
    .Q(\core_pipeline.pipeline_csr.mscratch[26] ));
 sky130_fd_sc_hd__dfxtp_1 _13639_ (.CLK(clknet_leaf_100_clk),
    .D(_00264_),
    .Q(\core_pipeline.pipeline_csr.mscratch[27] ));
 sky130_fd_sc_hd__dfxtp_1 _13640_ (.CLK(clknet_leaf_133_clk),
    .D(_00265_),
    .Q(\core_pipeline.pipeline_csr.mscratch[28] ));
 sky130_fd_sc_hd__dfxtp_1 _13641_ (.CLK(clknet_leaf_132_clk),
    .D(_00266_),
    .Q(\core_pipeline.pipeline_csr.mscratch[29] ));
 sky130_fd_sc_hd__dfxtp_1 _13642_ (.CLK(clknet_leaf_136_clk),
    .D(_00267_),
    .Q(\core_pipeline.pipeline_csr.mscratch[30] ));
 sky130_fd_sc_hd__dfxtp_1 _13643_ (.CLK(clknet_leaf_137_clk),
    .D(_00268_),
    .Q(\core_pipeline.pipeline_csr.mscratch[31] ));
 sky130_fd_sc_hd__dfxtp_1 _13644_ (.CLK(clknet_leaf_142_clk),
    .D(_00269_),
    .Q(\core_pipeline.pipeline_csr.mcause[0] ));
 sky130_fd_sc_hd__dfxtp_1 _13645_ (.CLK(clknet_leaf_142_clk),
    .D(_00270_),
    .Q(\core_pipeline.pipeline_csr.mcause[1] ));
 sky130_fd_sc_hd__dfxtp_1 _13646_ (.CLK(clknet_leaf_142_clk),
    .D(_00271_),
    .Q(\core_pipeline.pipeline_csr.mcause[2] ));
 sky130_fd_sc_hd__dfxtp_1 _13647_ (.CLK(clknet_leaf_148_clk),
    .D(_00272_),
    .Q(\core_pipeline.pipeline_csr.mcause[3] ));
 sky130_fd_sc_hd__dfxtp_1 _13648_ (.CLK(clknet_leaf_142_clk),
    .D(_00273_),
    .Q(\core_pipeline.pipeline_csr.minterupt ));
 sky130_fd_sc_hd__dfxtp_1 _13649_ (.CLK(clknet_leaf_91_clk),
    .D(_00274_),
    .Q(\core_pipeline.memory_to_writeback_load_data[0] ));
 sky130_fd_sc_hd__dfxtp_1 _13650_ (.CLK(clknet_leaf_93_clk),
    .D(_00275_),
    .Q(\core_pipeline.memory_to_writeback_load_data[1] ));
 sky130_fd_sc_hd__dfxtp_1 _13651_ (.CLK(clknet_leaf_92_clk),
    .D(_00276_),
    .Q(\core_pipeline.memory_to_writeback_load_data[2] ));
 sky130_fd_sc_hd__dfxtp_1 _13652_ (.CLK(clknet_leaf_93_clk),
    .D(_00277_),
    .Q(\core_pipeline.memory_to_writeback_load_data[3] ));
 sky130_fd_sc_hd__dfxtp_1 _13653_ (.CLK(clknet_leaf_88_clk),
    .D(_00278_),
    .Q(\core_pipeline.memory_to_writeback_load_data[4] ));
 sky130_fd_sc_hd__dfxtp_1 _13654_ (.CLK(clknet_leaf_93_clk),
    .D(_00279_),
    .Q(\core_pipeline.memory_to_writeback_load_data[5] ));
 sky130_fd_sc_hd__dfxtp_1 _13655_ (.CLK(clknet_leaf_88_clk),
    .D(_00280_),
    .Q(\core_pipeline.memory_to_writeback_load_data[6] ));
 sky130_fd_sc_hd__dfxtp_1 _13656_ (.CLK(clknet_leaf_90_clk),
    .D(_00281_),
    .Q(\core_pipeline.memory_to_writeback_load_data[7] ));
 sky130_fd_sc_hd__dfxtp_1 _13657_ (.CLK(clknet_leaf_80_clk),
    .D(_00282_),
    .Q(\core_pipeline.memory_to_writeback_load_data[8] ));
 sky130_fd_sc_hd__dfxtp_1 _13658_ (.CLK(clknet_leaf_80_clk),
    .D(_00283_),
    .Q(\core_pipeline.memory_to_writeback_load_data[9] ));
 sky130_fd_sc_hd__dfxtp_1 _13659_ (.CLK(clknet_leaf_80_clk),
    .D(_00284_),
    .Q(\core_pipeline.memory_to_writeback_load_data[10] ));
 sky130_fd_sc_hd__dfxtp_1 _13660_ (.CLK(clknet_leaf_86_clk),
    .D(_00285_),
    .Q(\core_pipeline.memory_to_writeback_load_data[11] ));
 sky130_fd_sc_hd__dfxtp_1 _13661_ (.CLK(clknet_leaf_80_clk),
    .D(_00286_),
    .Q(\core_pipeline.memory_to_writeback_load_data[12] ));
 sky130_fd_sc_hd__dfxtp_1 _13662_ (.CLK(clknet_leaf_86_clk),
    .D(_00287_),
    .Q(\core_pipeline.memory_to_writeback_load_data[13] ));
 sky130_fd_sc_hd__dfxtp_1 _13663_ (.CLK(clknet_leaf_80_clk),
    .D(_00288_),
    .Q(\core_pipeline.memory_to_writeback_load_data[14] ));
 sky130_fd_sc_hd__dfxtp_1 _13664_ (.CLK(clknet_leaf_79_clk),
    .D(_00289_),
    .Q(\core_pipeline.memory_to_writeback_load_data[15] ));
 sky130_fd_sc_hd__dfxtp_1 _13665_ (.CLK(clknet_leaf_79_clk),
    .D(_00290_),
    .Q(\core_pipeline.memory_to_writeback_load_data[16] ));
 sky130_fd_sc_hd__dfxtp_1 _13666_ (.CLK(clknet_leaf_105_clk),
    .D(_00291_),
    .Q(\core_pipeline.memory_to_writeback_load_data[17] ));
 sky130_fd_sc_hd__dfxtp_1 _13667_ (.CLK(clknet_leaf_80_clk),
    .D(_00292_),
    .Q(\core_pipeline.memory_to_writeback_load_data[18] ));
 sky130_fd_sc_hd__dfxtp_1 _13668_ (.CLK(clknet_leaf_79_clk),
    .D(_00293_),
    .Q(\core_pipeline.memory_to_writeback_load_data[19] ));
 sky130_fd_sc_hd__dfxtp_1 _13669_ (.CLK(clknet_leaf_96_clk),
    .D(_00294_),
    .Q(\core_pipeline.memory_to_writeback_load_data[20] ));
 sky130_fd_sc_hd__dfxtp_1 _13670_ (.CLK(clknet_leaf_96_clk),
    .D(_00295_),
    .Q(\core_pipeline.memory_to_writeback_load_data[21] ));
 sky130_fd_sc_hd__dfxtp_1 _13671_ (.CLK(clknet_leaf_104_clk),
    .D(_00296_),
    .Q(\core_pipeline.memory_to_writeback_load_data[22] ));
 sky130_fd_sc_hd__dfxtp_1 _13672_ (.CLK(clknet_leaf_87_clk),
    .D(_00297_),
    .Q(\core_pipeline.memory_to_writeback_load_data[23] ));
 sky130_fd_sc_hd__dfxtp_1 _13673_ (.CLK(clknet_leaf_79_clk),
    .D(_00298_),
    .Q(\core_pipeline.memory_to_writeback_load_data[24] ));
 sky130_fd_sc_hd__dfxtp_1 _13674_ (.CLK(clknet_leaf_79_clk),
    .D(_00299_),
    .Q(\core_pipeline.memory_to_writeback_load_data[25] ));
 sky130_fd_sc_hd__dfxtp_1 _13675_ (.CLK(clknet_leaf_87_clk),
    .D(_00300_),
    .Q(\core_pipeline.memory_to_writeback_load_data[26] ));
 sky130_fd_sc_hd__dfxtp_1 _13676_ (.CLK(clknet_leaf_96_clk),
    .D(_00301_),
    .Q(\core_pipeline.memory_to_writeback_load_data[27] ));
 sky130_fd_sc_hd__dfxtp_1 _13677_ (.CLK(clknet_leaf_95_clk),
    .D(_00302_),
    .Q(\core_pipeline.memory_to_writeback_load_data[28] ));
 sky130_fd_sc_hd__dfxtp_1 _13678_ (.CLK(clknet_leaf_88_clk),
    .D(_00303_),
    .Q(\core_pipeline.memory_to_writeback_load_data[29] ));
 sky130_fd_sc_hd__dfxtp_1 _13679_ (.CLK(clknet_leaf_95_clk),
    .D(_00304_),
    .Q(\core_pipeline.memory_to_writeback_load_data[30] ));
 sky130_fd_sc_hd__dfxtp_1 _13680_ (.CLK(clknet_leaf_88_clk),
    .D(_00305_),
    .Q(\core_pipeline.memory_to_writeback_load_data[31] ));
 sky130_fd_sc_hd__dfxtp_1 _13681_ (.CLK(clknet_leaf_245_clk),
    .D(_00306_),
    .Q(\core_pipeline.pipeline_registers.registers[31][0] ));
 sky130_fd_sc_hd__dfxtp_1 _13682_ (.CLK(clknet_leaf_165_clk),
    .D(_00307_),
    .Q(\core_pipeline.pipeline_registers.registers[31][1] ));
 sky130_fd_sc_hd__dfxtp_1 _13683_ (.CLK(clknet_leaf_192_clk),
    .D(_00308_),
    .Q(\core_pipeline.pipeline_registers.registers[31][2] ));
 sky130_fd_sc_hd__dfxtp_1 _13684_ (.CLK(clknet_leaf_237_clk),
    .D(_00309_),
    .Q(\core_pipeline.pipeline_registers.registers[31][3] ));
 sky130_fd_sc_hd__dfxtp_1 _13685_ (.CLK(clknet_leaf_245_clk),
    .D(_00310_),
    .Q(\core_pipeline.pipeline_registers.registers[31][4] ));
 sky130_fd_sc_hd__dfxtp_1 _13686_ (.CLK(clknet_leaf_201_clk),
    .D(_00311_),
    .Q(\core_pipeline.pipeline_registers.registers[31][5] ));
 sky130_fd_sc_hd__dfxtp_1 _13687_ (.CLK(clknet_leaf_205_clk),
    .D(_00312_),
    .Q(\core_pipeline.pipeline_registers.registers[31][6] ));
 sky130_fd_sc_hd__dfxtp_1 _13688_ (.CLK(clknet_leaf_234_clk),
    .D(_00313_),
    .Q(\core_pipeline.pipeline_registers.registers[31][7] ));
 sky130_fd_sc_hd__dfxtp_1 _13689_ (.CLK(clknet_leaf_241_clk),
    .D(_00314_),
    .Q(\core_pipeline.pipeline_registers.registers[31][8] ));
 sky130_fd_sc_hd__dfxtp_1 _13690_ (.CLK(clknet_leaf_248_clk),
    .D(_00315_),
    .Q(\core_pipeline.pipeline_registers.registers[31][9] ));
 sky130_fd_sc_hd__dfxtp_1 _13691_ (.CLK(clknet_leaf_23_clk),
    .D(_00316_),
    .Q(\core_pipeline.pipeline_registers.registers[31][10] ));
 sky130_fd_sc_hd__dfxtp_1 _13692_ (.CLK(clknet_leaf_247_clk),
    .D(_00317_),
    .Q(\core_pipeline.pipeline_registers.registers[31][11] ));
 sky130_fd_sc_hd__dfxtp_1 _13693_ (.CLK(clknet_leaf_229_clk),
    .D(_00318_),
    .Q(\core_pipeline.pipeline_registers.registers[31][12] ));
 sky130_fd_sc_hd__dfxtp_1 _13694_ (.CLK(clknet_leaf_21_clk),
    .D(_00319_),
    .Q(\core_pipeline.pipeline_registers.registers[31][13] ));
 sky130_fd_sc_hd__dfxtp_1 _13695_ (.CLK(clknet_leaf_6_clk),
    .D(_00320_),
    .Q(\core_pipeline.pipeline_registers.registers[31][14] ));
 sky130_fd_sc_hd__dfxtp_1 _13696_ (.CLK(clknet_leaf_26_clk),
    .D(_00321_),
    .Q(\core_pipeline.pipeline_registers.registers[31][15] ));
 sky130_fd_sc_hd__dfxtp_1 _13697_ (.CLK(clknet_leaf_242_clk),
    .D(_00322_),
    .Q(\core_pipeline.pipeline_registers.registers[31][16] ));
 sky130_fd_sc_hd__dfxtp_1 _13698_ (.CLK(clknet_leaf_196_clk),
    .D(_00323_),
    .Q(\core_pipeline.pipeline_registers.registers[31][17] ));
 sky130_fd_sc_hd__dfxtp_1 _13699_ (.CLK(clknet_leaf_181_clk),
    .D(_00324_),
    .Q(\core_pipeline.pipeline_registers.registers[31][18] ));
 sky130_fd_sc_hd__dfxtp_1 _13700_ (.CLK(clknet_leaf_194_clk),
    .D(_00325_),
    .Q(\core_pipeline.pipeline_registers.registers[31][19] ));
 sky130_fd_sc_hd__dfxtp_1 _13701_ (.CLK(clknet_leaf_189_clk),
    .D(_00326_),
    .Q(\core_pipeline.pipeline_registers.registers[31][20] ));
 sky130_fd_sc_hd__dfxtp_1 _13702_ (.CLK(clknet_leaf_173_clk),
    .D(_00327_),
    .Q(\core_pipeline.pipeline_registers.registers[31][21] ));
 sky130_fd_sc_hd__dfxtp_1 _13703_ (.CLK(clknet_leaf_197_clk),
    .D(_00328_),
    .Q(\core_pipeline.pipeline_registers.registers[31][22] ));
 sky130_fd_sc_hd__dfxtp_1 _13704_ (.CLK(clknet_leaf_217_clk),
    .D(_00329_),
    .Q(\core_pipeline.pipeline_registers.registers[31][23] ));
 sky130_fd_sc_hd__dfxtp_1 _13705_ (.CLK(clknet_leaf_226_clk),
    .D(_00330_),
    .Q(\core_pipeline.pipeline_registers.registers[31][24] ));
 sky130_fd_sc_hd__dfxtp_1 _13706_ (.CLK(clknet_leaf_24_clk),
    .D(_00331_),
    .Q(\core_pipeline.pipeline_registers.registers[31][25] ));
 sky130_fd_sc_hd__dfxtp_1 _13707_ (.CLK(clknet_leaf_28_clk),
    .D(_00332_),
    .Q(\core_pipeline.pipeline_registers.registers[31][26] ));
 sky130_fd_sc_hd__dfxtp_1 _13708_ (.CLK(clknet_leaf_165_clk),
    .D(_00333_),
    .Q(\core_pipeline.pipeline_registers.registers[31][27] ));
 sky130_fd_sc_hd__dfxtp_1 _13709_ (.CLK(clknet_leaf_183_clk),
    .D(_00334_),
    .Q(\core_pipeline.pipeline_registers.registers[31][28] ));
 sky130_fd_sc_hd__dfxtp_1 _13710_ (.CLK(clknet_leaf_197_clk),
    .D(_00335_),
    .Q(\core_pipeline.pipeline_registers.registers[31][29] ));
 sky130_fd_sc_hd__dfxtp_1 _13711_ (.CLK(clknet_leaf_207_clk),
    .D(_00336_),
    .Q(\core_pipeline.pipeline_registers.registers[31][30] ));
 sky130_fd_sc_hd__dfxtp_1 _13712_ (.CLK(clknet_leaf_175_clk),
    .D(_00337_),
    .Q(\core_pipeline.pipeline_registers.registers[31][31] ));
 sky130_fd_sc_hd__dfxtp_1 _13713_ (.CLK(clknet_leaf_43_clk),
    .D(_00338_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_sll[0] ));
 sky130_fd_sc_hd__dfxtp_1 _13714_ (.CLK(clknet_leaf_49_clk),
    .D(_00339_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_sll[1] ));
 sky130_fd_sc_hd__dfxtp_1 _13715_ (.CLK(clknet_leaf_49_clk),
    .D(_00340_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_sll[2] ));
 sky130_fd_sc_hd__dfxtp_1 _13716_ (.CLK(clknet_leaf_50_clk),
    .D(_00341_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_sll[3] ));
 sky130_fd_sc_hd__dfxtp_1 _13717_ (.CLK(clknet_leaf_50_clk),
    .D(_00342_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_sll[4] ));
 sky130_fd_sc_hd__dfxtp_1 _13718_ (.CLK(clknet_leaf_50_clk),
    .D(_00343_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_sll[5] ));
 sky130_fd_sc_hd__dfxtp_1 _13719_ (.CLK(clknet_leaf_52_clk),
    .D(_00344_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_sll[6] ));
 sky130_fd_sc_hd__dfxtp_2 _13720_ (.CLK(clknet_leaf_51_clk),
    .D(_00345_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_sll[7] ));
 sky130_fd_sc_hd__dfxtp_1 _13721_ (.CLK(clknet_leaf_60_clk),
    .D(_00346_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_sll[8] ));
 sky130_fd_sc_hd__dfxtp_1 _13722_ (.CLK(clknet_leaf_61_clk),
    .D(_00347_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_sll[9] ));
 sky130_fd_sc_hd__dfxtp_1 _13723_ (.CLK(clknet_leaf_60_clk),
    .D(_00348_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_sll[10] ));
 sky130_fd_sc_hd__dfxtp_1 _13724_ (.CLK(clknet_leaf_61_clk),
    .D(_00349_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_sll[11] ));
 sky130_fd_sc_hd__dfxtp_1 _13725_ (.CLK(clknet_leaf_61_clk),
    .D(_00350_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_sll[12] ));
 sky130_fd_sc_hd__dfxtp_1 _13726_ (.CLK(clknet_leaf_60_clk),
    .D(_00351_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_sll[13] ));
 sky130_fd_sc_hd__dfxtp_1 _13727_ (.CLK(clknet_leaf_60_clk),
    .D(_00352_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_sll[14] ));
 sky130_fd_sc_hd__dfxtp_1 _13728_ (.CLK(clknet_leaf_59_clk),
    .D(_00353_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_sll[15] ));
 sky130_fd_sc_hd__dfxtp_2 _13729_ (.CLK(clknet_leaf_222_clk),
    .D(_00354_),
    .Q(\core_pipeline.decode_to_execute_rd_address[4] ));
 sky130_fd_sc_hd__dfxtp_2 _13730_ (.CLK(clknet_leaf_222_clk),
    .D(_00355_),
    .Q(\core_pipeline.decode_to_execute_rd_address[3] ));
 sky130_fd_sc_hd__dfxtp_2 _13731_ (.CLK(clknet_leaf_154_clk),
    .D(_00356_),
    .Q(\core_pipeline.decode_to_execute_rd_address[2] ));
 sky130_fd_sc_hd__dfxtp_2 _13732_ (.CLK(clknet_leaf_222_clk),
    .D(_00357_),
    .Q(\core_pipeline.decode_to_execute_rd_address[1] ));
 sky130_fd_sc_hd__dfxtp_2 _13733_ (.CLK(clknet_leaf_222_clk),
    .D(_00358_),
    .Q(\core_pipeline.decode_to_execute_rd_address[0] ));
 sky130_fd_sc_hd__dfxtp_1 _13734_ (.CLK(clknet_leaf_222_clk),
    .D(_00359_),
    .Q(\core_pipeline.decode_to_execute_write_select[1] ));
 sky130_fd_sc_hd__dfxtp_1 _13735_ (.CLK(clknet_leaf_34_clk),
    .D(_00360_),
    .Q(\core_pipeline.decode_to_execute_write_select[0] ));
 sky130_fd_sc_hd__dfxtp_1 _13736_ (.CLK(clknet_leaf_154_clk),
    .D(_00361_),
    .Q(\core_pipeline.decode_to_execute_bypass_memory ));
 sky130_fd_sc_hd__dfxtp_2 _13737_ (.CLK(clknet_leaf_154_clk),
    .D(_00362_),
    .Q(\core_pipeline.decode_to_execute_csr_write ));
 sky130_fd_sc_hd__dfxtp_1 _13738_ (.CLK(clknet_leaf_154_clk),
    .D(_00363_),
    .Q(\core_pipeline.decode_to_execute_csr_read ));
 sky130_fd_sc_hd__dfxtp_4 _13739_ (.CLK(clknet_leaf_37_clk),
    .D(_00364_),
    .Q(\core_pipeline.decode_to_execute_alu_function_modifier ));
 sky130_fd_sc_hd__dfxtp_4 _13740_ (.CLK(clknet_leaf_37_clk),
    .D(_00365_),
    .Q(\core_pipeline.decode_to_execute_alu_function[2] ));
 sky130_fd_sc_hd__dfxtp_4 _13741_ (.CLK(clknet_leaf_45_clk),
    .D(_00366_),
    .Q(\core_pipeline.decode_to_execute_alu_function[1] ));
 sky130_fd_sc_hd__dfxtp_4 _13742_ (.CLK(clknet_leaf_37_clk),
    .D(_00367_),
    .Q(\core_pipeline.decode_to_execute_alu_function[0] ));
 sky130_fd_sc_hd__dfxtp_1 _13743_ (.CLK(clknet_leaf_35_clk),
    .D(_00368_),
    .Q(\core_pipeline.decode_to_execute_imm_data[31] ));
 sky130_fd_sc_hd__dfxtp_1 _13744_ (.CLK(clknet_leaf_89_clk),
    .D(_00369_),
    .Q(\core_pipeline.decode_to_execute_imm_data[30] ));
 sky130_fd_sc_hd__dfxtp_1 _13745_ (.CLK(clknet_leaf_85_clk),
    .D(_00370_),
    .Q(\core_pipeline.decode_to_execute_imm_data[29] ));
 sky130_fd_sc_hd__dfxtp_1 _13746_ (.CLK(clknet_leaf_86_clk),
    .D(_00371_),
    .Q(\core_pipeline.decode_to_execute_imm_data[28] ));
 sky130_fd_sc_hd__dfxtp_1 _13747_ (.CLK(clknet_leaf_89_clk),
    .D(_00372_),
    .Q(\core_pipeline.decode_to_execute_imm_data[27] ));
 sky130_fd_sc_hd__dfxtp_1 _13748_ (.CLK(clknet_leaf_85_clk),
    .D(_00373_),
    .Q(\core_pipeline.decode_to_execute_imm_data[26] ));
 sky130_fd_sc_hd__dfxtp_1 _13749_ (.CLK(clknet_leaf_85_clk),
    .D(_00374_),
    .Q(\core_pipeline.decode_to_execute_imm_data[25] ));
 sky130_fd_sc_hd__dfxtp_1 _13750_ (.CLK(clknet_leaf_85_clk),
    .D(_00375_),
    .Q(\core_pipeline.decode_to_execute_imm_data[24] ));
 sky130_fd_sc_hd__dfxtp_1 _13751_ (.CLK(clknet_leaf_86_clk),
    .D(_00376_),
    .Q(\core_pipeline.decode_to_execute_imm_data[23] ));
 sky130_fd_sc_hd__dfxtp_1 _13752_ (.CLK(clknet_leaf_86_clk),
    .D(_00377_),
    .Q(\core_pipeline.decode_to_execute_imm_data[22] ));
 sky130_fd_sc_hd__dfxtp_1 _13753_ (.CLK(clknet_leaf_89_clk),
    .D(_00378_),
    .Q(\core_pipeline.decode_to_execute_imm_data[21] ));
 sky130_fd_sc_hd__dfxtp_1 _13754_ (.CLK(clknet_leaf_85_clk),
    .D(_00379_),
    .Q(\core_pipeline.decode_to_execute_imm_data[20] ));
 sky130_fd_sc_hd__dfxtp_1 _13755_ (.CLK(clknet_leaf_84_clk),
    .D(_00380_),
    .Q(\core_pipeline.decode_to_execute_imm_data[19] ));
 sky130_fd_sc_hd__dfxtp_1 _13756_ (.CLK(clknet_leaf_84_clk),
    .D(_00381_),
    .Q(\core_pipeline.decode_to_execute_imm_data[18] ));
 sky130_fd_sc_hd__dfxtp_1 _13757_ (.CLK(clknet_leaf_84_clk),
    .D(_00382_),
    .Q(\core_pipeline.decode_to_execute_imm_data[17] ));
 sky130_fd_sc_hd__dfxtp_1 _13758_ (.CLK(clknet_leaf_84_clk),
    .D(_00383_),
    .Q(\core_pipeline.decode_to_execute_imm_data[16] ));
 sky130_fd_sc_hd__dfxtp_2 _13759_ (.CLK(clknet_leaf_84_clk),
    .D(_00384_),
    .Q(\core_pipeline.decode_to_execute_imm_data[15] ));
 sky130_fd_sc_hd__dfxtp_1 _13760_ (.CLK(clknet_leaf_84_clk),
    .D(_00385_),
    .Q(\core_pipeline.decode_to_execute_imm_data[14] ));
 sky130_fd_sc_hd__dfxtp_1 _13761_ (.CLK(clknet_leaf_84_clk),
    .D(_00386_),
    .Q(\core_pipeline.decode_to_execute_imm_data[13] ));
 sky130_fd_sc_hd__dfxtp_1 _13762_ (.CLK(clknet_leaf_84_clk),
    .D(_00387_),
    .Q(\core_pipeline.decode_to_execute_imm_data[12] ));
 sky130_fd_sc_hd__dfxtp_1 _13763_ (.CLK(clknet_leaf_41_clk),
    .D(_00388_),
    .Q(\core_pipeline.decode_to_execute_imm_data[11] ));
 sky130_fd_sc_hd__dfxtp_1 _13764_ (.CLK(clknet_leaf_84_clk),
    .D(_00389_),
    .Q(\core_pipeline.decode_to_execute_imm_data[10] ));
 sky130_fd_sc_hd__dfxtp_1 _13765_ (.CLK(clknet_leaf_89_clk),
    .D(_00390_),
    .Q(\core_pipeline.decode_to_execute_imm_data[9] ));
 sky130_fd_sc_hd__dfxtp_1 _13766_ (.CLK(clknet_leaf_84_clk),
    .D(_00391_),
    .Q(\core_pipeline.decode_to_execute_imm_data[8] ));
 sky130_fd_sc_hd__dfxtp_1 _13767_ (.CLK(clknet_leaf_36_clk),
    .D(_00392_),
    .Q(\core_pipeline.decode_to_execute_imm_data[7] ));
 sky130_fd_sc_hd__dfxtp_1 _13768_ (.CLK(clknet_leaf_40_clk),
    .D(_00393_),
    .Q(\core_pipeline.decode_to_execute_imm_data[6] ));
 sky130_fd_sc_hd__dfxtp_1 _13769_ (.CLK(clknet_leaf_37_clk),
    .D(_00394_),
    .Q(\core_pipeline.decode_to_execute_imm_data[5] ));
 sky130_fd_sc_hd__dfxtp_1 _13770_ (.CLK(clknet_leaf_39_clk),
    .D(_00395_),
    .Q(\core_pipeline.decode_to_execute_imm_data[4] ));
 sky130_fd_sc_hd__dfxtp_1 _13771_ (.CLK(clknet_leaf_36_clk),
    .D(_00396_),
    .Q(\core_pipeline.decode_to_execute_imm_data[3] ));
 sky130_fd_sc_hd__dfxtp_1 _13772_ (.CLK(clknet_leaf_35_clk),
    .D(_00397_),
    .Q(\core_pipeline.decode_to_execute_imm_data[2] ));
 sky130_fd_sc_hd__dfxtp_1 _13773_ (.CLK(clknet_leaf_37_clk),
    .D(_00398_),
    .Q(\core_pipeline.decode_to_execute_imm_data[1] ));
 sky130_fd_sc_hd__dfxtp_2 _13774_ (.CLK(clknet_leaf_38_clk),
    .D(_00399_),
    .Q(\core_pipeline.decode_to_execute_imm_data[0] ));
 sky130_fd_sc_hd__dfxtp_4 _13775_ (.CLK(clknet_leaf_137_clk),
    .D(_00400_),
    .Q(\core_pipeline.decode_to_execute_csr_data[31] ));
 sky130_fd_sc_hd__dfxtp_4 _13776_ (.CLK(clknet_leaf_133_clk),
    .D(_00401_),
    .Q(\core_pipeline.decode_to_execute_csr_data[30] ));
 sky130_fd_sc_hd__dfxtp_4 _13777_ (.CLK(clknet_leaf_132_clk),
    .D(_00402_),
    .Q(\core_pipeline.decode_to_execute_csr_data[29] ));
 sky130_fd_sc_hd__dfxtp_4 _13778_ (.CLK(clknet_leaf_133_clk),
    .D(_00403_),
    .Q(\core_pipeline.decode_to_execute_csr_data[28] ));
 sky130_fd_sc_hd__dfxtp_4 _13779_ (.CLK(clknet_leaf_132_clk),
    .D(_00404_),
    .Q(\core_pipeline.decode_to_execute_csr_data[27] ));
 sky130_fd_sc_hd__dfxtp_4 _13780_ (.CLK(clknet_leaf_132_clk),
    .D(_00405_),
    .Q(\core_pipeline.decode_to_execute_csr_data[26] ));
 sky130_fd_sc_hd__dfxtp_4 _13781_ (.CLK(clknet_leaf_130_clk),
    .D(_00406_),
    .Q(\core_pipeline.decode_to_execute_csr_data[25] ));
 sky130_fd_sc_hd__dfxtp_4 _13782_ (.CLK(clknet_leaf_130_clk),
    .D(_00407_),
    .Q(\core_pipeline.decode_to_execute_csr_data[24] ));
 sky130_fd_sc_hd__dfxtp_4 _13783_ (.CLK(clknet_leaf_129_clk),
    .D(_00408_),
    .Q(\core_pipeline.decode_to_execute_csr_data[23] ));
 sky130_fd_sc_hd__dfxtp_4 _13784_ (.CLK(clknet_leaf_129_clk),
    .D(_00409_),
    .Q(\core_pipeline.decode_to_execute_csr_data[22] ));
 sky130_fd_sc_hd__dfxtp_4 _13785_ (.CLK(clknet_leaf_119_clk),
    .D(_00410_),
    .Q(\core_pipeline.decode_to_execute_csr_data[21] ));
 sky130_fd_sc_hd__dfxtp_4 _13786_ (.CLK(clknet_leaf_130_clk),
    .D(_00411_),
    .Q(\core_pipeline.decode_to_execute_csr_data[20] ));
 sky130_fd_sc_hd__dfxtp_4 _13787_ (.CLK(clknet_leaf_120_clk),
    .D(_00412_),
    .Q(\core_pipeline.decode_to_execute_csr_data[19] ));
 sky130_fd_sc_hd__dfxtp_4 _13788_ (.CLK(clknet_leaf_119_clk),
    .D(_00413_),
    .Q(\core_pipeline.decode_to_execute_csr_data[18] ));
 sky130_fd_sc_hd__dfxtp_4 _13789_ (.CLK(clknet_leaf_123_clk),
    .D(_00414_),
    .Q(\core_pipeline.decode_to_execute_csr_data[17] ));
 sky130_fd_sc_hd__dfxtp_2 _13790_ (.CLK(clknet_leaf_72_clk),
    .D(_00415_),
    .Q(\core_pipeline.decode_to_execute_csr_data[16] ));
 sky130_fd_sc_hd__dfxtp_4 _13791_ (.CLK(clknet_leaf_74_clk),
    .D(_00416_),
    .Q(\core_pipeline.decode_to_execute_csr_data[15] ));
 sky130_fd_sc_hd__dfxtp_2 _13792_ (.CLK(clknet_leaf_78_clk),
    .D(_00417_),
    .Q(\core_pipeline.decode_to_execute_csr_data[14] ));
 sky130_fd_sc_hd__dfxtp_2 _13793_ (.CLK(clknet_leaf_72_clk),
    .D(_00418_),
    .Q(\core_pipeline.decode_to_execute_csr_data[13] ));
 sky130_fd_sc_hd__dfxtp_2 _13794_ (.CLK(clknet_leaf_73_clk),
    .D(_00419_),
    .Q(\core_pipeline.decode_to_execute_csr_data[12] ));
 sky130_fd_sc_hd__dfxtp_4 _13795_ (.CLK(clknet_leaf_145_clk),
    .D(_00420_),
    .Q(\core_pipeline.decode_to_execute_csr_data[11] ));
 sky130_fd_sc_hd__dfxtp_1 _13796_ (.CLK(clknet_leaf_82_clk),
    .D(_00421_),
    .Q(\core_pipeline.decode_to_execute_csr_data[10] ));
 sky130_fd_sc_hd__dfxtp_1 _13797_ (.CLK(clknet_leaf_82_clk),
    .D(_00422_),
    .Q(\core_pipeline.decode_to_execute_csr_data[9] ));
 sky130_fd_sc_hd__dfxtp_4 _13798_ (.CLK(clknet_leaf_131_clk),
    .D(_00423_),
    .Q(\core_pipeline.decode_to_execute_csr_data[8] ));
 sky130_fd_sc_hd__dfxtp_4 _13799_ (.CLK(clknet_leaf_146_clk),
    .D(_00424_),
    .Q(\core_pipeline.decode_to_execute_csr_data[7] ));
 sky130_fd_sc_hd__dfxtp_1 _13800_ (.CLK(clknet_leaf_85_clk),
    .D(_00425_),
    .Q(\core_pipeline.decode_to_execute_csr_data[6] ));
 sky130_fd_sc_hd__dfxtp_2 _13801_ (.CLK(clknet_leaf_94_clk),
    .D(_00426_),
    .Q(\core_pipeline.decode_to_execute_csr_data[5] ));
 sky130_fd_sc_hd__dfxtp_1 _13802_ (.CLK(clknet_leaf_39_clk),
    .D(_00427_),
    .Q(\core_pipeline.decode_to_execute_csr_data[4] ));
 sky130_fd_sc_hd__dfxtp_2 _13803_ (.CLK(clknet_leaf_148_clk),
    .D(_00428_),
    .Q(\core_pipeline.decode_to_execute_csr_data[3] ));
 sky130_fd_sc_hd__dfxtp_4 _13804_ (.CLK(clknet_leaf_142_clk),
    .D(_00429_),
    .Q(\core_pipeline.decode_to_execute_csr_data[2] ));
 sky130_fd_sc_hd__dfxtp_2 _13805_ (.CLK(clknet_leaf_37_clk),
    .D(_00430_),
    .Q(\core_pipeline.decode_to_execute_csr_data[1] ));
 sky130_fd_sc_hd__dfxtp_1 _13806_ (.CLK(clknet_leaf_38_clk),
    .D(_00431_),
    .Q(\core_pipeline.decode_to_execute_csr_data[0] ));
 sky130_fd_sc_hd__dfxtp_1 _13807_ (.CLK(clknet_leaf_156_clk),
    .D(_00432_),
    .Q(\core_pipeline.decode_to_execute_exception ));
 sky130_fd_sc_hd__dfxtp_1 _13808_ (.CLK(clknet_leaf_157_clk),
    .D(_00433_),
    .Q(\core_pipeline.decode_to_execute_ecause[3] ));
 sky130_fd_sc_hd__dfxtp_1 _13809_ (.CLK(clknet_leaf_157_clk),
    .D(_00434_),
    .Q(\core_pipeline.decode_to_execute_ecause[1] ));
 sky130_fd_sc_hd__dfxtp_1 _13810_ (.CLK(clknet_leaf_157_clk),
    .D(_00435_),
    .Q(\core_pipeline.decode_to_execute_ecause[0] ));
 sky130_fd_sc_hd__dfxtp_1 _13811_ (.CLK(clknet_leaf_255_clk),
    .D(_00436_),
    .Q(\core_pipeline.pipeline_registers.registers[10][0] ));
 sky130_fd_sc_hd__dfxtp_1 _13812_ (.CLK(clknet_leaf_160_clk),
    .D(_00437_),
    .Q(\core_pipeline.pipeline_registers.registers[10][1] ));
 sky130_fd_sc_hd__dfxtp_1 _13813_ (.CLK(clknet_leaf_200_clk),
    .D(_00438_),
    .Q(\core_pipeline.pipeline_registers.registers[10][2] ));
 sky130_fd_sc_hd__dfxtp_1 _13814_ (.CLK(clknet_leaf_246_clk),
    .D(_00439_),
    .Q(\core_pipeline.pipeline_registers.registers[10][3] ));
 sky130_fd_sc_hd__dfxtp_1 _13815_ (.CLK(clknet_leaf_256_clk),
    .D(_00440_),
    .Q(\core_pipeline.pipeline_registers.registers[10][4] ));
 sky130_fd_sc_hd__dfxtp_1 _13816_ (.CLK(clknet_leaf_200_clk),
    .D(_00441_),
    .Q(\core_pipeline.pipeline_registers.registers[10][5] ));
 sky130_fd_sc_hd__dfxtp_1 _13817_ (.CLK(clknet_leaf_240_clk),
    .D(_00442_),
    .Q(\core_pipeline.pipeline_registers.registers[10][6] ));
 sky130_fd_sc_hd__dfxtp_1 _13818_ (.CLK(clknet_leaf_2_clk),
    .D(_00443_),
    .Q(\core_pipeline.pipeline_registers.registers[10][7] ));
 sky130_fd_sc_hd__dfxtp_1 _13819_ (.CLK(clknet_leaf_240_clk),
    .D(_00444_),
    .Q(\core_pipeline.pipeline_registers.registers[10][8] ));
 sky130_fd_sc_hd__dfxtp_1 _13820_ (.CLK(clknet_leaf_11_clk),
    .D(_00445_),
    .Q(\core_pipeline.pipeline_registers.registers[10][9] ));
 sky130_fd_sc_hd__dfxtp_1 _13821_ (.CLK(clknet_leaf_14_clk),
    .D(_00446_),
    .Q(\core_pipeline.pipeline_registers.registers[10][10] ));
 sky130_fd_sc_hd__dfxtp_1 _13822_ (.CLK(clknet_leaf_2_clk),
    .D(_00447_),
    .Q(\core_pipeline.pipeline_registers.registers[10][11] ));
 sky130_fd_sc_hd__dfxtp_1 _13823_ (.CLK(clknet_leaf_248_clk),
    .D(_00448_),
    .Q(\core_pipeline.pipeline_registers.registers[10][12] ));
 sky130_fd_sc_hd__dfxtp_1 _13824_ (.CLK(clknet_leaf_11_clk),
    .D(_00449_),
    .Q(\core_pipeline.pipeline_registers.registers[10][13] ));
 sky130_fd_sc_hd__dfxtp_1 _13825_ (.CLK(clknet_leaf_14_clk),
    .D(_00450_),
    .Q(\core_pipeline.pipeline_registers.registers[10][14] ));
 sky130_fd_sc_hd__dfxtp_1 _13826_ (.CLK(clknet_leaf_46_clk),
    .D(_00451_),
    .Q(\core_pipeline.pipeline_registers.registers[10][15] ));
 sky130_fd_sc_hd__dfxtp_1 _13827_ (.CLK(clknet_leaf_252_clk),
    .D(_00452_),
    .Q(\core_pipeline.pipeline_registers.registers[10][16] ));
 sky130_fd_sc_hd__dfxtp_1 _13828_ (.CLK(clknet_leaf_196_clk),
    .D(_00453_),
    .Q(\core_pipeline.pipeline_registers.registers[10][17] ));
 sky130_fd_sc_hd__dfxtp_1 _13829_ (.CLK(clknet_leaf_186_clk),
    .D(_00454_),
    .Q(\core_pipeline.pipeline_registers.registers[10][18] ));
 sky130_fd_sc_hd__dfxtp_1 _13830_ (.CLK(clknet_leaf_191_clk),
    .D(_00455_),
    .Q(\core_pipeline.pipeline_registers.registers[10][19] ));
 sky130_fd_sc_hd__dfxtp_1 _13831_ (.CLK(clknet_leaf_189_clk),
    .D(_00456_),
    .Q(\core_pipeline.pipeline_registers.registers[10][20] ));
 sky130_fd_sc_hd__dfxtp_1 _13832_ (.CLK(clknet_leaf_169_clk),
    .D(_00457_),
    .Q(\core_pipeline.pipeline_registers.registers[10][21] ));
 sky130_fd_sc_hd__dfxtp_1 _13833_ (.CLK(clknet_leaf_204_clk),
    .D(_00458_),
    .Q(\core_pipeline.pipeline_registers.registers[10][22] ));
 sky130_fd_sc_hd__dfxtp_1 _13834_ (.CLK(clknet_leaf_225_clk),
    .D(_00459_),
    .Q(\core_pipeline.pipeline_registers.registers[10][23] ));
 sky130_fd_sc_hd__dfxtp_1 _13835_ (.CLK(clknet_leaf_235_clk),
    .D(_00460_),
    .Q(\core_pipeline.pipeline_registers.registers[10][24] ));
 sky130_fd_sc_hd__dfxtp_1 _13836_ (.CLK(clknet_leaf_12_clk),
    .D(_00461_),
    .Q(\core_pipeline.pipeline_registers.registers[10][25] ));
 sky130_fd_sc_hd__dfxtp_1 _13837_ (.CLK(clknet_leaf_17_clk),
    .D(_00462_),
    .Q(\core_pipeline.pipeline_registers.registers[10][26] ));
 sky130_fd_sc_hd__dfxtp_1 _13838_ (.CLK(clknet_leaf_170_clk),
    .D(_00463_),
    .Q(\core_pipeline.pipeline_registers.registers[10][27] ));
 sky130_fd_sc_hd__dfxtp_1 _13839_ (.CLK(clknet_leaf_183_clk),
    .D(_00464_),
    .Q(\core_pipeline.pipeline_registers.registers[10][28] ));
 sky130_fd_sc_hd__dfxtp_1 _13840_ (.CLK(clknet_leaf_214_clk),
    .D(_00465_),
    .Q(\core_pipeline.pipeline_registers.registers[10][29] ));
 sky130_fd_sc_hd__dfxtp_1 _13841_ (.CLK(clknet_leaf_236_clk),
    .D(_00466_),
    .Q(\core_pipeline.pipeline_registers.registers[10][30] ));
 sky130_fd_sc_hd__dfxtp_1 _13842_ (.CLK(clknet_leaf_176_clk),
    .D(_00467_),
    .Q(\core_pipeline.pipeline_registers.registers[10][31] ));
 sky130_fd_sc_hd__dfxtp_1 _13843_ (.CLK(clknet_leaf_254_clk),
    .D(_00468_),
    .Q(\core_pipeline.pipeline_registers.registers[2][0] ));
 sky130_fd_sc_hd__dfxtp_1 _13844_ (.CLK(clknet_leaf_160_clk),
    .D(_00469_),
    .Q(\core_pipeline.pipeline_registers.registers[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 _13845_ (.CLK(clknet_leaf_197_clk),
    .D(_00470_),
    .Q(\core_pipeline.pipeline_registers.registers[2][2] ));
 sky130_fd_sc_hd__dfxtp_1 _13846_ (.CLK(clknet_leaf_238_clk),
    .D(_00471_),
    .Q(\core_pipeline.pipeline_registers.registers[2][3] ));
 sky130_fd_sc_hd__dfxtp_1 _13847_ (.CLK(clknet_leaf_256_clk),
    .D(_00472_),
    .Q(\core_pipeline.pipeline_registers.registers[2][4] ));
 sky130_fd_sc_hd__dfxtp_1 _13848_ (.CLK(clknet_leaf_199_clk),
    .D(_00473_),
    .Q(\core_pipeline.pipeline_registers.registers[2][5] ));
 sky130_fd_sc_hd__dfxtp_1 _13849_ (.CLK(clknet_leaf_239_clk),
    .D(_00474_),
    .Q(\core_pipeline.pipeline_registers.registers[2][6] ));
 sky130_fd_sc_hd__dfxtp_1 _13850_ (.CLK(clknet_leaf_1_clk),
    .D(_00475_),
    .Q(\core_pipeline.pipeline_registers.registers[2][7] ));
 sky130_fd_sc_hd__dfxtp_1 _13851_ (.CLK(clknet_leaf_242_clk),
    .D(_00476_),
    .Q(\core_pipeline.pipeline_registers.registers[2][8] ));
 sky130_fd_sc_hd__dfxtp_1 _13852_ (.CLK(clknet_leaf_3_clk),
    .D(_00477_),
    .Q(\core_pipeline.pipeline_registers.registers[2][9] ));
 sky130_fd_sc_hd__dfxtp_1 _13853_ (.CLK(clknet_leaf_49_clk),
    .D(_00478_),
    .Q(\core_pipeline.pipeline_registers.registers[2][10] ));
 sky130_fd_sc_hd__dfxtp_1 _13854_ (.CLK(clknet_leaf_4_clk),
    .D(_00479_),
    .Q(\core_pipeline.pipeline_registers.registers[2][11] ));
 sky130_fd_sc_hd__dfxtp_1 _13855_ (.CLK(clknet_leaf_231_clk),
    .D(_00480_),
    .Q(\core_pipeline.pipeline_registers.registers[2][12] ));
 sky130_fd_sc_hd__dfxtp_1 _13856_ (.CLK(clknet_leaf_16_clk),
    .D(_00481_),
    .Q(\core_pipeline.pipeline_registers.registers[2][13] ));
 sky130_fd_sc_hd__dfxtp_1 _13857_ (.CLK(clknet_leaf_49_clk),
    .D(_00482_),
    .Q(\core_pipeline.pipeline_registers.registers[2][14] ));
 sky130_fd_sc_hd__dfxtp_1 _13858_ (.CLK(clknet_leaf_19_clk),
    .D(_00483_),
    .Q(\core_pipeline.pipeline_registers.registers[2][15] ));
 sky130_fd_sc_hd__dfxtp_1 _13859_ (.CLK(clknet_leaf_251_clk),
    .D(_00484_),
    .Q(\core_pipeline.pipeline_registers.registers[2][16] ));
 sky130_fd_sc_hd__dfxtp_1 _13860_ (.CLK(clknet_leaf_196_clk),
    .D(_00485_),
    .Q(\core_pipeline.pipeline_registers.registers[2][17] ));
 sky130_fd_sc_hd__dfxtp_1 _13861_ (.CLK(clknet_leaf_175_clk),
    .D(_00486_),
    .Q(\core_pipeline.pipeline_registers.registers[2][18] ));
 sky130_fd_sc_hd__dfxtp_1 _13862_ (.CLK(clknet_leaf_192_clk),
    .D(_00487_),
    .Q(\core_pipeline.pipeline_registers.registers[2][19] ));
 sky130_fd_sc_hd__dfxtp_1 _13863_ (.CLK(clknet_leaf_187_clk),
    .D(_00488_),
    .Q(\core_pipeline.pipeline_registers.registers[2][20] ));
 sky130_fd_sc_hd__dfxtp_1 _13864_ (.CLK(clknet_leaf_172_clk),
    .D(_00489_),
    .Q(\core_pipeline.pipeline_registers.registers[2][21] ));
 sky130_fd_sc_hd__dfxtp_1 _13865_ (.CLK(clknet_leaf_202_clk),
    .D(_00490_),
    .Q(\core_pipeline.pipeline_registers.registers[2][22] ));
 sky130_fd_sc_hd__dfxtp_1 _13866_ (.CLK(clknet_leaf_218_clk),
    .D(_00491_),
    .Q(\core_pipeline.pipeline_registers.registers[2][23] ));
 sky130_fd_sc_hd__dfxtp_1 _13867_ (.CLK(clknet_leaf_228_clk),
    .D(_00492_),
    .Q(\core_pipeline.pipeline_registers.registers[2][24] ));
 sky130_fd_sc_hd__dfxtp_1 _13868_ (.CLK(clknet_leaf_13_clk),
    .D(_00493_),
    .Q(\core_pipeline.pipeline_registers.registers[2][25] ));
 sky130_fd_sc_hd__dfxtp_1 _13869_ (.CLK(clknet_leaf_48_clk),
    .D(_00494_),
    .Q(\core_pipeline.pipeline_registers.registers[2][26] ));
 sky130_fd_sc_hd__dfxtp_1 _13870_ (.CLK(clknet_leaf_171_clk),
    .D(_00495_),
    .Q(\core_pipeline.pipeline_registers.registers[2][27] ));
 sky130_fd_sc_hd__dfxtp_1 _13871_ (.CLK(clknet_leaf_184_clk),
    .D(_00496_),
    .Q(\core_pipeline.pipeline_registers.registers[2][28] ));
 sky130_fd_sc_hd__dfxtp_1 _13872_ (.CLK(clknet_leaf_215_clk),
    .D(_00497_),
    .Q(\core_pipeline.pipeline_registers.registers[2][29] ));
 sky130_fd_sc_hd__dfxtp_1 _13873_ (.CLK(clknet_leaf_208_clk),
    .D(_00498_),
    .Q(\core_pipeline.pipeline_registers.registers[2][30] ));
 sky130_fd_sc_hd__dfxtp_1 _13874_ (.CLK(clknet_leaf_172_clk),
    .D(_00499_),
    .Q(\core_pipeline.pipeline_registers.registers[2][31] ));
 sky130_fd_sc_hd__dfxtp_1 _13875_ (.CLK(clknet_leaf_245_clk),
    .D(_00500_),
    .Q(\core_pipeline.pipeline_registers.registers[28][0] ));
 sky130_fd_sc_hd__dfxtp_1 _13876_ (.CLK(clknet_leaf_164_clk),
    .D(_00501_),
    .Q(\core_pipeline.pipeline_registers.registers[28][1] ));
 sky130_fd_sc_hd__dfxtp_1 _13877_ (.CLK(clknet_leaf_199_clk),
    .D(_00502_),
    .Q(\core_pipeline.pipeline_registers.registers[28][2] ));
 sky130_fd_sc_hd__dfxtp_1 _13878_ (.CLK(clknet_leaf_237_clk),
    .D(_00503_),
    .Q(\core_pipeline.pipeline_registers.registers[28][3] ));
 sky130_fd_sc_hd__dfxtp_1 _13879_ (.CLK(clknet_leaf_251_clk),
    .D(_00504_),
    .Q(\core_pipeline.pipeline_registers.registers[28][4] ));
 sky130_fd_sc_hd__dfxtp_1 _13880_ (.CLK(clknet_leaf_202_clk),
    .D(_00505_),
    .Q(\core_pipeline.pipeline_registers.registers[28][5] ));
 sky130_fd_sc_hd__dfxtp_1 _13881_ (.CLK(clknet_leaf_206_clk),
    .D(_00506_),
    .Q(\core_pipeline.pipeline_registers.registers[28][6] ));
 sky130_fd_sc_hd__dfxtp_1 _13882_ (.CLK(clknet_leaf_232_clk),
    .D(_00507_),
    .Q(\core_pipeline.pipeline_registers.registers[28][7] ));
 sky130_fd_sc_hd__dfxtp_1 _13883_ (.CLK(clknet_leaf_242_clk),
    .D(_00508_),
    .Q(\core_pipeline.pipeline_registers.registers[28][8] ));
 sky130_fd_sc_hd__dfxtp_1 _13884_ (.CLK(clknet_leaf_25_clk),
    .D(_00509_),
    .Q(\core_pipeline.pipeline_registers.registers[28][9] ));
 sky130_fd_sc_hd__dfxtp_1 _13885_ (.CLK(clknet_leaf_7_clk),
    .D(_00510_),
    .Q(\core_pipeline.pipeline_registers.registers[28][10] ));
 sky130_fd_sc_hd__dfxtp_1 _13886_ (.CLK(clknet_leaf_247_clk),
    .D(_00511_),
    .Q(\core_pipeline.pipeline_registers.registers[28][11] ));
 sky130_fd_sc_hd__dfxtp_1 _13887_ (.CLK(clknet_leaf_229_clk),
    .D(_00512_),
    .Q(\core_pipeline.pipeline_registers.registers[28][12] ));
 sky130_fd_sc_hd__dfxtp_1 _13888_ (.CLK(clknet_leaf_22_clk),
    .D(_00513_),
    .Q(\core_pipeline.pipeline_registers.registers[28][13] ));
 sky130_fd_sc_hd__dfxtp_1 _13889_ (.CLK(clknet_leaf_7_clk),
    .D(_00514_),
    .Q(\core_pipeline.pipeline_registers.registers[28][14] ));
 sky130_fd_sc_hd__dfxtp_1 _13890_ (.CLK(clknet_leaf_25_clk),
    .D(_00515_),
    .Q(\core_pipeline.pipeline_registers.registers[28][15] ));
 sky130_fd_sc_hd__dfxtp_1 _13891_ (.CLK(clknet_leaf_245_clk),
    .D(_00516_),
    .Q(\core_pipeline.pipeline_registers.registers[28][16] ));
 sky130_fd_sc_hd__dfxtp_1 _13892_ (.CLK(clknet_leaf_195_clk),
    .D(_00517_),
    .Q(\core_pipeline.pipeline_registers.registers[28][17] ));
 sky130_fd_sc_hd__dfxtp_1 _13893_ (.CLK(clknet_leaf_181_clk),
    .D(_00518_),
    .Q(\core_pipeline.pipeline_registers.registers[28][18] ));
 sky130_fd_sc_hd__dfxtp_1 _13894_ (.CLK(clknet_leaf_194_clk),
    .D(_00519_),
    .Q(\core_pipeline.pipeline_registers.registers[28][19] ));
 sky130_fd_sc_hd__dfxtp_1 _13895_ (.CLK(clknet_leaf_189_clk),
    .D(_00520_),
    .Q(\core_pipeline.pipeline_registers.registers[28][20] ));
 sky130_fd_sc_hd__dfxtp_1 _13896_ (.CLK(clknet_leaf_177_clk),
    .D(_00521_),
    .Q(\core_pipeline.pipeline_registers.registers[28][21] ));
 sky130_fd_sc_hd__dfxtp_1 _13897_ (.CLK(clknet_leaf_211_clk),
    .D(_00522_),
    .Q(\core_pipeline.pipeline_registers.registers[28][22] ));
 sky130_fd_sc_hd__dfxtp_1 _13898_ (.CLK(clknet_leaf_216_clk),
    .D(_00523_),
    .Q(\core_pipeline.pipeline_registers.registers[28][23] ));
 sky130_fd_sc_hd__dfxtp_1 _13899_ (.CLK(clknet_leaf_225_clk),
    .D(_00524_),
    .Q(\core_pipeline.pipeline_registers.registers[28][24] ));
 sky130_fd_sc_hd__dfxtp_1 _13900_ (.CLK(clknet_leaf_7_clk),
    .D(_00525_),
    .Q(\core_pipeline.pipeline_registers.registers[28][25] ));
 sky130_fd_sc_hd__dfxtp_1 _13901_ (.CLK(clknet_leaf_21_clk),
    .D(_00526_),
    .Q(\core_pipeline.pipeline_registers.registers[28][26] ));
 sky130_fd_sc_hd__dfxtp_1 _13902_ (.CLK(clknet_leaf_169_clk),
    .D(_00527_),
    .Q(\core_pipeline.pipeline_registers.registers[28][27] ));
 sky130_fd_sc_hd__dfxtp_1 _13903_ (.CLK(clknet_leaf_182_clk),
    .D(_00528_),
    .Q(\core_pipeline.pipeline_registers.registers[28][28] ));
 sky130_fd_sc_hd__dfxtp_1 _13904_ (.CLK(clknet_leaf_212_clk),
    .D(_00529_),
    .Q(\core_pipeline.pipeline_registers.registers[28][29] ));
 sky130_fd_sc_hd__dfxtp_1 _13905_ (.CLK(clknet_leaf_208_clk),
    .D(_00530_),
    .Q(\core_pipeline.pipeline_registers.registers[28][30] ));
 sky130_fd_sc_hd__dfxtp_1 _13906_ (.CLK(clknet_leaf_176_clk),
    .D(_00531_),
    .Q(\core_pipeline.pipeline_registers.registers[28][31] ));
 sky130_fd_sc_hd__dfxtp_1 _13907_ (.CLK(clknet_leaf_20_clk),
    .D(_00532_),
    .Q(\core_pipeline.decode_to_execute_rs2_data[0] ));
 sky130_fd_sc_hd__dfxtp_1 _13908_ (.CLK(clknet_leaf_221_clk),
    .D(_00533_),
    .Q(\core_pipeline.decode_to_execute_rs2_data[1] ));
 sky130_fd_sc_hd__dfxtp_1 _13909_ (.CLK(clknet_leaf_220_clk),
    .D(_00534_),
    .Q(\core_pipeline.decode_to_execute_rs2_data[2] ));
 sky130_fd_sc_hd__dfxtp_1 _13910_ (.CLK(clknet_leaf_26_clk),
    .D(_00535_),
    .Q(\core_pipeline.decode_to_execute_rs2_data[3] ));
 sky130_fd_sc_hd__dfxtp_1 _13911_ (.CLK(clknet_leaf_28_clk),
    .D(_00536_),
    .Q(\core_pipeline.decode_to_execute_rs2_data[4] ));
 sky130_fd_sc_hd__dfxtp_1 _13912_ (.CLK(clknet_leaf_221_clk),
    .D(_00537_),
    .Q(\core_pipeline.decode_to_execute_rs2_data[5] ));
 sky130_fd_sc_hd__dfxtp_1 _13913_ (.CLK(clknet_leaf_225_clk),
    .D(_00538_),
    .Q(\core_pipeline.decode_to_execute_rs2_data[6] ));
 sky130_fd_sc_hd__dfxtp_1 _13914_ (.CLK(clknet_leaf_30_clk),
    .D(_00539_),
    .Q(\core_pipeline.decode_to_execute_rs2_data[7] ));
 sky130_fd_sc_hd__dfxtp_1 _13915_ (.CLK(clknet_leaf_228_clk),
    .D(_00540_),
    .Q(\core_pipeline.decode_to_execute_rs2_data[8] ));
 sky130_fd_sc_hd__dfxtp_1 _13916_ (.CLK(clknet_leaf_26_clk),
    .D(_00541_),
    .Q(\core_pipeline.decode_to_execute_rs2_data[9] ));
 sky130_fd_sc_hd__dfxtp_1 _13917_ (.CLK(clknet_leaf_28_clk),
    .D(_00542_),
    .Q(\core_pipeline.decode_to_execute_rs2_data[10] ));
 sky130_fd_sc_hd__dfxtp_1 _13918_ (.CLK(clknet_leaf_28_clk),
    .D(_00543_),
    .Q(\core_pipeline.decode_to_execute_rs2_data[11] ));
 sky130_fd_sc_hd__dfxtp_2 _13919_ (.CLK(clknet_leaf_27_clk),
    .D(_00544_),
    .Q(\core_pipeline.decode_to_execute_rs2_data[12] ));
 sky130_fd_sc_hd__dfxtp_1 _13920_ (.CLK(clknet_leaf_19_clk),
    .D(_00545_),
    .Q(\core_pipeline.decode_to_execute_rs2_data[13] ));
 sky130_fd_sc_hd__dfxtp_1 _13921_ (.CLK(clknet_leaf_26_clk),
    .D(_00546_),
    .Q(\core_pipeline.decode_to_execute_rs2_data[14] ));
 sky130_fd_sc_hd__dfxtp_1 _13922_ (.CLK(clknet_leaf_20_clk),
    .D(_00547_),
    .Q(\core_pipeline.decode_to_execute_rs2_data[15] ));
 sky130_fd_sc_hd__dfxtp_2 _13923_ (.CLK(clknet_leaf_246_clk),
    .D(_00548_),
    .Q(\core_pipeline.decode_to_execute_rs2_data[16] ));
 sky130_fd_sc_hd__dfxtp_2 _13924_ (.CLK(clknet_leaf_213_clk),
    .D(_00549_),
    .Q(\core_pipeline.decode_to_execute_rs2_data[17] ));
 sky130_fd_sc_hd__dfxtp_2 _13925_ (.CLK(clknet_leaf_180_clk),
    .D(_00550_),
    .Q(\core_pipeline.decode_to_execute_rs2_data[18] ));
 sky130_fd_sc_hd__dfxtp_2 _13926_ (.CLK(clknet_leaf_164_clk),
    .D(_00551_),
    .Q(\core_pipeline.decode_to_execute_rs2_data[19] ));
 sky130_fd_sc_hd__dfxtp_4 _13927_ (.CLK(clknet_leaf_179_clk),
    .D(_00552_),
    .Q(\core_pipeline.decode_to_execute_rs2_data[20] ));
 sky130_fd_sc_hd__dfxtp_2 _13928_ (.CLK(clknet_leaf_170_clk),
    .D(_00553_),
    .Q(\core_pipeline.decode_to_execute_rs2_data[21] ));
 sky130_fd_sc_hd__dfxtp_2 _13929_ (.CLK(clknet_leaf_210_clk),
    .D(_00554_),
    .Q(\core_pipeline.decode_to_execute_rs2_data[22] ));
 sky130_fd_sc_hd__dfxtp_1 _13930_ (.CLK(clknet_leaf_219_clk),
    .D(_00555_),
    .Q(\core_pipeline.decode_to_execute_rs2_data[23] ));
 sky130_fd_sc_hd__dfxtp_1 _13931_ (.CLK(clknet_leaf_227_clk),
    .D(_00556_),
    .Q(\core_pipeline.decode_to_execute_rs2_data[24] ));
 sky130_fd_sc_hd__dfxtp_2 _13932_ (.CLK(clknet_leaf_21_clk),
    .D(_00557_),
    .Q(\core_pipeline.decode_to_execute_rs2_data[25] ));
 sky130_fd_sc_hd__dfxtp_1 _13933_ (.CLK(clknet_leaf_21_clk),
    .D(_00558_),
    .Q(\core_pipeline.decode_to_execute_rs2_data[26] ));
 sky130_fd_sc_hd__dfxtp_2 _13934_ (.CLK(clknet_leaf_168_clk),
    .D(_00559_),
    .Q(\core_pipeline.decode_to_execute_rs2_data[27] ));
 sky130_fd_sc_hd__dfxtp_2 _13935_ (.CLK(clknet_leaf_176_clk),
    .D(_00560_),
    .Q(\core_pipeline.decode_to_execute_rs2_data[28] ));
 sky130_fd_sc_hd__dfxtp_1 _13936_ (.CLK(clknet_leaf_215_clk),
    .D(_00561_),
    .Q(\core_pipeline.decode_to_execute_rs2_data[29] ));
 sky130_fd_sc_hd__dfxtp_1 _13937_ (.CLK(clknet_leaf_225_clk),
    .D(_00562_),
    .Q(\core_pipeline.decode_to_execute_rs2_data[30] ));
 sky130_fd_sc_hd__dfxtp_1 _13938_ (.CLK(clknet_leaf_161_clk),
    .D(_00563_),
    .Q(\core_pipeline.decode_to_execute_rs2_data[31] ));
 sky130_fd_sc_hd__dfxtp_1 _13939_ (.CLK(clknet_leaf_245_clk),
    .D(_00564_),
    .Q(\core_pipeline.pipeline_registers.registers[30][0] ));
 sky130_fd_sc_hd__dfxtp_1 _13940_ (.CLK(clknet_leaf_164_clk),
    .D(_00565_),
    .Q(\core_pipeline.pipeline_registers.registers[30][1] ));
 sky130_fd_sc_hd__dfxtp_1 _13941_ (.CLK(clknet_leaf_193_clk),
    .D(_00566_),
    .Q(\core_pipeline.pipeline_registers.registers[30][2] ));
 sky130_fd_sc_hd__dfxtp_1 _13942_ (.CLK(clknet_leaf_237_clk),
    .D(_00567_),
    .Q(\core_pipeline.pipeline_registers.registers[30][3] ));
 sky130_fd_sc_hd__dfxtp_1 _13943_ (.CLK(clknet_leaf_245_clk),
    .D(_00568_),
    .Q(\core_pipeline.pipeline_registers.registers[30][4] ));
 sky130_fd_sc_hd__dfxtp_1 _13944_ (.CLK(clknet_leaf_202_clk),
    .D(_00569_),
    .Q(\core_pipeline.pipeline_registers.registers[30][5] ));
 sky130_fd_sc_hd__dfxtp_1 _13945_ (.CLK(clknet_leaf_205_clk),
    .D(_00570_),
    .Q(\core_pipeline.pipeline_registers.registers[30][6] ));
 sky130_fd_sc_hd__dfxtp_1 _13946_ (.CLK(clknet_leaf_235_clk),
    .D(_00571_),
    .Q(\core_pipeline.pipeline_registers.registers[30][7] ));
 sky130_fd_sc_hd__dfxtp_1 _13947_ (.CLK(clknet_leaf_242_clk),
    .D(_00572_),
    .Q(\core_pipeline.pipeline_registers.registers[30][8] ));
 sky130_fd_sc_hd__dfxtp_1 _13948_ (.CLK(clknet_leaf_231_clk),
    .D(_00573_),
    .Q(\core_pipeline.pipeline_registers.registers[30][9] ));
 sky130_fd_sc_hd__dfxtp_1 _13949_ (.CLK(clknet_leaf_22_clk),
    .D(_00574_),
    .Q(\core_pipeline.pipeline_registers.registers[30][10] ));
 sky130_fd_sc_hd__dfxtp_1 _13950_ (.CLK(clknet_leaf_246_clk),
    .D(_00575_),
    .Q(\core_pipeline.pipeline_registers.registers[30][11] ));
 sky130_fd_sc_hd__dfxtp_1 _13951_ (.CLK(clknet_leaf_229_clk),
    .D(_00576_),
    .Q(\core_pipeline.pipeline_registers.registers[30][12] ));
 sky130_fd_sc_hd__dfxtp_1 _13952_ (.CLK(clknet_leaf_21_clk),
    .D(_00577_),
    .Q(\core_pipeline.pipeline_registers.registers[30][13] ));
 sky130_fd_sc_hd__dfxtp_1 _13953_ (.CLK(clknet_leaf_6_clk),
    .D(_00578_),
    .Q(\core_pipeline.pipeline_registers.registers[30][14] ));
 sky130_fd_sc_hd__dfxtp_1 _13954_ (.CLK(clknet_leaf_26_clk),
    .D(_00579_),
    .Q(\core_pipeline.pipeline_registers.registers[30][15] ));
 sky130_fd_sc_hd__dfxtp_1 _13955_ (.CLK(clknet_leaf_242_clk),
    .D(_00580_),
    .Q(\core_pipeline.pipeline_registers.registers[30][16] ));
 sky130_fd_sc_hd__dfxtp_1 _13956_ (.CLK(clknet_leaf_196_clk),
    .D(_00581_),
    .Q(\core_pipeline.pipeline_registers.registers[30][17] ));
 sky130_fd_sc_hd__dfxtp_1 _13957_ (.CLK(clknet_leaf_181_clk),
    .D(_00582_),
    .Q(\core_pipeline.pipeline_registers.registers[30][18] ));
 sky130_fd_sc_hd__dfxtp_1 _13958_ (.CLK(clknet_leaf_194_clk),
    .D(_00583_),
    .Q(\core_pipeline.pipeline_registers.registers[30][19] ));
 sky130_fd_sc_hd__dfxtp_1 _13959_ (.CLK(clknet_leaf_189_clk),
    .D(_00584_),
    .Q(\core_pipeline.pipeline_registers.registers[30][20] ));
 sky130_fd_sc_hd__dfxtp_1 _13960_ (.CLK(clknet_leaf_173_clk),
    .D(_00585_),
    .Q(\core_pipeline.pipeline_registers.registers[30][21] ));
 sky130_fd_sc_hd__dfxtp_1 _13961_ (.CLK(clknet_leaf_197_clk),
    .D(_00586_),
    .Q(\core_pipeline.pipeline_registers.registers[30][22] ));
 sky130_fd_sc_hd__dfxtp_1 _13962_ (.CLK(clknet_leaf_217_clk),
    .D(_00587_),
    .Q(\core_pipeline.pipeline_registers.registers[30][23] ));
 sky130_fd_sc_hd__dfxtp_1 _13963_ (.CLK(clknet_leaf_225_clk),
    .D(_00588_),
    .Q(\core_pipeline.pipeline_registers.registers[30][24] ));
 sky130_fd_sc_hd__dfxtp_1 _13964_ (.CLK(clknet_leaf_24_clk),
    .D(_00589_),
    .Q(\core_pipeline.pipeline_registers.registers[30][25] ));
 sky130_fd_sc_hd__dfxtp_1 _13965_ (.CLK(clknet_leaf_24_clk),
    .D(_00590_),
    .Q(\core_pipeline.pipeline_registers.registers[30][26] ));
 sky130_fd_sc_hd__dfxtp_1 _13966_ (.CLK(clknet_leaf_165_clk),
    .D(_00591_),
    .Q(\core_pipeline.pipeline_registers.registers[30][27] ));
 sky130_fd_sc_hd__dfxtp_1 _13967_ (.CLK(clknet_leaf_183_clk),
    .D(_00592_),
    .Q(\core_pipeline.pipeline_registers.registers[30][28] ));
 sky130_fd_sc_hd__dfxtp_1 _13968_ (.CLK(clknet_leaf_197_clk),
    .D(_00593_),
    .Q(\core_pipeline.pipeline_registers.registers[30][29] ));
 sky130_fd_sc_hd__dfxtp_1 _13969_ (.CLK(clknet_leaf_207_clk),
    .D(_00594_),
    .Q(\core_pipeline.pipeline_registers.registers[30][30] ));
 sky130_fd_sc_hd__dfxtp_1 _13970_ (.CLK(clknet_leaf_175_clk),
    .D(_00595_),
    .Q(\core_pipeline.pipeline_registers.registers[30][31] ));
 sky130_fd_sc_hd__dfxtp_1 _13971_ (.CLK(clknet_leaf_244_clk),
    .D(_00596_),
    .Q(\core_pipeline.pipeline_registers.registers[27][0] ));
 sky130_fd_sc_hd__dfxtp_1 _13972_ (.CLK(clknet_leaf_163_clk),
    .D(_00597_),
    .Q(\core_pipeline.pipeline_registers.registers[27][1] ));
 sky130_fd_sc_hd__dfxtp_1 _13973_ (.CLK(clknet_leaf_200_clk),
    .D(_00598_),
    .Q(\core_pipeline.pipeline_registers.registers[27][2] ));
 sky130_fd_sc_hd__dfxtp_1 _13974_ (.CLK(clknet_leaf_239_clk),
    .D(_00599_),
    .Q(\core_pipeline.pipeline_registers.registers[27][3] ));
 sky130_fd_sc_hd__dfxtp_1 _13975_ (.CLK(clknet_leaf_249_clk),
    .D(_00600_),
    .Q(\core_pipeline.pipeline_registers.registers[27][4] ));
 sky130_fd_sc_hd__dfxtp_1 _13976_ (.CLK(clknet_leaf_201_clk),
    .D(_00601_),
    .Q(\core_pipeline.pipeline_registers.registers[27][5] ));
 sky130_fd_sc_hd__dfxtp_1 _13977_ (.CLK(clknet_leaf_204_clk),
    .D(_00602_),
    .Q(\core_pipeline.pipeline_registers.registers[27][6] ));
 sky130_fd_sc_hd__dfxtp_1 _13978_ (.CLK(clknet_leaf_234_clk),
    .D(_00603_),
    .Q(\core_pipeline.pipeline_registers.registers[27][7] ));
 sky130_fd_sc_hd__dfxtp_1 _13979_ (.CLK(clknet_leaf_243_clk),
    .D(_00604_),
    .Q(\core_pipeline.pipeline_registers.registers[27][8] ));
 sky130_fd_sc_hd__dfxtp_1 _13980_ (.CLK(clknet_leaf_7_clk),
    .D(_00605_),
    .Q(\core_pipeline.pipeline_registers.registers[27][9] ));
 sky130_fd_sc_hd__dfxtp_1 _13981_ (.CLK(clknet_leaf_8_clk),
    .D(_00606_),
    .Q(\core_pipeline.pipeline_registers.registers[27][10] ));
 sky130_fd_sc_hd__dfxtp_1 _13982_ (.CLK(clknet_leaf_247_clk),
    .D(_00607_),
    .Q(\core_pipeline.pipeline_registers.registers[27][11] ));
 sky130_fd_sc_hd__dfxtp_1 _13983_ (.CLK(clknet_leaf_228_clk),
    .D(_00608_),
    .Q(\core_pipeline.pipeline_registers.registers[27][12] ));
 sky130_fd_sc_hd__dfxtp_1 _13984_ (.CLK(clknet_leaf_9_clk),
    .D(_00609_),
    .Q(\core_pipeline.pipeline_registers.registers[27][13] ));
 sky130_fd_sc_hd__dfxtp_1 _13985_ (.CLK(clknet_leaf_6_clk),
    .D(_00610_),
    .Q(\core_pipeline.pipeline_registers.registers[27][14] ));
 sky130_fd_sc_hd__dfxtp_1 _13986_ (.CLK(clknet_leaf_25_clk),
    .D(_00611_),
    .Q(\core_pipeline.pipeline_registers.registers[27][15] ));
 sky130_fd_sc_hd__dfxtp_1 _13987_ (.CLK(clknet_leaf_243_clk),
    .D(_00612_),
    .Q(\core_pipeline.pipeline_registers.registers[27][16] ));
 sky130_fd_sc_hd__dfxtp_1 _13988_ (.CLK(clknet_leaf_197_clk),
    .D(_00613_),
    .Q(\core_pipeline.pipeline_registers.registers[27][17] ));
 sky130_fd_sc_hd__dfxtp_1 _13989_ (.CLK(clknet_leaf_181_clk),
    .D(_00614_),
    .Q(\core_pipeline.pipeline_registers.registers[27][18] ));
 sky130_fd_sc_hd__dfxtp_1 _13990_ (.CLK(clknet_leaf_194_clk),
    .D(_00615_),
    .Q(\core_pipeline.pipeline_registers.registers[27][19] ));
 sky130_fd_sc_hd__dfxtp_1 _13991_ (.CLK(clknet_leaf_189_clk),
    .D(_00616_),
    .Q(\core_pipeline.pipeline_registers.registers[27][20] ));
 sky130_fd_sc_hd__dfxtp_1 _13992_ (.CLK(clknet_leaf_165_clk),
    .D(_00617_),
    .Q(\core_pipeline.pipeline_registers.registers[27][21] ));
 sky130_fd_sc_hd__dfxtp_1 _13993_ (.CLK(clknet_leaf_198_clk),
    .D(_00618_),
    .Q(\core_pipeline.pipeline_registers.registers[27][22] ));
 sky130_fd_sc_hd__dfxtp_1 _13994_ (.CLK(clknet_leaf_214_clk),
    .D(_00619_),
    .Q(\core_pipeline.pipeline_registers.registers[27][23] ));
 sky130_fd_sc_hd__dfxtp_1 _13995_ (.CLK(clknet_leaf_226_clk),
    .D(_00620_),
    .Q(\core_pipeline.pipeline_registers.registers[27][24] ));
 sky130_fd_sc_hd__dfxtp_1 _13996_ (.CLK(clknet_leaf_24_clk),
    .D(_00621_),
    .Q(\core_pipeline.pipeline_registers.registers[27][25] ));
 sky130_fd_sc_hd__dfxtp_1 _13997_ (.CLK(clknet_leaf_25_clk),
    .D(_00622_),
    .Q(\core_pipeline.pipeline_registers.registers[27][26] ));
 sky130_fd_sc_hd__dfxtp_1 _13998_ (.CLK(clknet_leaf_165_clk),
    .D(_00623_),
    .Q(\core_pipeline.pipeline_registers.registers[27][27] ));
 sky130_fd_sc_hd__dfxtp_1 _13999_ (.CLK(clknet_leaf_182_clk),
    .D(_00624_),
    .Q(\core_pipeline.pipeline_registers.registers[27][28] ));
 sky130_fd_sc_hd__dfxtp_1 _14000_ (.CLK(clknet_leaf_211_clk),
    .D(_00625_),
    .Q(\core_pipeline.pipeline_registers.registers[27][29] ));
 sky130_fd_sc_hd__dfxtp_1 _14001_ (.CLK(clknet_leaf_208_clk),
    .D(_00626_),
    .Q(\core_pipeline.pipeline_registers.registers[27][30] ));
 sky130_fd_sc_hd__dfxtp_1 _14002_ (.CLK(clknet_leaf_178_clk),
    .D(_00627_),
    .Q(\core_pipeline.pipeline_registers.registers[27][31] ));
 sky130_fd_sc_hd__dfxtp_1 _14003_ (.CLK(clknet_leaf_244_clk),
    .D(_00628_),
    .Q(\core_pipeline.pipeline_registers.registers[26][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14004_ (.CLK(clknet_leaf_163_clk),
    .D(_00629_),
    .Q(\core_pipeline.pipeline_registers.registers[26][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14005_ (.CLK(clknet_leaf_200_clk),
    .D(_00630_),
    .Q(\core_pipeline.pipeline_registers.registers[26][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14006_ (.CLK(clknet_leaf_239_clk),
    .D(_00631_),
    .Q(\core_pipeline.pipeline_registers.registers[26][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14007_ (.CLK(clknet_leaf_249_clk),
    .D(_00632_),
    .Q(\core_pipeline.pipeline_registers.registers[26][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14008_ (.CLK(clknet_leaf_201_clk),
    .D(_00633_),
    .Q(\core_pipeline.pipeline_registers.registers[26][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14009_ (.CLK(clknet_leaf_204_clk),
    .D(_00634_),
    .Q(\core_pipeline.pipeline_registers.registers[26][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14010_ (.CLK(clknet_leaf_234_clk),
    .D(_00635_),
    .Q(\core_pipeline.pipeline_registers.registers[26][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14011_ (.CLK(clknet_leaf_243_clk),
    .D(_00636_),
    .Q(\core_pipeline.pipeline_registers.registers[26][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14012_ (.CLK(clknet_leaf_7_clk),
    .D(_00637_),
    .Q(\core_pipeline.pipeline_registers.registers[26][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14013_ (.CLK(clknet_leaf_8_clk),
    .D(_00638_),
    .Q(\core_pipeline.pipeline_registers.registers[26][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14014_ (.CLK(clknet_leaf_247_clk),
    .D(_00639_),
    .Q(\core_pipeline.pipeline_registers.registers[26][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14015_ (.CLK(clknet_leaf_228_clk),
    .D(_00640_),
    .Q(\core_pipeline.pipeline_registers.registers[26][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14016_ (.CLK(clknet_leaf_8_clk),
    .D(_00641_),
    .Q(\core_pipeline.pipeline_registers.registers[26][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14017_ (.CLK(clknet_leaf_6_clk),
    .D(_00642_),
    .Q(\core_pipeline.pipeline_registers.registers[26][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14018_ (.CLK(clknet_leaf_230_clk),
    .D(_00643_),
    .Q(\core_pipeline.pipeline_registers.registers[26][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14019_ (.CLK(clknet_leaf_243_clk),
    .D(_00644_),
    .Q(\core_pipeline.pipeline_registers.registers[26][16] ));
 sky130_fd_sc_hd__dfxtp_1 _14020_ (.CLK(clknet_leaf_195_clk),
    .D(_00645_),
    .Q(\core_pipeline.pipeline_registers.registers[26][17] ));
 sky130_fd_sc_hd__dfxtp_1 _14021_ (.CLK(clknet_leaf_182_clk),
    .D(_00646_),
    .Q(\core_pipeline.pipeline_registers.registers[26][18] ));
 sky130_fd_sc_hd__dfxtp_1 _14022_ (.CLK(clknet_leaf_193_clk),
    .D(_00647_),
    .Q(\core_pipeline.pipeline_registers.registers[26][19] ));
 sky130_fd_sc_hd__dfxtp_1 _14023_ (.CLK(clknet_leaf_191_clk),
    .D(_00648_),
    .Q(\core_pipeline.pipeline_registers.registers[26][20] ));
 sky130_fd_sc_hd__dfxtp_1 _14024_ (.CLK(clknet_leaf_165_clk),
    .D(_00649_),
    .Q(\core_pipeline.pipeline_registers.registers[26][21] ));
 sky130_fd_sc_hd__dfxtp_1 _14025_ (.CLK(clknet_leaf_198_clk),
    .D(_00650_),
    .Q(\core_pipeline.pipeline_registers.registers[26][22] ));
 sky130_fd_sc_hd__dfxtp_1 _14026_ (.CLK(clknet_leaf_214_clk),
    .D(_00651_),
    .Q(\core_pipeline.pipeline_registers.registers[26][23] ));
 sky130_fd_sc_hd__dfxtp_1 _14027_ (.CLK(clknet_leaf_236_clk),
    .D(_00652_),
    .Q(\core_pipeline.pipeline_registers.registers[26][24] ));
 sky130_fd_sc_hd__dfxtp_1 _14028_ (.CLK(clknet_leaf_24_clk),
    .D(_00653_),
    .Q(\core_pipeline.pipeline_registers.registers[26][25] ));
 sky130_fd_sc_hd__dfxtp_1 _14029_ (.CLK(clknet_leaf_25_clk),
    .D(_00654_),
    .Q(\core_pipeline.pipeline_registers.registers[26][26] ));
 sky130_fd_sc_hd__dfxtp_1 _14030_ (.CLK(clknet_leaf_165_clk),
    .D(_00655_),
    .Q(\core_pipeline.pipeline_registers.registers[26][27] ));
 sky130_fd_sc_hd__dfxtp_1 _14031_ (.CLK(clknet_leaf_194_clk),
    .D(_00656_),
    .Q(\core_pipeline.pipeline_registers.registers[26][28] ));
 sky130_fd_sc_hd__dfxtp_1 _14032_ (.CLK(clknet_leaf_212_clk),
    .D(_00657_),
    .Q(\core_pipeline.pipeline_registers.registers[26][29] ));
 sky130_fd_sc_hd__dfxtp_1 _14033_ (.CLK(clknet_leaf_208_clk),
    .D(_00658_),
    .Q(\core_pipeline.pipeline_registers.registers[26][30] ));
 sky130_fd_sc_hd__dfxtp_1 _14034_ (.CLK(clknet_leaf_178_clk),
    .D(_00659_),
    .Q(\core_pipeline.pipeline_registers.registers[26][31] ));
 sky130_fd_sc_hd__dfxtp_1 _14035_ (.CLK(clknet_leaf_244_clk),
    .D(_00660_),
    .Q(\core_pipeline.pipeline_registers.registers[25][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14036_ (.CLK(clknet_leaf_163_clk),
    .D(_00661_),
    .Q(\core_pipeline.pipeline_registers.registers[25][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14037_ (.CLK(clknet_leaf_199_clk),
    .D(_00662_),
    .Q(\core_pipeline.pipeline_registers.registers[25][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14038_ (.CLK(clknet_leaf_238_clk),
    .D(_00663_),
    .Q(\core_pipeline.pipeline_registers.registers[25][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14039_ (.CLK(clknet_leaf_251_clk),
    .D(_00664_),
    .Q(\core_pipeline.pipeline_registers.registers[25][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14040_ (.CLK(clknet_leaf_203_clk),
    .D(_00665_),
    .Q(\core_pipeline.pipeline_registers.registers[25][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14041_ (.CLK(clknet_leaf_205_clk),
    .D(_00666_),
    .Q(\core_pipeline.pipeline_registers.registers[25][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14042_ (.CLK(clknet_leaf_233_clk),
    .D(_00667_),
    .Q(\core_pipeline.pipeline_registers.registers[25][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14043_ (.CLK(clknet_leaf_243_clk),
    .D(_00668_),
    .Q(\core_pipeline.pipeline_registers.registers[25][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14044_ (.CLK(clknet_leaf_7_clk),
    .D(_00669_),
    .Q(\core_pipeline.pipeline_registers.registers[25][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14045_ (.CLK(clknet_leaf_8_clk),
    .D(_00670_),
    .Q(\core_pipeline.pipeline_registers.registers[25][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14046_ (.CLK(clknet_leaf_247_clk),
    .D(_00671_),
    .Q(\core_pipeline.pipeline_registers.registers[25][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14047_ (.CLK(clknet_leaf_232_clk),
    .D(_00672_),
    .Q(\core_pipeline.pipeline_registers.registers[25][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14048_ (.CLK(clknet_leaf_22_clk),
    .D(_00673_),
    .Q(\core_pipeline.pipeline_registers.registers[25][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14049_ (.CLK(clknet_leaf_8_clk),
    .D(_00674_),
    .Q(\core_pipeline.pipeline_registers.registers[25][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14050_ (.CLK(clknet_leaf_25_clk),
    .D(_00675_),
    .Q(\core_pipeline.pipeline_registers.registers[25][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14051_ (.CLK(clknet_leaf_243_clk),
    .D(_00676_),
    .Q(\core_pipeline.pipeline_registers.registers[25][16] ));
 sky130_fd_sc_hd__dfxtp_1 _14052_ (.CLK(clknet_leaf_197_clk),
    .D(_00677_),
    .Q(\core_pipeline.pipeline_registers.registers[25][17] ));
 sky130_fd_sc_hd__dfxtp_1 _14053_ (.CLK(clknet_leaf_196_clk),
    .D(_00678_),
    .Q(\core_pipeline.pipeline_registers.registers[25][18] ));
 sky130_fd_sc_hd__dfxtp_1 _14054_ (.CLK(clknet_leaf_193_clk),
    .D(_00679_),
    .Q(\core_pipeline.pipeline_registers.registers[25][19] ));
 sky130_fd_sc_hd__dfxtp_1 _14055_ (.CLK(clknet_leaf_191_clk),
    .D(_00680_),
    .Q(\core_pipeline.pipeline_registers.registers[25][20] ));
 sky130_fd_sc_hd__dfxtp_1 _14056_ (.CLK(clknet_leaf_165_clk),
    .D(_00681_),
    .Q(\core_pipeline.pipeline_registers.registers[25][21] ));
 sky130_fd_sc_hd__dfxtp_1 _14057_ (.CLK(clknet_leaf_198_clk),
    .D(_00682_),
    .Q(\core_pipeline.pipeline_registers.registers[25][22] ));
 sky130_fd_sc_hd__dfxtp_1 _14058_ (.CLK(clknet_leaf_217_clk),
    .D(_00683_),
    .Q(\core_pipeline.pipeline_registers.registers[25][23] ));
 sky130_fd_sc_hd__dfxtp_1 _14059_ (.CLK(clknet_leaf_226_clk),
    .D(_00684_),
    .Q(\core_pipeline.pipeline_registers.registers[25][24] ));
 sky130_fd_sc_hd__dfxtp_1 _14060_ (.CLK(clknet_leaf_24_clk),
    .D(_00685_),
    .Q(\core_pipeline.pipeline_registers.registers[25][25] ));
 sky130_fd_sc_hd__dfxtp_1 _14061_ (.CLK(clknet_leaf_23_clk),
    .D(_00686_),
    .Q(\core_pipeline.pipeline_registers.registers[25][26] ));
 sky130_fd_sc_hd__dfxtp_1 _14062_ (.CLK(clknet_leaf_166_clk),
    .D(_00687_),
    .Q(\core_pipeline.pipeline_registers.registers[25][27] ));
 sky130_fd_sc_hd__dfxtp_1 _14063_ (.CLK(clknet_leaf_182_clk),
    .D(_00688_),
    .Q(\core_pipeline.pipeline_registers.registers[25][28] ));
 sky130_fd_sc_hd__dfxtp_1 _14064_ (.CLK(clknet_leaf_212_clk),
    .D(_00689_),
    .Q(\core_pipeline.pipeline_registers.registers[25][29] ));
 sky130_fd_sc_hd__dfxtp_1 _14065_ (.CLK(clknet_leaf_208_clk),
    .D(_00690_),
    .Q(\core_pipeline.pipeline_registers.registers[25][30] ));
 sky130_fd_sc_hd__dfxtp_1 _14066_ (.CLK(clknet_leaf_179_clk),
    .D(_00691_),
    .Q(\core_pipeline.pipeline_registers.registers[25][31] ));
 sky130_fd_sc_hd__dfxtp_1 _14067_ (.CLK(clknet_leaf_244_clk),
    .D(_00692_),
    .Q(\core_pipeline.pipeline_registers.registers[24][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14068_ (.CLK(clknet_leaf_164_clk),
    .D(_00693_),
    .Q(\core_pipeline.pipeline_registers.registers[24][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14069_ (.CLK(clknet_leaf_200_clk),
    .D(_00694_),
    .Q(\core_pipeline.pipeline_registers.registers[24][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14070_ (.CLK(clknet_leaf_238_clk),
    .D(_00695_),
    .Q(\core_pipeline.pipeline_registers.registers[24][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14071_ (.CLK(clknet_leaf_249_clk),
    .D(_00696_),
    .Q(\core_pipeline.pipeline_registers.registers[24][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14072_ (.CLK(clknet_leaf_203_clk),
    .D(_00697_),
    .Q(\core_pipeline.pipeline_registers.registers[24][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14073_ (.CLK(clknet_leaf_205_clk),
    .D(_00698_),
    .Q(\core_pipeline.pipeline_registers.registers[24][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14074_ (.CLK(clknet_leaf_234_clk),
    .D(_00699_),
    .Q(\core_pipeline.pipeline_registers.registers[24][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14075_ (.CLK(clknet_leaf_242_clk),
    .D(_00700_),
    .Q(\core_pipeline.pipeline_registers.registers[24][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14076_ (.CLK(clknet_leaf_248_clk),
    .D(_00701_),
    .Q(\core_pipeline.pipeline_registers.registers[24][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14077_ (.CLK(clknet_leaf_8_clk),
    .D(_00702_),
    .Q(\core_pipeline.pipeline_registers.registers[24][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14078_ (.CLK(clknet_leaf_249_clk),
    .D(_00703_),
    .Q(\core_pipeline.pipeline_registers.registers[24][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14079_ (.CLK(clknet_leaf_229_clk),
    .D(_00704_),
    .Q(\core_pipeline.pipeline_registers.registers[24][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14080_ (.CLK(clknet_leaf_22_clk),
    .D(_00705_),
    .Q(\core_pipeline.pipeline_registers.registers[24][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14081_ (.CLK(clknet_leaf_8_clk),
    .D(_00706_),
    .Q(\core_pipeline.pipeline_registers.registers[24][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14082_ (.CLK(clknet_leaf_25_clk),
    .D(_00707_),
    .Q(\core_pipeline.pipeline_registers.registers[24][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14083_ (.CLK(clknet_leaf_243_clk),
    .D(_00708_),
    .Q(\core_pipeline.pipeline_registers.registers[24][16] ));
 sky130_fd_sc_hd__dfxtp_1 _14084_ (.CLK(clknet_leaf_197_clk),
    .D(_00709_),
    .Q(\core_pipeline.pipeline_registers.registers[24][17] ));
 sky130_fd_sc_hd__dfxtp_1 _14085_ (.CLK(clknet_leaf_195_clk),
    .D(_00710_),
    .Q(\core_pipeline.pipeline_registers.registers[24][18] ));
 sky130_fd_sc_hd__dfxtp_1 _14086_ (.CLK(clknet_leaf_193_clk),
    .D(_00711_),
    .Q(\core_pipeline.pipeline_registers.registers[24][19] ));
 sky130_fd_sc_hd__dfxtp_1 _14087_ (.CLK(clknet_leaf_191_clk),
    .D(_00712_),
    .Q(\core_pipeline.pipeline_registers.registers[24][20] ));
 sky130_fd_sc_hd__dfxtp_1 _14088_ (.CLK(clknet_leaf_165_clk),
    .D(_00713_),
    .Q(\core_pipeline.pipeline_registers.registers[24][21] ));
 sky130_fd_sc_hd__dfxtp_1 _14089_ (.CLK(clknet_leaf_198_clk),
    .D(_00714_),
    .Q(\core_pipeline.pipeline_registers.registers[24][22] ));
 sky130_fd_sc_hd__dfxtp_1 _14090_ (.CLK(clknet_leaf_217_clk),
    .D(_00715_),
    .Q(\core_pipeline.pipeline_registers.registers[24][23] ));
 sky130_fd_sc_hd__dfxtp_1 _14091_ (.CLK(clknet_leaf_226_clk),
    .D(_00716_),
    .Q(\core_pipeline.pipeline_registers.registers[24][24] ));
 sky130_fd_sc_hd__dfxtp_1 _14092_ (.CLK(clknet_leaf_24_clk),
    .D(_00717_),
    .Q(\core_pipeline.pipeline_registers.registers[24][25] ));
 sky130_fd_sc_hd__dfxtp_1 _14093_ (.CLK(clknet_leaf_23_clk),
    .D(_00718_),
    .Q(\core_pipeline.pipeline_registers.registers[24][26] ));
 sky130_fd_sc_hd__dfxtp_1 _14094_ (.CLK(clknet_leaf_166_clk),
    .D(_00719_),
    .Q(\core_pipeline.pipeline_registers.registers[24][27] ));
 sky130_fd_sc_hd__dfxtp_1 _14095_ (.CLK(clknet_leaf_182_clk),
    .D(_00720_),
    .Q(\core_pipeline.pipeline_registers.registers[24][28] ));
 sky130_fd_sc_hd__dfxtp_1 _14096_ (.CLK(clknet_leaf_212_clk),
    .D(_00721_),
    .Q(\core_pipeline.pipeline_registers.registers[24][29] ));
 sky130_fd_sc_hd__dfxtp_1 _14097_ (.CLK(clknet_leaf_208_clk),
    .D(_00722_),
    .Q(\core_pipeline.pipeline_registers.registers[24][30] ));
 sky130_fd_sc_hd__dfxtp_1 _14098_ (.CLK(clknet_leaf_180_clk),
    .D(_00723_),
    .Q(\core_pipeline.pipeline_registers.registers[24][31] ));
 sky130_fd_sc_hd__dfxtp_1 _14099_ (.CLK(clknet_leaf_253_clk),
    .D(_00724_),
    .Q(\core_pipeline.pipeline_registers.registers[23][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14100_ (.CLK(clknet_leaf_161_clk),
    .D(_00725_),
    .Q(\core_pipeline.pipeline_registers.registers[23][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14101_ (.CLK(clknet_leaf_197_clk),
    .D(_00726_),
    .Q(\core_pipeline.pipeline_registers.registers[23][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14102_ (.CLK(clknet_leaf_234_clk),
    .D(_00727_),
    .Q(\core_pipeline.pipeline_registers.registers[23][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14103_ (.CLK(clknet_leaf_254_clk),
    .D(_00728_),
    .Q(\core_pipeline.pipeline_registers.registers[23][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14104_ (.CLK(clknet_leaf_202_clk),
    .D(_00729_),
    .Q(\core_pipeline.pipeline_registers.registers[23][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14105_ (.CLK(clknet_leaf_239_clk),
    .D(_00730_),
    .Q(\core_pipeline.pipeline_registers.registers[23][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14106_ (.CLK(clknet_leaf_233_clk),
    .D(_00731_),
    .Q(\core_pipeline.pipeline_registers.registers[23][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14107_ (.CLK(clknet_leaf_246_clk),
    .D(_00732_),
    .Q(\core_pipeline.pipeline_registers.registers[23][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14108_ (.CLK(clknet_leaf_4_clk),
    .D(_00733_),
    .Q(\core_pipeline.pipeline_registers.registers[23][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14109_ (.CLK(clknet_leaf_10_clk),
    .D(_00734_),
    .Q(\core_pipeline.pipeline_registers.registers[23][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14110_ (.CLK(clknet_leaf_249_clk),
    .D(_00735_),
    .Q(\core_pipeline.pipeline_registers.registers[23][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14111_ (.CLK(clknet_leaf_231_clk),
    .D(_00736_),
    .Q(\core_pipeline.pipeline_registers.registers[23][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14112_ (.CLK(clknet_leaf_12_clk),
    .D(_00737_),
    .Q(\core_pipeline.pipeline_registers.registers[23][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14113_ (.CLK(clknet_leaf_4_clk),
    .D(_00738_),
    .Q(\core_pipeline.pipeline_registers.registers[23][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14114_ (.CLK(clknet_leaf_21_clk),
    .D(_00739_),
    .Q(\core_pipeline.pipeline_registers.registers[23][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14115_ (.CLK(clknet_leaf_245_clk),
    .D(_00740_),
    .Q(\core_pipeline.pipeline_registers.registers[23][16] ));
 sky130_fd_sc_hd__dfxtp_1 _14116_ (.CLK(clknet_leaf_162_clk),
    .D(_00741_),
    .Q(\core_pipeline.pipeline_registers.registers[23][17] ));
 sky130_fd_sc_hd__dfxtp_1 _14117_ (.CLK(clknet_leaf_180_clk),
    .D(_00742_),
    .Q(\core_pipeline.pipeline_registers.registers[23][18] ));
 sky130_fd_sc_hd__dfxtp_1 _14118_ (.CLK(clknet_leaf_195_clk),
    .D(_00743_),
    .Q(\core_pipeline.pipeline_registers.registers[23][19] ));
 sky130_fd_sc_hd__dfxtp_1 _14119_ (.CLK(clknet_leaf_190_clk),
    .D(_00744_),
    .Q(\core_pipeline.pipeline_registers.registers[23][20] ));
 sky130_fd_sc_hd__dfxtp_1 _14120_ (.CLK(clknet_leaf_169_clk),
    .D(_00745_),
    .Q(\core_pipeline.pipeline_registers.registers[23][21] ));
 sky130_fd_sc_hd__dfxtp_1 _14121_ (.CLK(clknet_leaf_207_clk),
    .D(_00746_),
    .Q(\core_pipeline.pipeline_registers.registers[23][22] ));
 sky130_fd_sc_hd__dfxtp_1 _14122_ (.CLK(clknet_leaf_218_clk),
    .D(_00747_),
    .Q(\core_pipeline.pipeline_registers.registers[23][23] ));
 sky130_fd_sc_hd__dfxtp_1 _14123_ (.CLK(clknet_leaf_227_clk),
    .D(_00748_),
    .Q(\core_pipeline.pipeline_registers.registers[23][24] ));
 sky130_fd_sc_hd__dfxtp_1 _14124_ (.CLK(clknet_leaf_10_clk),
    .D(_00749_),
    .Q(\core_pipeline.pipeline_registers.registers[23][25] ));
 sky130_fd_sc_hd__dfxtp_1 _14125_ (.CLK(clknet_leaf_18_clk),
    .D(_00750_),
    .Q(\core_pipeline.pipeline_registers.registers[23][26] ));
 sky130_fd_sc_hd__dfxtp_1 _14126_ (.CLK(clknet_leaf_166_clk),
    .D(_00751_),
    .Q(\core_pipeline.pipeline_registers.registers[23][27] ));
 sky130_fd_sc_hd__dfxtp_1 _14127_ (.CLK(clknet_leaf_181_clk),
    .D(_00752_),
    .Q(\core_pipeline.pipeline_registers.registers[23][28] ));
 sky130_fd_sc_hd__dfxtp_1 _14128_ (.CLK(clknet_leaf_210_clk),
    .D(_00753_),
    .Q(\core_pipeline.pipeline_registers.registers[23][29] ));
 sky130_fd_sc_hd__dfxtp_1 _14129_ (.CLK(clknet_leaf_209_clk),
    .D(_00754_),
    .Q(\core_pipeline.pipeline_registers.registers[23][30] ));
 sky130_fd_sc_hd__dfxtp_1 _14130_ (.CLK(clknet_leaf_177_clk),
    .D(_00755_),
    .Q(\core_pipeline.pipeline_registers.registers[23][31] ));
 sky130_fd_sc_hd__dfxtp_1 _14131_ (.CLK(clknet_leaf_251_clk),
    .D(_00756_),
    .Q(\core_pipeline.pipeline_registers.registers[21][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14132_ (.CLK(clknet_leaf_161_clk),
    .D(_00757_),
    .Q(\core_pipeline.pipeline_registers.registers[21][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14133_ (.CLK(clknet_leaf_199_clk),
    .D(_00758_),
    .Q(\core_pipeline.pipeline_registers.registers[21][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14134_ (.CLK(clknet_leaf_237_clk),
    .D(_00759_),
    .Q(\core_pipeline.pipeline_registers.registers[21][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14135_ (.CLK(clknet_leaf_254_clk),
    .D(_00760_),
    .Q(\core_pipeline.pipeline_registers.registers[21][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14136_ (.CLK(clknet_leaf_202_clk),
    .D(_00761_),
    .Q(\core_pipeline.pipeline_registers.registers[21][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14137_ (.CLK(clknet_leaf_206_clk),
    .D(_00762_),
    .Q(\core_pipeline.pipeline_registers.registers[21][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14138_ (.CLK(clknet_leaf_233_clk),
    .D(_00763_),
    .Q(\core_pipeline.pipeline_registers.registers[21][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14139_ (.CLK(clknet_leaf_242_clk),
    .D(_00764_),
    .Q(\core_pipeline.pipeline_registers.registers[21][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14140_ (.CLK(clknet_leaf_6_clk),
    .D(_00765_),
    .Q(\core_pipeline.pipeline_registers.registers[21][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14141_ (.CLK(clknet_leaf_10_clk),
    .D(_00766_),
    .Q(\core_pipeline.pipeline_registers.registers[21][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14142_ (.CLK(clknet_leaf_249_clk),
    .D(_00767_),
    .Q(\core_pipeline.pipeline_registers.registers[21][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14143_ (.CLK(clknet_leaf_231_clk),
    .D(_00768_),
    .Q(\core_pipeline.pipeline_registers.registers[21][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14144_ (.CLK(clknet_leaf_13_clk),
    .D(_00769_),
    .Q(\core_pipeline.pipeline_registers.registers[21][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14145_ (.CLK(clknet_leaf_4_clk),
    .D(_00770_),
    .Q(\core_pipeline.pipeline_registers.registers[21][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14146_ (.CLK(clknet_leaf_20_clk),
    .D(_00771_),
    .Q(\core_pipeline.pipeline_registers.registers[21][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14147_ (.CLK(clknet_leaf_246_clk),
    .D(_00772_),
    .Q(\core_pipeline.pipeline_registers.registers[21][16] ));
 sky130_fd_sc_hd__dfxtp_1 _14148_ (.CLK(clknet_leaf_162_clk),
    .D(_00773_),
    .Q(\core_pipeline.pipeline_registers.registers[21][17] ));
 sky130_fd_sc_hd__dfxtp_1 _14149_ (.CLK(clknet_leaf_179_clk),
    .D(_00774_),
    .Q(\core_pipeline.pipeline_registers.registers[21][18] ));
 sky130_fd_sc_hd__dfxtp_1 _14150_ (.CLK(clknet_leaf_194_clk),
    .D(_00775_),
    .Q(\core_pipeline.pipeline_registers.registers[21][19] ));
 sky130_fd_sc_hd__dfxtp_1 _14151_ (.CLK(clknet_leaf_190_clk),
    .D(_00776_),
    .Q(\core_pipeline.pipeline_registers.registers[21][20] ));
 sky130_fd_sc_hd__dfxtp_1 _14152_ (.CLK(clknet_leaf_169_clk),
    .D(_00777_),
    .Q(\core_pipeline.pipeline_registers.registers[21][21] ));
 sky130_fd_sc_hd__dfxtp_1 _14153_ (.CLK(clknet_leaf_207_clk),
    .D(_00778_),
    .Q(\core_pipeline.pipeline_registers.registers[21][22] ));
 sky130_fd_sc_hd__dfxtp_1 _14154_ (.CLK(clknet_leaf_209_clk),
    .D(_00779_),
    .Q(\core_pipeline.pipeline_registers.registers[21][23] ));
 sky130_fd_sc_hd__dfxtp_1 _14155_ (.CLK(clknet_leaf_224_clk),
    .D(_00780_),
    .Q(\core_pipeline.pipeline_registers.registers[21][24] ));
 sky130_fd_sc_hd__dfxtp_1 _14156_ (.CLK(clknet_leaf_10_clk),
    .D(_00781_),
    .Q(\core_pipeline.pipeline_registers.registers[21][25] ));
 sky130_fd_sc_hd__dfxtp_1 _14157_ (.CLK(clknet_leaf_18_clk),
    .D(_00782_),
    .Q(\core_pipeline.pipeline_registers.registers[21][26] ));
 sky130_fd_sc_hd__dfxtp_1 _14158_ (.CLK(clknet_leaf_165_clk),
    .D(_00783_),
    .Q(\core_pipeline.pipeline_registers.registers[21][27] ));
 sky130_fd_sc_hd__dfxtp_1 _14159_ (.CLK(clknet_leaf_184_clk),
    .D(_00784_),
    .Q(\core_pipeline.pipeline_registers.registers[21][28] ));
 sky130_fd_sc_hd__dfxtp_1 _14160_ (.CLK(clknet_leaf_211_clk),
    .D(_00785_),
    .Q(\core_pipeline.pipeline_registers.registers[21][29] ));
 sky130_fd_sc_hd__dfxtp_1 _14161_ (.CLK(clknet_leaf_209_clk),
    .D(_00786_),
    .Q(\core_pipeline.pipeline_registers.registers[21][30] ));
 sky130_fd_sc_hd__dfxtp_1 _14162_ (.CLK(clknet_leaf_177_clk),
    .D(_00787_),
    .Q(\core_pipeline.pipeline_registers.registers[21][31] ));
 sky130_fd_sc_hd__dfxtp_1 _14163_ (.CLK(clknet_leaf_253_clk),
    .D(_00788_),
    .Q(\core_pipeline.pipeline_registers.registers[22][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14164_ (.CLK(clknet_leaf_161_clk),
    .D(_00789_),
    .Q(\core_pipeline.pipeline_registers.registers[22][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14165_ (.CLK(clknet_leaf_198_clk),
    .D(_00790_),
    .Q(\core_pipeline.pipeline_registers.registers[22][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14166_ (.CLK(clknet_leaf_234_clk),
    .D(_00791_),
    .Q(\core_pipeline.pipeline_registers.registers[22][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14167_ (.CLK(clknet_leaf_254_clk),
    .D(_00792_),
    .Q(\core_pipeline.pipeline_registers.registers[22][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14168_ (.CLK(clknet_leaf_202_clk),
    .D(_00793_),
    .Q(\core_pipeline.pipeline_registers.registers[22][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14169_ (.CLK(clknet_leaf_239_clk),
    .D(_00794_),
    .Q(\core_pipeline.pipeline_registers.registers[22][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14170_ (.CLK(clknet_leaf_246_clk),
    .D(_00795_),
    .Q(\core_pipeline.pipeline_registers.registers[22][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14171_ (.CLK(clknet_leaf_246_clk),
    .D(_00796_),
    .Q(\core_pipeline.pipeline_registers.registers[22][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14172_ (.CLK(clknet_leaf_4_clk),
    .D(_00797_),
    .Q(\core_pipeline.pipeline_registers.registers[22][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14173_ (.CLK(clknet_leaf_10_clk),
    .D(_00798_),
    .Q(\core_pipeline.pipeline_registers.registers[22][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14174_ (.CLK(clknet_leaf_249_clk),
    .D(_00799_),
    .Q(\core_pipeline.pipeline_registers.registers[22][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14175_ (.CLK(clknet_leaf_230_clk),
    .D(_00800_),
    .Q(\core_pipeline.pipeline_registers.registers[22][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14176_ (.CLK(clknet_leaf_13_clk),
    .D(_00801_),
    .Q(\core_pipeline.pipeline_registers.registers[22][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14177_ (.CLK(clknet_leaf_4_clk),
    .D(_00802_),
    .Q(\core_pipeline.pipeline_registers.registers[22][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14178_ (.CLK(clknet_leaf_21_clk),
    .D(_00803_),
    .Q(\core_pipeline.pipeline_registers.registers[22][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14179_ (.CLK(clknet_leaf_245_clk),
    .D(_00804_),
    .Q(\core_pipeline.pipeline_registers.registers[22][16] ));
 sky130_fd_sc_hd__dfxtp_1 _14180_ (.CLK(clknet_leaf_162_clk),
    .D(_00805_),
    .Q(\core_pipeline.pipeline_registers.registers[22][17] ));
 sky130_fd_sc_hd__dfxtp_1 _14181_ (.CLK(clknet_leaf_180_clk),
    .D(_00806_),
    .Q(\core_pipeline.pipeline_registers.registers[22][18] ));
 sky130_fd_sc_hd__dfxtp_1 _14182_ (.CLK(clknet_leaf_193_clk),
    .D(_00807_),
    .Q(\core_pipeline.pipeline_registers.registers[22][19] ));
 sky130_fd_sc_hd__dfxtp_1 _14183_ (.CLK(clknet_leaf_190_clk),
    .D(_00808_),
    .Q(\core_pipeline.pipeline_registers.registers[22][20] ));
 sky130_fd_sc_hd__dfxtp_1 _14184_ (.CLK(clknet_leaf_169_clk),
    .D(_00809_),
    .Q(\core_pipeline.pipeline_registers.registers[22][21] ));
 sky130_fd_sc_hd__dfxtp_1 _14185_ (.CLK(clknet_leaf_207_clk),
    .D(_00810_),
    .Q(\core_pipeline.pipeline_registers.registers[22][22] ));
 sky130_fd_sc_hd__dfxtp_1 _14186_ (.CLK(clknet_leaf_209_clk),
    .D(_00811_),
    .Q(\core_pipeline.pipeline_registers.registers[22][23] ));
 sky130_fd_sc_hd__dfxtp_1 _14187_ (.CLK(clknet_leaf_227_clk),
    .D(_00812_),
    .Q(\core_pipeline.pipeline_registers.registers[22][24] ));
 sky130_fd_sc_hd__dfxtp_1 _14188_ (.CLK(clknet_leaf_10_clk),
    .D(_00813_),
    .Q(\core_pipeline.pipeline_registers.registers[22][25] ));
 sky130_fd_sc_hd__dfxtp_1 _14189_ (.CLK(clknet_leaf_18_clk),
    .D(_00814_),
    .Q(\core_pipeline.pipeline_registers.registers[22][26] ));
 sky130_fd_sc_hd__dfxtp_1 _14190_ (.CLK(clknet_leaf_166_clk),
    .D(_00815_),
    .Q(\core_pipeline.pipeline_registers.registers[22][27] ));
 sky130_fd_sc_hd__dfxtp_1 _14191_ (.CLK(clknet_leaf_181_clk),
    .D(_00816_),
    .Q(\core_pipeline.pipeline_registers.registers[22][28] ));
 sky130_fd_sc_hd__dfxtp_1 _14192_ (.CLK(clknet_leaf_210_clk),
    .D(_00817_),
    .Q(\core_pipeline.pipeline_registers.registers[22][29] ));
 sky130_fd_sc_hd__dfxtp_1 _14193_ (.CLK(clknet_leaf_208_clk),
    .D(_00818_),
    .Q(\core_pipeline.pipeline_registers.registers[22][30] ));
 sky130_fd_sc_hd__dfxtp_1 _14194_ (.CLK(clknet_leaf_177_clk),
    .D(_00819_),
    .Q(\core_pipeline.pipeline_registers.registers[22][31] ));
 sky130_fd_sc_hd__dfxtp_2 _14195_ (.CLK(clknet_leaf_35_clk),
    .D(_00820_),
    .Q(\core_pipeline.pipeline_decode.alu_select_a_out[1] ));
 sky130_fd_sc_hd__dfxtp_1 _14196_ (.CLK(clknet_leaf_254_clk),
    .D(_00821_),
    .Q(\core_pipeline.pipeline_registers.registers[3][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14197_ (.CLK(clknet_leaf_160_clk),
    .D(_00822_),
    .Q(\core_pipeline.pipeline_registers.registers[3][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14198_ (.CLK(clknet_leaf_197_clk),
    .D(_00823_),
    .Q(\core_pipeline.pipeline_registers.registers[3][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14199_ (.CLK(clknet_leaf_238_clk),
    .D(_00824_),
    .Q(\core_pipeline.pipeline_registers.registers[3][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14200_ (.CLK(clknet_leaf_256_clk),
    .D(_00825_),
    .Q(\core_pipeline.pipeline_registers.registers[3][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14201_ (.CLK(clknet_leaf_199_clk),
    .D(_00826_),
    .Q(\core_pipeline.pipeline_registers.registers[3][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14202_ (.CLK(clknet_leaf_239_clk),
    .D(_00827_),
    .Q(\core_pipeline.pipeline_registers.registers[3][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14203_ (.CLK(clknet_leaf_1_clk),
    .D(_00828_),
    .Q(\core_pipeline.pipeline_registers.registers[3][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14204_ (.CLK(clknet_leaf_241_clk),
    .D(_00829_),
    .Q(\core_pipeline.pipeline_registers.registers[3][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14205_ (.CLK(clknet_leaf_3_clk),
    .D(_00830_),
    .Q(\core_pipeline.pipeline_registers.registers[3][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14206_ (.CLK(clknet_leaf_48_clk),
    .D(_00831_),
    .Q(\core_pipeline.pipeline_registers.registers[3][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14207_ (.CLK(clknet_leaf_4_clk),
    .D(_00832_),
    .Q(\core_pipeline.pipeline_registers.registers[3][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14208_ (.CLK(clknet_leaf_231_clk),
    .D(_00833_),
    .Q(\core_pipeline.pipeline_registers.registers[3][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14209_ (.CLK(clknet_leaf_16_clk),
    .D(_00834_),
    .Q(\core_pipeline.pipeline_registers.registers[3][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14210_ (.CLK(clknet_leaf_49_clk),
    .D(_00835_),
    .Q(\core_pipeline.pipeline_registers.registers[3][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14211_ (.CLK(clknet_leaf_19_clk),
    .D(_00836_),
    .Q(\core_pipeline.pipeline_registers.registers[3][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14212_ (.CLK(clknet_leaf_251_clk),
    .D(_00837_),
    .Q(\core_pipeline.pipeline_registers.registers[3][16] ));
 sky130_fd_sc_hd__dfxtp_1 _14213_ (.CLK(clknet_leaf_196_clk),
    .D(_00838_),
    .Q(\core_pipeline.pipeline_registers.registers[3][17] ));
 sky130_fd_sc_hd__dfxtp_1 _14214_ (.CLK(clknet_leaf_175_clk),
    .D(_00839_),
    .Q(\core_pipeline.pipeline_registers.registers[3][18] ));
 sky130_fd_sc_hd__dfxtp_1 _14215_ (.CLK(clknet_leaf_192_clk),
    .D(_00840_),
    .Q(\core_pipeline.pipeline_registers.registers[3][19] ));
 sky130_fd_sc_hd__dfxtp_1 _14216_ (.CLK(clknet_leaf_187_clk),
    .D(_00841_),
    .Q(\core_pipeline.pipeline_registers.registers[3][20] ));
 sky130_fd_sc_hd__dfxtp_1 _14217_ (.CLK(clknet_leaf_172_clk),
    .D(_00842_),
    .Q(\core_pipeline.pipeline_registers.registers[3][21] ));
 sky130_fd_sc_hd__dfxtp_1 _14218_ (.CLK(clknet_leaf_207_clk),
    .D(_00843_),
    .Q(\core_pipeline.pipeline_registers.registers[3][22] ));
 sky130_fd_sc_hd__dfxtp_1 _14219_ (.CLK(clknet_leaf_218_clk),
    .D(_00844_),
    .Q(\core_pipeline.pipeline_registers.registers[3][23] ));
 sky130_fd_sc_hd__dfxtp_1 _14220_ (.CLK(clknet_leaf_227_clk),
    .D(_00845_),
    .Q(\core_pipeline.pipeline_registers.registers[3][24] ));
 sky130_fd_sc_hd__dfxtp_1 _14221_ (.CLK(clknet_leaf_13_clk),
    .D(_00846_),
    .Q(\core_pipeline.pipeline_registers.registers[3][25] ));
 sky130_fd_sc_hd__dfxtp_1 _14222_ (.CLK(clknet_leaf_48_clk),
    .D(_00847_),
    .Q(\core_pipeline.pipeline_registers.registers[3][26] ));
 sky130_fd_sc_hd__dfxtp_1 _14223_ (.CLK(clknet_leaf_171_clk),
    .D(_00848_),
    .Q(\core_pipeline.pipeline_registers.registers[3][27] ));
 sky130_fd_sc_hd__dfxtp_1 _14224_ (.CLK(clknet_leaf_184_clk),
    .D(_00849_),
    .Q(\core_pipeline.pipeline_registers.registers[3][28] ));
 sky130_fd_sc_hd__dfxtp_1 _14225_ (.CLK(clknet_leaf_162_clk),
    .D(_00850_),
    .Q(\core_pipeline.pipeline_registers.registers[3][29] ));
 sky130_fd_sc_hd__dfxtp_1 _14226_ (.CLK(clknet_leaf_208_clk),
    .D(_00851_),
    .Q(\core_pipeline.pipeline_registers.registers[3][30] ));
 sky130_fd_sc_hd__dfxtp_1 _14227_ (.CLK(clknet_leaf_172_clk),
    .D(_00852_),
    .Q(\core_pipeline.pipeline_registers.registers[3][31] ));
 sky130_fd_sc_hd__dfxtp_1 _14228_ (.CLK(clknet_leaf_253_clk),
    .D(_00853_),
    .Q(\core_pipeline.pipeline_registers.registers[4][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14229_ (.CLK(clknet_leaf_166_clk),
    .D(_00854_),
    .Q(\core_pipeline.pipeline_registers.registers[4][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14230_ (.CLK(clknet_leaf_193_clk),
    .D(_00855_),
    .Q(\core_pipeline.pipeline_registers.registers[4][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14231_ (.CLK(clknet_leaf_237_clk),
    .D(_00856_),
    .Q(\core_pipeline.pipeline_registers.registers[4][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14232_ (.CLK(clknet_leaf_254_clk),
    .D(_00857_),
    .Q(\core_pipeline.pipeline_registers.registers[4][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14233_ (.CLK(clknet_leaf_199_clk),
    .D(_00858_),
    .Q(\core_pipeline.pipeline_registers.registers[4][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14234_ (.CLK(clknet_leaf_205_clk),
    .D(_00859_),
    .Q(\core_pipeline.pipeline_registers.registers[4][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14235_ (.CLK(clknet_leaf_5_clk),
    .D(_00860_),
    .Q(\core_pipeline.pipeline_registers.registers[4][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14236_ (.CLK(clknet_leaf_239_clk),
    .D(_00861_),
    .Q(\core_pipeline.pipeline_registers.registers[4][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14237_ (.CLK(clknet_leaf_3_clk),
    .D(_00862_),
    .Q(\core_pipeline.pipeline_registers.registers[4][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14238_ (.CLK(clknet_leaf_16_clk),
    .D(_00863_),
    .Q(\core_pipeline.pipeline_registers.registers[4][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14239_ (.CLK(clknet_leaf_4_clk),
    .D(_00864_),
    .Q(\core_pipeline.pipeline_registers.registers[4][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14240_ (.CLK(clknet_leaf_247_clk),
    .D(_00865_),
    .Q(\core_pipeline.pipeline_registers.registers[4][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14241_ (.CLK(clknet_leaf_17_clk),
    .D(_00866_),
    .Q(\core_pipeline.pipeline_registers.registers[4][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14242_ (.CLK(clknet_leaf_49_clk),
    .D(_00867_),
    .Q(\core_pipeline.pipeline_registers.registers[4][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14243_ (.CLK(clknet_leaf_46_clk),
    .D(_00868_),
    .Q(\core_pipeline.pipeline_registers.registers[4][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14244_ (.CLK(clknet_leaf_252_clk),
    .D(_00869_),
    .Q(\core_pipeline.pipeline_registers.registers[4][16] ));
 sky130_fd_sc_hd__dfxtp_1 _14245_ (.CLK(clknet_leaf_180_clk),
    .D(_00870_),
    .Q(\core_pipeline.pipeline_registers.registers[4][17] ));
 sky130_fd_sc_hd__dfxtp_1 _14246_ (.CLK(clknet_leaf_175_clk),
    .D(_00871_),
    .Q(\core_pipeline.pipeline_registers.registers[4][18] ));
 sky130_fd_sc_hd__dfxtp_1 _14247_ (.CLK(clknet_leaf_191_clk),
    .D(_00872_),
    .Q(\core_pipeline.pipeline_registers.registers[4][19] ));
 sky130_fd_sc_hd__dfxtp_1 _14248_ (.CLK(clknet_leaf_188_clk),
    .D(_00873_),
    .Q(\core_pipeline.pipeline_registers.registers[4][20] ));
 sky130_fd_sc_hd__dfxtp_1 _14249_ (.CLK(clknet_leaf_171_clk),
    .D(_00874_),
    .Q(\core_pipeline.pipeline_registers.registers[4][21] ));
 sky130_fd_sc_hd__dfxtp_1 _14250_ (.CLK(clknet_leaf_203_clk),
    .D(_00875_),
    .Q(\core_pipeline.pipeline_registers.registers[4][22] ));
 sky130_fd_sc_hd__dfxtp_1 _14251_ (.CLK(clknet_leaf_216_clk),
    .D(_00876_),
    .Q(\core_pipeline.pipeline_registers.registers[4][23] ));
 sky130_fd_sc_hd__dfxtp_1 _14252_ (.CLK(clknet_leaf_226_clk),
    .D(_00877_),
    .Q(\core_pipeline.pipeline_registers.registers[4][24] ));
 sky130_fd_sc_hd__dfxtp_1 _14253_ (.CLK(clknet_leaf_13_clk),
    .D(_00878_),
    .Q(\core_pipeline.pipeline_registers.registers[4][25] ));
 sky130_fd_sc_hd__dfxtp_1 _14254_ (.CLK(clknet_leaf_19_clk),
    .D(_00879_),
    .Q(\core_pipeline.pipeline_registers.registers[4][26] ));
 sky130_fd_sc_hd__dfxtp_1 _14255_ (.CLK(clknet_leaf_138_clk),
    .D(_00880_),
    .Q(\core_pipeline.pipeline_registers.registers[4][27] ));
 sky130_fd_sc_hd__dfxtp_1 _14256_ (.CLK(clknet_leaf_185_clk),
    .D(_00881_),
    .Q(\core_pipeline.pipeline_registers.registers[4][28] ));
 sky130_fd_sc_hd__dfxtp_1 _14257_ (.CLK(clknet_leaf_214_clk),
    .D(_00882_),
    .Q(\core_pipeline.pipeline_registers.registers[4][29] ));
 sky130_fd_sc_hd__dfxtp_1 _14258_ (.CLK(clknet_leaf_209_clk),
    .D(_00883_),
    .Q(\core_pipeline.pipeline_registers.registers[4][30] ));
 sky130_fd_sc_hd__dfxtp_1 _14259_ (.CLK(clknet_leaf_174_clk),
    .D(_00884_),
    .Q(\core_pipeline.pipeline_registers.registers[4][31] ));
 sky130_fd_sc_hd__dfxtp_1 _14260_ (.CLK(clknet_leaf_252_clk),
    .D(_00885_),
    .Q(\core_pipeline.pipeline_registers.registers[5][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14261_ (.CLK(clknet_leaf_159_clk),
    .D(_00886_),
    .Q(\core_pipeline.pipeline_registers.registers[5][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14262_ (.CLK(clknet_leaf_193_clk),
    .D(_00887_),
    .Q(\core_pipeline.pipeline_registers.registers[5][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14263_ (.CLK(clknet_leaf_234_clk),
    .D(_00888_),
    .Q(\core_pipeline.pipeline_registers.registers[5][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14264_ (.CLK(clknet_leaf_254_clk),
    .D(_00889_),
    .Q(\core_pipeline.pipeline_registers.registers[5][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14265_ (.CLK(clknet_leaf_201_clk),
    .D(_00890_),
    .Q(\core_pipeline.pipeline_registers.registers[5][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14266_ (.CLK(clknet_leaf_239_clk),
    .D(_00891_),
    .Q(\core_pipeline.pipeline_registers.registers[5][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14267_ (.CLK(clknet_leaf_5_clk),
    .D(_00892_),
    .Q(\core_pipeline.pipeline_registers.registers[5][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14268_ (.CLK(clknet_leaf_240_clk),
    .D(_00893_),
    .Q(\core_pipeline.pipeline_registers.registers[5][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14269_ (.CLK(clknet_leaf_3_clk),
    .D(_00894_),
    .Q(\core_pipeline.pipeline_registers.registers[5][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14270_ (.CLK(clknet_leaf_15_clk),
    .D(_00895_),
    .Q(\core_pipeline.pipeline_registers.registers[5][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14271_ (.CLK(clknet_leaf_3_clk),
    .D(_00896_),
    .Q(\core_pipeline.pipeline_registers.registers[5][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14272_ (.CLK(clknet_leaf_231_clk),
    .D(_00897_),
    .Q(\core_pipeline.pipeline_registers.registers[5][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14273_ (.CLK(clknet_leaf_16_clk),
    .D(_00898_),
    .Q(\core_pipeline.pipeline_registers.registers[5][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14274_ (.CLK(clknet_leaf_49_clk),
    .D(_00899_),
    .Q(\core_pipeline.pipeline_registers.registers[5][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14275_ (.CLK(clknet_leaf_46_clk),
    .D(_00900_),
    .Q(\core_pipeline.pipeline_registers.registers[5][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14276_ (.CLK(clknet_leaf_252_clk),
    .D(_00901_),
    .Q(\core_pipeline.pipeline_registers.registers[5][16] ));
 sky130_fd_sc_hd__dfxtp_1 _14277_ (.CLK(clknet_leaf_163_clk),
    .D(_00902_),
    .Q(\core_pipeline.pipeline_registers.registers[5][17] ));
 sky130_fd_sc_hd__dfxtp_1 _14278_ (.CLK(clknet_leaf_175_clk),
    .D(_00903_),
    .Q(\core_pipeline.pipeline_registers.registers[5][18] ));
 sky130_fd_sc_hd__dfxtp_1 _14279_ (.CLK(clknet_leaf_191_clk),
    .D(_00904_),
    .Q(\core_pipeline.pipeline_registers.registers[5][19] ));
 sky130_fd_sc_hd__dfxtp_1 _14280_ (.CLK(clknet_leaf_187_clk),
    .D(_00905_),
    .Q(\core_pipeline.pipeline_registers.registers[5][20] ));
 sky130_fd_sc_hd__dfxtp_1 _14281_ (.CLK(clknet_leaf_171_clk),
    .D(_00906_),
    .Q(\core_pipeline.pipeline_registers.registers[5][21] ));
 sky130_fd_sc_hd__dfxtp_1 _14282_ (.CLK(clknet_leaf_203_clk),
    .D(_00907_),
    .Q(\core_pipeline.pipeline_registers.registers[5][22] ));
 sky130_fd_sc_hd__dfxtp_1 _14283_ (.CLK(clknet_leaf_216_clk),
    .D(_00908_),
    .Q(\core_pipeline.pipeline_registers.registers[5][23] ));
 sky130_fd_sc_hd__dfxtp_1 _14284_ (.CLK(clknet_leaf_227_clk),
    .D(_00909_),
    .Q(\core_pipeline.pipeline_registers.registers[5][24] ));
 sky130_fd_sc_hd__dfxtp_1 _14285_ (.CLK(clknet_leaf_13_clk),
    .D(_00910_),
    .Q(\core_pipeline.pipeline_registers.registers[5][25] ));
 sky130_fd_sc_hd__dfxtp_1 _14286_ (.CLK(clknet_leaf_19_clk),
    .D(_00911_),
    .Q(\core_pipeline.pipeline_registers.registers[5][26] ));
 sky130_fd_sc_hd__dfxtp_1 _14287_ (.CLK(clknet_leaf_138_clk),
    .D(_00912_),
    .Q(\core_pipeline.pipeline_registers.registers[5][27] ));
 sky130_fd_sc_hd__dfxtp_1 _14288_ (.CLK(clknet_leaf_185_clk),
    .D(_00913_),
    .Q(\core_pipeline.pipeline_registers.registers[5][28] ));
 sky130_fd_sc_hd__dfxtp_1 _14289_ (.CLK(clknet_leaf_215_clk),
    .D(_00914_),
    .Q(\core_pipeline.pipeline_registers.registers[5][29] ));
 sky130_fd_sc_hd__dfxtp_1 _14290_ (.CLK(clknet_leaf_226_clk),
    .D(_00915_),
    .Q(\core_pipeline.pipeline_registers.registers[5][30] ));
 sky130_fd_sc_hd__dfxtp_1 _14291_ (.CLK(clknet_leaf_174_clk),
    .D(_00916_),
    .Q(\core_pipeline.pipeline_registers.registers[5][31] ));
 sky130_fd_sc_hd__dfxtp_1 _14292_ (.CLK(clknet_leaf_253_clk),
    .D(_00917_),
    .Q(\core_pipeline.pipeline_registers.registers[6][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14293_ (.CLK(clknet_leaf_159_clk),
    .D(_00918_),
    .Q(\core_pipeline.pipeline_registers.registers[6][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14294_ (.CLK(clknet_leaf_199_clk),
    .D(_00919_),
    .Q(\core_pipeline.pipeline_registers.registers[6][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14295_ (.CLK(clknet_leaf_234_clk),
    .D(_00920_),
    .Q(\core_pipeline.pipeline_registers.registers[6][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14296_ (.CLK(clknet_leaf_1_clk),
    .D(_00921_),
    .Q(\core_pipeline.pipeline_registers.registers[6][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14297_ (.CLK(clknet_leaf_201_clk),
    .D(_00922_),
    .Q(\core_pipeline.pipeline_registers.registers[6][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14298_ (.CLK(clknet_leaf_239_clk),
    .D(_00923_),
    .Q(\core_pipeline.pipeline_registers.registers[6][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14299_ (.CLK(clknet_leaf_5_clk),
    .D(_00924_),
    .Q(\core_pipeline.pipeline_registers.registers[6][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14300_ (.CLK(clknet_leaf_241_clk),
    .D(_00925_),
    .Q(\core_pipeline.pipeline_registers.registers[6][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14301_ (.CLK(clknet_leaf_3_clk),
    .D(_00926_),
    .Q(\core_pipeline.pipeline_registers.registers[6][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14302_ (.CLK(clknet_leaf_49_clk),
    .D(_00927_),
    .Q(\core_pipeline.pipeline_registers.registers[6][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14303_ (.CLK(clknet_leaf_3_clk),
    .D(_00928_),
    .Q(\core_pipeline.pipeline_registers.registers[6][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14304_ (.CLK(clknet_leaf_248_clk),
    .D(_00929_),
    .Q(\core_pipeline.pipeline_registers.registers[6][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14305_ (.CLK(clknet_leaf_15_clk),
    .D(_00930_),
    .Q(\core_pipeline.pipeline_registers.registers[6][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14306_ (.CLK(clknet_leaf_49_clk),
    .D(_00931_),
    .Q(\core_pipeline.pipeline_registers.registers[6][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14307_ (.CLK(clknet_leaf_46_clk),
    .D(_00932_),
    .Q(\core_pipeline.pipeline_registers.registers[6][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14308_ (.CLK(clknet_leaf_252_clk),
    .D(_00933_),
    .Q(\core_pipeline.pipeline_registers.registers[6][16] ));
 sky130_fd_sc_hd__dfxtp_1 _14309_ (.CLK(clknet_leaf_163_clk),
    .D(_00934_),
    .Q(\core_pipeline.pipeline_registers.registers[6][17] ));
 sky130_fd_sc_hd__dfxtp_1 _14310_ (.CLK(clknet_leaf_175_clk),
    .D(_00935_),
    .Q(\core_pipeline.pipeline_registers.registers[6][18] ));
 sky130_fd_sc_hd__dfxtp_1 _14311_ (.CLK(clknet_leaf_192_clk),
    .D(_00936_),
    .Q(\core_pipeline.pipeline_registers.registers[6][19] ));
 sky130_fd_sc_hd__dfxtp_1 _14312_ (.CLK(clknet_leaf_187_clk),
    .D(_00937_),
    .Q(\core_pipeline.pipeline_registers.registers[6][20] ));
 sky130_fd_sc_hd__dfxtp_1 _14313_ (.CLK(clknet_leaf_170_clk),
    .D(_00938_),
    .Q(\core_pipeline.pipeline_registers.registers[6][21] ));
 sky130_fd_sc_hd__dfxtp_1 _14314_ (.CLK(clknet_leaf_204_clk),
    .D(_00939_),
    .Q(\core_pipeline.pipeline_registers.registers[6][22] ));
 sky130_fd_sc_hd__dfxtp_1 _14315_ (.CLK(clknet_leaf_218_clk),
    .D(_00940_),
    .Q(\core_pipeline.pipeline_registers.registers[6][23] ));
 sky130_fd_sc_hd__dfxtp_1 _14316_ (.CLK(clknet_leaf_228_clk),
    .D(_00941_),
    .Q(\core_pipeline.pipeline_registers.registers[6][24] ));
 sky130_fd_sc_hd__dfxtp_1 _14317_ (.CLK(clknet_leaf_12_clk),
    .D(_00942_),
    .Q(\core_pipeline.pipeline_registers.registers[6][25] ));
 sky130_fd_sc_hd__dfxtp_1 _14318_ (.CLK(clknet_leaf_16_clk),
    .D(_00943_),
    .Q(\core_pipeline.pipeline_registers.registers[6][26] ));
 sky130_fd_sc_hd__dfxtp_1 _14319_ (.CLK(clknet_leaf_138_clk),
    .D(_00944_),
    .Q(\core_pipeline.pipeline_registers.registers[6][27] ));
 sky130_fd_sc_hd__dfxtp_1 _14320_ (.CLK(clknet_leaf_186_clk),
    .D(_00945_),
    .Q(\core_pipeline.pipeline_registers.registers[6][28] ));
 sky130_fd_sc_hd__dfxtp_1 _14321_ (.CLK(clknet_leaf_215_clk),
    .D(_00946_),
    .Q(\core_pipeline.pipeline_registers.registers[6][29] ));
 sky130_fd_sc_hd__dfxtp_1 _14322_ (.CLK(clknet_leaf_236_clk),
    .D(_00947_),
    .Q(\core_pipeline.pipeline_registers.registers[6][30] ));
 sky130_fd_sc_hd__dfxtp_1 _14323_ (.CLK(clknet_leaf_174_clk),
    .D(_00948_),
    .Q(\core_pipeline.pipeline_registers.registers[6][31] ));
 sky130_fd_sc_hd__dfxtp_1 _14324_ (.CLK(clknet_leaf_253_clk),
    .D(_00949_),
    .Q(\core_pipeline.pipeline_registers.registers[7][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14325_ (.CLK(clknet_leaf_159_clk),
    .D(_00950_),
    .Q(\core_pipeline.pipeline_registers.registers[7][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14326_ (.CLK(clknet_leaf_199_clk),
    .D(_00951_),
    .Q(\core_pipeline.pipeline_registers.registers[7][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14327_ (.CLK(clknet_leaf_234_clk),
    .D(_00952_),
    .Q(\core_pipeline.pipeline_registers.registers[7][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14328_ (.CLK(clknet_leaf_1_clk),
    .D(_00953_),
    .Q(\core_pipeline.pipeline_registers.registers[7][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14329_ (.CLK(clknet_leaf_201_clk),
    .D(_00954_),
    .Q(\core_pipeline.pipeline_registers.registers[7][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14330_ (.CLK(clknet_leaf_239_clk),
    .D(_00955_),
    .Q(\core_pipeline.pipeline_registers.registers[7][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14331_ (.CLK(clknet_leaf_4_clk),
    .D(_00956_),
    .Q(\core_pipeline.pipeline_registers.registers[7][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14332_ (.CLK(clknet_leaf_241_clk),
    .D(_00957_),
    .Q(\core_pipeline.pipeline_registers.registers[7][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14333_ (.CLK(clknet_leaf_3_clk),
    .D(_00958_),
    .Q(\core_pipeline.pipeline_registers.registers[7][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14334_ (.CLK(clknet_leaf_16_clk),
    .D(_00959_),
    .Q(\core_pipeline.pipeline_registers.registers[7][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14335_ (.CLK(clknet_leaf_3_clk),
    .D(_00960_),
    .Q(\core_pipeline.pipeline_registers.registers[7][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14336_ (.CLK(clknet_leaf_247_clk),
    .D(_00961_),
    .Q(\core_pipeline.pipeline_registers.registers[7][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14337_ (.CLK(clknet_leaf_14_clk),
    .D(_00962_),
    .Q(\core_pipeline.pipeline_registers.registers[7][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14338_ (.CLK(clknet_leaf_49_clk),
    .D(_00963_),
    .Q(\core_pipeline.pipeline_registers.registers[7][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14339_ (.CLK(clknet_leaf_46_clk),
    .D(_00964_),
    .Q(\core_pipeline.pipeline_registers.registers[7][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14340_ (.CLK(clknet_leaf_252_clk),
    .D(_00965_),
    .Q(\core_pipeline.pipeline_registers.registers[7][16] ));
 sky130_fd_sc_hd__dfxtp_1 _14341_ (.CLK(clknet_leaf_163_clk),
    .D(_00966_),
    .Q(\core_pipeline.pipeline_registers.registers[7][17] ));
 sky130_fd_sc_hd__dfxtp_1 _14342_ (.CLK(clknet_leaf_175_clk),
    .D(_00967_),
    .Q(\core_pipeline.pipeline_registers.registers[7][18] ));
 sky130_fd_sc_hd__dfxtp_1 _14343_ (.CLK(clknet_leaf_191_clk),
    .D(_00968_),
    .Q(\core_pipeline.pipeline_registers.registers[7][19] ));
 sky130_fd_sc_hd__dfxtp_1 _14344_ (.CLK(clknet_leaf_189_clk),
    .D(_00969_),
    .Q(\core_pipeline.pipeline_registers.registers[7][20] ));
 sky130_fd_sc_hd__dfxtp_1 _14345_ (.CLK(clknet_leaf_170_clk),
    .D(_00970_),
    .Q(\core_pipeline.pipeline_registers.registers[7][21] ));
 sky130_fd_sc_hd__dfxtp_1 _14346_ (.CLK(clknet_leaf_203_clk),
    .D(_00971_),
    .Q(\core_pipeline.pipeline_registers.registers[7][22] ));
 sky130_fd_sc_hd__dfxtp_1 _14347_ (.CLK(clknet_leaf_216_clk),
    .D(_00972_),
    .Q(\core_pipeline.pipeline_registers.registers[7][23] ));
 sky130_fd_sc_hd__dfxtp_1 _14348_ (.CLK(clknet_leaf_227_clk),
    .D(_00973_),
    .Q(\core_pipeline.pipeline_registers.registers[7][24] ));
 sky130_fd_sc_hd__dfxtp_1 _14349_ (.CLK(clknet_leaf_12_clk),
    .D(_00974_),
    .Q(\core_pipeline.pipeline_registers.registers[7][25] ));
 sky130_fd_sc_hd__dfxtp_1 _14350_ (.CLK(clknet_leaf_17_clk),
    .D(_00975_),
    .Q(\core_pipeline.pipeline_registers.registers[7][26] ));
 sky130_fd_sc_hd__dfxtp_1 _14351_ (.CLK(clknet_leaf_138_clk),
    .D(_00976_),
    .Q(\core_pipeline.pipeline_registers.registers[7][27] ));
 sky130_fd_sc_hd__dfxtp_1 _14352_ (.CLK(clknet_leaf_184_clk),
    .D(_00977_),
    .Q(\core_pipeline.pipeline_registers.registers[7][28] ));
 sky130_fd_sc_hd__dfxtp_1 _14353_ (.CLK(clknet_leaf_215_clk),
    .D(_00978_),
    .Q(\core_pipeline.pipeline_registers.registers[7][29] ));
 sky130_fd_sc_hd__dfxtp_1 _14354_ (.CLK(clknet_leaf_236_clk),
    .D(_00979_),
    .Q(\core_pipeline.pipeline_registers.registers[7][30] ));
 sky130_fd_sc_hd__dfxtp_1 _14355_ (.CLK(clknet_leaf_174_clk),
    .D(_00980_),
    .Q(\core_pipeline.pipeline_registers.registers[7][31] ));
 sky130_fd_sc_hd__dfxtp_1 _14356_ (.CLK(clknet_leaf_253_clk),
    .D(_00981_),
    .Q(\core_pipeline.pipeline_registers.registers[8][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14357_ (.CLK(clknet_leaf_164_clk),
    .D(_00982_),
    .Q(\core_pipeline.pipeline_registers.registers[8][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14358_ (.CLK(clknet_leaf_192_clk),
    .D(_00983_),
    .Q(\core_pipeline.pipeline_registers.registers[8][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14359_ (.CLK(clknet_leaf_233_clk),
    .D(_00984_),
    .Q(\core_pipeline.pipeline_registers.registers[8][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14360_ (.CLK(clknet_leaf_256_clk),
    .D(_00985_),
    .Q(\core_pipeline.pipeline_registers.registers[8][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14361_ (.CLK(clknet_leaf_200_clk),
    .D(_00986_),
    .Q(\core_pipeline.pipeline_registers.registers[8][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14362_ (.CLK(clknet_leaf_205_clk),
    .D(_00987_),
    .Q(\core_pipeline.pipeline_registers.registers[8][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14363_ (.CLK(clknet_leaf_2_clk),
    .D(_00988_),
    .Q(\core_pipeline.pipeline_registers.registers[8][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14364_ (.CLK(clknet_leaf_240_clk),
    .D(_00989_),
    .Q(\core_pipeline.pipeline_registers.registers[8][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14365_ (.CLK(clknet_leaf_11_clk),
    .D(_00990_),
    .Q(\core_pipeline.pipeline_registers.registers[8][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14366_ (.CLK(clknet_leaf_14_clk),
    .D(_00991_),
    .Q(\core_pipeline.pipeline_registers.registers[8][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14367_ (.CLK(clknet_leaf_2_clk),
    .D(_00992_),
    .Q(\core_pipeline.pipeline_registers.registers[8][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14368_ (.CLK(clknet_leaf_248_clk),
    .D(_00993_),
    .Q(\core_pipeline.pipeline_registers.registers[8][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14369_ (.CLK(clknet_leaf_10_clk),
    .D(_00994_),
    .Q(\core_pipeline.pipeline_registers.registers[8][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14370_ (.CLK(clknet_leaf_15_clk),
    .D(_00995_),
    .Q(\core_pipeline.pipeline_registers.registers[8][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14371_ (.CLK(clknet_leaf_20_clk),
    .D(_00996_),
    .Q(\core_pipeline.pipeline_registers.registers[8][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14372_ (.CLK(clknet_leaf_244_clk),
    .D(_00997_),
    .Q(\core_pipeline.pipeline_registers.registers[8][16] ));
 sky130_fd_sc_hd__dfxtp_1 _14373_ (.CLK(clknet_leaf_196_clk),
    .D(_00998_),
    .Q(\core_pipeline.pipeline_registers.registers[8][17] ));
 sky130_fd_sc_hd__dfxtp_1 _14374_ (.CLK(clknet_leaf_186_clk),
    .D(_00999_),
    .Q(\core_pipeline.pipeline_registers.registers[8][18] ));
 sky130_fd_sc_hd__dfxtp_1 _14375_ (.CLK(clknet_leaf_191_clk),
    .D(_01000_),
    .Q(\core_pipeline.pipeline_registers.registers[8][19] ));
 sky130_fd_sc_hd__dfxtp_1 _14376_ (.CLK(clknet_leaf_188_clk),
    .D(_01001_),
    .Q(\core_pipeline.pipeline_registers.registers[8][20] ));
 sky130_fd_sc_hd__dfxtp_1 _14377_ (.CLK(clknet_leaf_172_clk),
    .D(_01002_),
    .Q(\core_pipeline.pipeline_registers.registers[8][21] ));
 sky130_fd_sc_hd__dfxtp_1 _14378_ (.CLK(clknet_leaf_203_clk),
    .D(_01003_),
    .Q(\core_pipeline.pipeline_registers.registers[8][22] ));
 sky130_fd_sc_hd__dfxtp_1 _14379_ (.CLK(clknet_leaf_218_clk),
    .D(_01004_),
    .Q(\core_pipeline.pipeline_registers.registers[8][23] ));
 sky130_fd_sc_hd__dfxtp_1 _14380_ (.CLK(clknet_leaf_236_clk),
    .D(_01005_),
    .Q(\core_pipeline.pipeline_registers.registers[8][24] ));
 sky130_fd_sc_hd__dfxtp_1 _14381_ (.CLK(clknet_leaf_12_clk),
    .D(_01006_),
    .Q(\core_pipeline.pipeline_registers.registers[8][25] ));
 sky130_fd_sc_hd__dfxtp_1 _14382_ (.CLK(clknet_leaf_17_clk),
    .D(_01007_),
    .Q(\core_pipeline.pipeline_registers.registers[8][26] ));
 sky130_fd_sc_hd__dfxtp_1 _14383_ (.CLK(clknet_leaf_138_clk),
    .D(_01008_),
    .Q(\core_pipeline.pipeline_registers.registers[8][27] ));
 sky130_fd_sc_hd__dfxtp_1 _14384_ (.CLK(clknet_leaf_184_clk),
    .D(_01009_),
    .Q(\core_pipeline.pipeline_registers.registers[8][28] ));
 sky130_fd_sc_hd__dfxtp_1 _14385_ (.CLK(clknet_leaf_213_clk),
    .D(_01010_),
    .Q(\core_pipeline.pipeline_registers.registers[8][29] ));
 sky130_fd_sc_hd__dfxtp_1 _14386_ (.CLK(clknet_leaf_208_clk),
    .D(_01011_),
    .Q(\core_pipeline.pipeline_registers.registers[8][30] ));
 sky130_fd_sc_hd__dfxtp_1 _14387_ (.CLK(clknet_leaf_174_clk),
    .D(_01012_),
    .Q(\core_pipeline.pipeline_registers.registers[8][31] ));
 sky130_fd_sc_hd__dfxtp_1 _14388_ (.CLK(clknet_leaf_151_clk),
    .D(_01013_),
    .Q(\core_pipeline.pipeline_fetch.pc[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14389_ (.CLK(clknet_leaf_152_clk),
    .D(_01014_),
    .Q(\core_pipeline.pipeline_fetch.pc[1] ));
 sky130_fd_sc_hd__dfxtp_1 _14390_ (.CLK(clknet_leaf_245_clk),
    .D(_01015_),
    .Q(\core_pipeline.pipeline_registers.registers[29][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14391_ (.CLK(clknet_leaf_164_clk),
    .D(_01016_),
    .Q(\core_pipeline.pipeline_registers.registers[29][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14392_ (.CLK(clknet_leaf_199_clk),
    .D(_01017_),
    .Q(\core_pipeline.pipeline_registers.registers[29][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14393_ (.CLK(clknet_leaf_237_clk),
    .D(_01018_),
    .Q(\core_pipeline.pipeline_registers.registers[29][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14394_ (.CLK(clknet_leaf_251_clk),
    .D(_01019_),
    .Q(\core_pipeline.pipeline_registers.registers[29][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14395_ (.CLK(clknet_leaf_202_clk),
    .D(_01020_),
    .Q(\core_pipeline.pipeline_registers.registers[29][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14396_ (.CLK(clknet_leaf_205_clk),
    .D(_01021_),
    .Q(\core_pipeline.pipeline_registers.registers[29][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14397_ (.CLK(clknet_leaf_235_clk),
    .D(_01022_),
    .Q(\core_pipeline.pipeline_registers.registers[29][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14398_ (.CLK(clknet_leaf_242_clk),
    .D(_01023_),
    .Q(\core_pipeline.pipeline_registers.registers[29][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14399_ (.CLK(clknet_leaf_231_clk),
    .D(_01024_),
    .Q(\core_pipeline.pipeline_registers.registers[29][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14400_ (.CLK(clknet_leaf_8_clk),
    .D(_01025_),
    .Q(\core_pipeline.pipeline_registers.registers[29][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14401_ (.CLK(clknet_leaf_247_clk),
    .D(_01026_),
    .Q(\core_pipeline.pipeline_registers.registers[29][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14402_ (.CLK(clknet_leaf_229_clk),
    .D(_01027_),
    .Q(\core_pipeline.pipeline_registers.registers[29][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14403_ (.CLK(clknet_leaf_22_clk),
    .D(_01028_),
    .Q(\core_pipeline.pipeline_registers.registers[29][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14404_ (.CLK(clknet_leaf_7_clk),
    .D(_01029_),
    .Q(\core_pipeline.pipeline_registers.registers[29][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14405_ (.CLK(clknet_leaf_24_clk),
    .D(_01030_),
    .Q(\core_pipeline.pipeline_registers.registers[29][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14406_ (.CLK(clknet_leaf_245_clk),
    .D(_01031_),
    .Q(\core_pipeline.pipeline_registers.registers[29][16] ));
 sky130_fd_sc_hd__dfxtp_1 _14407_ (.CLK(clknet_leaf_195_clk),
    .D(_01032_),
    .Q(\core_pipeline.pipeline_registers.registers[29][17] ));
 sky130_fd_sc_hd__dfxtp_1 _14408_ (.CLK(clknet_leaf_181_clk),
    .D(_01033_),
    .Q(\core_pipeline.pipeline_registers.registers[29][18] ));
 sky130_fd_sc_hd__dfxtp_1 _14409_ (.CLK(clknet_leaf_194_clk),
    .D(_01034_),
    .Q(\core_pipeline.pipeline_registers.registers[29][19] ));
 sky130_fd_sc_hd__dfxtp_1 _14410_ (.CLK(clknet_leaf_190_clk),
    .D(_01035_),
    .Q(\core_pipeline.pipeline_registers.registers[29][20] ));
 sky130_fd_sc_hd__dfxtp_1 _14411_ (.CLK(clknet_leaf_177_clk),
    .D(_01036_),
    .Q(\core_pipeline.pipeline_registers.registers[29][21] ));
 sky130_fd_sc_hd__dfxtp_1 _14412_ (.CLK(clknet_leaf_211_clk),
    .D(_01037_),
    .Q(\core_pipeline.pipeline_registers.registers[29][22] ));
 sky130_fd_sc_hd__dfxtp_1 _14413_ (.CLK(clknet_leaf_216_clk),
    .D(_01038_),
    .Q(\core_pipeline.pipeline_registers.registers[29][23] ));
 sky130_fd_sc_hd__dfxtp_1 _14414_ (.CLK(clknet_leaf_225_clk),
    .D(_01039_),
    .Q(\core_pipeline.pipeline_registers.registers[29][24] ));
 sky130_fd_sc_hd__dfxtp_1 _14415_ (.CLK(clknet_leaf_7_clk),
    .D(_01040_),
    .Q(\core_pipeline.pipeline_registers.registers[29][25] ));
 sky130_fd_sc_hd__dfxtp_1 _14416_ (.CLK(clknet_leaf_21_clk),
    .D(_01041_),
    .Q(\core_pipeline.pipeline_registers.registers[29][26] ));
 sky130_fd_sc_hd__dfxtp_1 _14417_ (.CLK(clknet_leaf_169_clk),
    .D(_01042_),
    .Q(\core_pipeline.pipeline_registers.registers[29][27] ));
 sky130_fd_sc_hd__dfxtp_1 _14418_ (.CLK(clknet_leaf_182_clk),
    .D(_01043_),
    .Q(\core_pipeline.pipeline_registers.registers[29][28] ));
 sky130_fd_sc_hd__dfxtp_1 _14419_ (.CLK(clknet_leaf_212_clk),
    .D(_01044_),
    .Q(\core_pipeline.pipeline_registers.registers[29][29] ));
 sky130_fd_sc_hd__dfxtp_1 _14420_ (.CLK(clknet_leaf_208_clk),
    .D(_01045_),
    .Q(\core_pipeline.pipeline_registers.registers[29][30] ));
 sky130_fd_sc_hd__dfxtp_1 _14421_ (.CLK(clknet_leaf_178_clk),
    .D(_01046_),
    .Q(\core_pipeline.pipeline_registers.registers[29][31] ));
 sky130_fd_sc_hd__dfxtp_1 _14422_ (.CLK(clknet_leaf_254_clk),
    .D(_01047_),
    .Q(\core_pipeline.pipeline_registers.registers[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14423_ (.CLK(clknet_leaf_159_clk),
    .D(_01048_),
    .Q(\core_pipeline.pipeline_registers.registers[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14424_ (.CLK(clknet_leaf_195_clk),
    .D(_01049_),
    .Q(\core_pipeline.pipeline_registers.registers[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14425_ (.CLK(clknet_leaf_238_clk),
    .D(_01050_),
    .Q(\core_pipeline.pipeline_registers.registers[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14426_ (.CLK(clknet_leaf_1_clk),
    .D(_01051_),
    .Q(\core_pipeline.pipeline_registers.registers[1][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14427_ (.CLK(clknet_leaf_199_clk),
    .D(_01052_),
    .Q(\core_pipeline.pipeline_registers.registers[1][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14428_ (.CLK(clknet_leaf_239_clk),
    .D(_01053_),
    .Q(\core_pipeline.pipeline_registers.registers[1][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14429_ (.CLK(clknet_leaf_1_clk),
    .D(_01054_),
    .Q(\core_pipeline.pipeline_registers.registers[1][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14430_ (.CLK(clknet_leaf_238_clk),
    .D(_01055_),
    .Q(\core_pipeline.pipeline_registers.registers[1][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14431_ (.CLK(clknet_leaf_4_clk),
    .D(_01056_),
    .Q(\core_pipeline.pipeline_registers.registers[1][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14432_ (.CLK(clknet_leaf_48_clk),
    .D(_01057_),
    .Q(\core_pipeline.pipeline_registers.registers[1][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14433_ (.CLK(clknet_leaf_4_clk),
    .D(_01058_),
    .Q(\core_pipeline.pipeline_registers.registers[1][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14434_ (.CLK(clknet_leaf_247_clk),
    .D(_01059_),
    .Q(\core_pipeline.pipeline_registers.registers[1][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14435_ (.CLK(clknet_leaf_48_clk),
    .D(_01060_),
    .Q(\core_pipeline.pipeline_registers.registers[1][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14436_ (.CLK(clknet_leaf_48_clk),
    .D(_01061_),
    .Q(\core_pipeline.pipeline_registers.registers[1][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14437_ (.CLK(clknet_leaf_19_clk),
    .D(_01062_),
    .Q(\core_pipeline.pipeline_registers.registers[1][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14438_ (.CLK(clknet_leaf_251_clk),
    .D(_01063_),
    .Q(\core_pipeline.pipeline_registers.registers[1][16] ));
 sky130_fd_sc_hd__dfxtp_1 _14439_ (.CLK(clknet_leaf_180_clk),
    .D(_01064_),
    .Q(\core_pipeline.pipeline_registers.registers[1][17] ));
 sky130_fd_sc_hd__dfxtp_1 _14440_ (.CLK(clknet_leaf_175_clk),
    .D(_01065_),
    .Q(\core_pipeline.pipeline_registers.registers[1][18] ));
 sky130_fd_sc_hd__dfxtp_1 _14441_ (.CLK(clknet_leaf_193_clk),
    .D(_01066_),
    .Q(\core_pipeline.pipeline_registers.registers[1][19] ));
 sky130_fd_sc_hd__dfxtp_1 _14442_ (.CLK(clknet_leaf_187_clk),
    .D(_01067_),
    .Q(\core_pipeline.pipeline_registers.registers[1][20] ));
 sky130_fd_sc_hd__dfxtp_1 _14443_ (.CLK(clknet_leaf_171_clk),
    .D(_01068_),
    .Q(\core_pipeline.pipeline_registers.registers[1][21] ));
 sky130_fd_sc_hd__dfxtp_1 _14444_ (.CLK(clknet_leaf_202_clk),
    .D(_01069_),
    .Q(\core_pipeline.pipeline_registers.registers[1][22] ));
 sky130_fd_sc_hd__dfxtp_1 _14445_ (.CLK(clknet_leaf_219_clk),
    .D(_01070_),
    .Q(\core_pipeline.pipeline_registers.registers[1][23] ));
 sky130_fd_sc_hd__dfxtp_1 _14446_ (.CLK(clknet_leaf_227_clk),
    .D(_01071_),
    .Q(\core_pipeline.pipeline_registers.registers[1][24] ));
 sky130_fd_sc_hd__dfxtp_1 _14447_ (.CLK(clknet_leaf_13_clk),
    .D(_01072_),
    .Q(\core_pipeline.pipeline_registers.registers[1][25] ));
 sky130_fd_sc_hd__dfxtp_1 _14448_ (.CLK(clknet_leaf_48_clk),
    .D(_01073_),
    .Q(\core_pipeline.pipeline_registers.registers[1][26] ));
 sky130_fd_sc_hd__dfxtp_1 _14449_ (.CLK(clknet_leaf_138_clk),
    .D(_01074_),
    .Q(\core_pipeline.pipeline_registers.registers[1][27] ));
 sky130_fd_sc_hd__dfxtp_1 _14450_ (.CLK(clknet_leaf_184_clk),
    .D(_01075_),
    .Q(\core_pipeline.pipeline_registers.registers[1][28] ));
 sky130_fd_sc_hd__dfxtp_1 _14451_ (.CLK(clknet_leaf_161_clk),
    .D(_01076_),
    .Q(\core_pipeline.pipeline_registers.registers[1][29] ));
 sky130_fd_sc_hd__dfxtp_1 _14452_ (.CLK(clknet_leaf_209_clk),
    .D(_01077_),
    .Q(\core_pipeline.pipeline_registers.registers[1][30] ));
 sky130_fd_sc_hd__dfxtp_1 _14453_ (.CLK(clknet_leaf_172_clk),
    .D(_01078_),
    .Q(\core_pipeline.pipeline_registers.registers[1][31] ));
 sky130_fd_sc_hd__dfxtp_1 _14454_ (.CLK(clknet_leaf_253_clk),
    .D(_01079_),
    .Q(\core_pipeline.pipeline_registers.registers[0][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14455_ (.CLK(clknet_leaf_159_clk),
    .D(_01080_),
    .Q(\core_pipeline.pipeline_registers.registers[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14456_ (.CLK(clknet_leaf_195_clk),
    .D(_01081_),
    .Q(\core_pipeline.pipeline_registers.registers[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14457_ (.CLK(clknet_leaf_238_clk),
    .D(_01082_),
    .Q(\core_pipeline.pipeline_registers.registers[0][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14458_ (.CLK(clknet_leaf_254_clk),
    .D(_01083_),
    .Q(\core_pipeline.pipeline_registers.registers[0][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14459_ (.CLK(clknet_leaf_199_clk),
    .D(_01084_),
    .Q(\core_pipeline.pipeline_registers.registers[0][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14460_ (.CLK(clknet_leaf_205_clk),
    .D(_01085_),
    .Q(\core_pipeline.pipeline_registers.registers[0][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14461_ (.CLK(clknet_leaf_250_clk),
    .D(_01086_),
    .Q(\core_pipeline.pipeline_registers.registers[0][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14462_ (.CLK(clknet_leaf_239_clk),
    .D(_01087_),
    .Q(\core_pipeline.pipeline_registers.registers[0][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14463_ (.CLK(clknet_leaf_4_clk),
    .D(_01088_),
    .Q(\core_pipeline.pipeline_registers.registers[0][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14464_ (.CLK(clknet_leaf_48_clk),
    .D(_01089_),
    .Q(\core_pipeline.pipeline_registers.registers[0][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14465_ (.CLK(clknet_leaf_4_clk),
    .D(_01090_),
    .Q(\core_pipeline.pipeline_registers.registers[0][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14466_ (.CLK(clknet_leaf_233_clk),
    .D(_01091_),
    .Q(\core_pipeline.pipeline_registers.registers[0][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14467_ (.CLK(clknet_leaf_16_clk),
    .D(_01092_),
    .Q(\core_pipeline.pipeline_registers.registers[0][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14468_ (.CLK(clknet_leaf_49_clk),
    .D(_01093_),
    .Q(\core_pipeline.pipeline_registers.registers[0][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14469_ (.CLK(clknet_leaf_20_clk),
    .D(_01094_),
    .Q(\core_pipeline.pipeline_registers.registers[0][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14470_ (.CLK(clknet_leaf_244_clk),
    .D(_01095_),
    .Q(\core_pipeline.pipeline_registers.registers[0][16] ));
 sky130_fd_sc_hd__dfxtp_1 _14471_ (.CLK(clknet_leaf_181_clk),
    .D(_01096_),
    .Q(\core_pipeline.pipeline_registers.registers[0][17] ));
 sky130_fd_sc_hd__dfxtp_1 _14472_ (.CLK(clknet_leaf_175_clk),
    .D(_01097_),
    .Q(\core_pipeline.pipeline_registers.registers[0][18] ));
 sky130_fd_sc_hd__dfxtp_1 _14473_ (.CLK(clknet_leaf_193_clk),
    .D(_01098_),
    .Q(\core_pipeline.pipeline_registers.registers[0][19] ));
 sky130_fd_sc_hd__dfxtp_1 _14474_ (.CLK(clknet_leaf_188_clk),
    .D(_01099_),
    .Q(\core_pipeline.pipeline_registers.registers[0][20] ));
 sky130_fd_sc_hd__dfxtp_1 _14475_ (.CLK(clknet_leaf_172_clk),
    .D(_01100_),
    .Q(\core_pipeline.pipeline_registers.registers[0][21] ));
 sky130_fd_sc_hd__dfxtp_1 _14476_ (.CLK(clknet_leaf_202_clk),
    .D(_01101_),
    .Q(\core_pipeline.pipeline_registers.registers[0][22] ));
 sky130_fd_sc_hd__dfxtp_1 _14477_ (.CLK(clknet_leaf_220_clk),
    .D(_01102_),
    .Q(\core_pipeline.pipeline_registers.registers[0][23] ));
 sky130_fd_sc_hd__dfxtp_1 _14478_ (.CLK(clknet_leaf_227_clk),
    .D(_01103_),
    .Q(\core_pipeline.pipeline_registers.registers[0][24] ));
 sky130_fd_sc_hd__dfxtp_1 _14479_ (.CLK(clknet_leaf_18_clk),
    .D(_01104_),
    .Q(\core_pipeline.pipeline_registers.registers[0][25] ));
 sky130_fd_sc_hd__dfxtp_1 _14480_ (.CLK(clknet_leaf_47_clk),
    .D(_01105_),
    .Q(\core_pipeline.pipeline_registers.registers[0][26] ));
 sky130_fd_sc_hd__dfxtp_1 _14481_ (.CLK(clknet_leaf_171_clk),
    .D(_01106_),
    .Q(\core_pipeline.pipeline_registers.registers[0][27] ));
 sky130_fd_sc_hd__dfxtp_1 _14482_ (.CLK(clknet_leaf_185_clk),
    .D(_01107_),
    .Q(\core_pipeline.pipeline_registers.registers[0][28] ));
 sky130_fd_sc_hd__dfxtp_1 _14483_ (.CLK(clknet_leaf_161_clk),
    .D(_01108_),
    .Q(\core_pipeline.pipeline_registers.registers[0][29] ));
 sky130_fd_sc_hd__dfxtp_1 _14484_ (.CLK(clknet_leaf_209_clk),
    .D(_01109_),
    .Q(\core_pipeline.pipeline_registers.registers[0][30] ));
 sky130_fd_sc_hd__dfxtp_1 _14485_ (.CLK(clknet_leaf_172_clk),
    .D(_01110_),
    .Q(\core_pipeline.pipeline_registers.registers[0][31] ));
 sky130_fd_sc_hd__dfxtp_1 _14486_ (.CLK(clknet_leaf_140_clk),
    .D(_01111_),
    .Q(\core_pipeline.pipeline_csr.mtimecmp[32] ));
 sky130_fd_sc_hd__dfxtp_2 _14487_ (.CLK(clknet_leaf_139_clk),
    .D(_01112_),
    .Q(\core_pipeline.pipeline_csr.mtimecmp[33] ));
 sky130_fd_sc_hd__dfxtp_1 _14488_ (.CLK(clknet_leaf_139_clk),
    .D(_01113_),
    .Q(\core_pipeline.pipeline_csr.mtimecmp[34] ));
 sky130_fd_sc_hd__dfxtp_2 _14489_ (.CLK(clknet_leaf_143_clk),
    .D(_01114_),
    .Q(\core_pipeline.pipeline_csr.mtimecmp[35] ));
 sky130_fd_sc_hd__dfxtp_2 _14490_ (.CLK(clknet_leaf_143_clk),
    .D(_01115_),
    .Q(\core_pipeline.pipeline_csr.mtimecmp[36] ));
 sky130_fd_sc_hd__dfxtp_2 _14491_ (.CLK(clknet_leaf_143_clk),
    .D(_01116_),
    .Q(\core_pipeline.pipeline_csr.mtimecmp[37] ));
 sky130_fd_sc_hd__dfxtp_1 _14492_ (.CLK(clknet_leaf_144_clk),
    .D(_01117_),
    .Q(\core_pipeline.pipeline_csr.mtimecmp[38] ));
 sky130_fd_sc_hd__dfxtp_1 _14493_ (.CLK(clknet_leaf_145_clk),
    .D(_01118_),
    .Q(\core_pipeline.pipeline_csr.mtimecmp[39] ));
 sky130_fd_sc_hd__dfxtp_1 _14494_ (.CLK(clknet_leaf_118_clk),
    .D(_01119_),
    .Q(\core_pipeline.pipeline_csr.mtimecmp[40] ));
 sky130_fd_sc_hd__dfxtp_1 _14495_ (.CLK(clknet_leaf_119_clk),
    .D(_01120_),
    .Q(\core_pipeline.pipeline_csr.mtimecmp[41] ));
 sky130_fd_sc_hd__dfxtp_1 _14496_ (.CLK(clknet_leaf_117_clk),
    .D(_01121_),
    .Q(\core_pipeline.pipeline_csr.mtimecmp[42] ));
 sky130_fd_sc_hd__dfxtp_2 _14497_ (.CLK(clknet_leaf_144_clk),
    .D(_01122_),
    .Q(\core_pipeline.pipeline_csr.mtimecmp[43] ));
 sky130_fd_sc_hd__dfxtp_2 _14498_ (.CLK(clknet_leaf_114_clk),
    .D(_01123_),
    .Q(\core_pipeline.pipeline_csr.mtimecmp[44] ));
 sky130_fd_sc_hd__dfxtp_2 _14499_ (.CLK(clknet_leaf_114_clk),
    .D(_01124_),
    .Q(\core_pipeline.pipeline_csr.mtimecmp[45] ));
 sky130_fd_sc_hd__dfxtp_1 _14500_ (.CLK(clknet_leaf_121_clk),
    .D(_01125_),
    .Q(\core_pipeline.pipeline_csr.mtimecmp[46] ));
 sky130_fd_sc_hd__dfxtp_1 _14501_ (.CLK(clknet_leaf_121_clk),
    .D(_01126_),
    .Q(\core_pipeline.pipeline_csr.mtimecmp[47] ));
 sky130_fd_sc_hd__dfxtp_1 _14502_ (.CLK(clknet_leaf_124_clk),
    .D(_01127_),
    .Q(\core_pipeline.pipeline_csr.mtimecmp[48] ));
 sky130_fd_sc_hd__dfxtp_1 _14503_ (.CLK(clknet_leaf_124_clk),
    .D(_01128_),
    .Q(\core_pipeline.pipeline_csr.mtimecmp[49] ));
 sky130_fd_sc_hd__dfxtp_1 _14504_ (.CLK(clknet_leaf_123_clk),
    .D(_01129_),
    .Q(\core_pipeline.pipeline_csr.mtimecmp[50] ));
 sky130_fd_sc_hd__dfxtp_1 _14505_ (.CLK(clknet_leaf_120_clk),
    .D(_01130_),
    .Q(\core_pipeline.pipeline_csr.mtimecmp[51] ));
 sky130_fd_sc_hd__dfxtp_1 _14506_ (.CLK(clknet_leaf_126_clk),
    .D(_01131_),
    .Q(\core_pipeline.pipeline_csr.mtimecmp[52] ));
 sky130_fd_sc_hd__dfxtp_1 _14507_ (.CLK(clknet_leaf_129_clk),
    .D(_01132_),
    .Q(\core_pipeline.pipeline_csr.mtimecmp[53] ));
 sky130_fd_sc_hd__dfxtp_1 _14508_ (.CLK(clknet_leaf_129_clk),
    .D(_01133_),
    .Q(\core_pipeline.pipeline_csr.mtimecmp[54] ));
 sky130_fd_sc_hd__dfxtp_1 _14509_ (.CLK(clknet_leaf_129_clk),
    .D(_01134_),
    .Q(\core_pipeline.pipeline_csr.mtimecmp[55] ));
 sky130_fd_sc_hd__dfxtp_2 _14510_ (.CLK(clknet_leaf_129_clk),
    .D(_01135_),
    .Q(\core_pipeline.pipeline_csr.mtimecmp[56] ));
 sky130_fd_sc_hd__dfxtp_1 _14511_ (.CLK(clknet_leaf_128_clk),
    .D(_01136_),
    .Q(\core_pipeline.pipeline_csr.mtimecmp[57] ));
 sky130_fd_sc_hd__dfxtp_1 _14512_ (.CLK(clknet_leaf_132_clk),
    .D(_01137_),
    .Q(\core_pipeline.pipeline_csr.mtimecmp[58] ));
 sky130_fd_sc_hd__dfxtp_1 _14513_ (.CLK(clknet_leaf_134_clk),
    .D(_01138_),
    .Q(\core_pipeline.pipeline_csr.mtimecmp[59] ));
 sky130_fd_sc_hd__dfxtp_1 _14514_ (.CLK(clknet_leaf_133_clk),
    .D(_01139_),
    .Q(\core_pipeline.pipeline_csr.mtimecmp[60] ));
 sky130_fd_sc_hd__dfxtp_1 _14515_ (.CLK(clknet_leaf_133_clk),
    .D(_01140_),
    .Q(\core_pipeline.pipeline_csr.mtimecmp[61] ));
 sky130_fd_sc_hd__dfxtp_1 _14516_ (.CLK(clknet_leaf_137_clk),
    .D(_01141_),
    .Q(\core_pipeline.pipeline_csr.mtimecmp[62] ));
 sky130_fd_sc_hd__dfxtp_1 _14517_ (.CLK(clknet_leaf_137_clk),
    .D(_01142_),
    .Q(\core_pipeline.pipeline_csr.mtimecmp[63] ));
 sky130_fd_sc_hd__dfxtp_1 _14518_ (.CLK(clknet_leaf_251_clk),
    .D(_01143_),
    .Q(\core_pipeline.pipeline_registers.registers[20][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14519_ (.CLK(clknet_leaf_161_clk),
    .D(_01144_),
    .Q(\core_pipeline.pipeline_registers.registers[20][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14520_ (.CLK(clknet_leaf_199_clk),
    .D(_01145_),
    .Q(\core_pipeline.pipeline_registers.registers[20][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14521_ (.CLK(clknet_leaf_236_clk),
    .D(_01146_),
    .Q(\core_pipeline.pipeline_registers.registers[20][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14522_ (.CLK(clknet_leaf_250_clk),
    .D(_01147_),
    .Q(\core_pipeline.pipeline_registers.registers[20][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14523_ (.CLK(clknet_leaf_202_clk),
    .D(_01148_),
    .Q(\core_pipeline.pipeline_registers.registers[20][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14524_ (.CLK(clknet_leaf_206_clk),
    .D(_01149_),
    .Q(\core_pipeline.pipeline_registers.registers[20][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14525_ (.CLK(clknet_leaf_233_clk),
    .D(_01150_),
    .Q(\core_pipeline.pipeline_registers.registers[20][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14526_ (.CLK(clknet_leaf_242_clk),
    .D(_01151_),
    .Q(\core_pipeline.pipeline_registers.registers[20][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14527_ (.CLK(clknet_leaf_6_clk),
    .D(_01152_),
    .Q(\core_pipeline.pipeline_registers.registers[20][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14528_ (.CLK(clknet_leaf_10_clk),
    .D(_01153_),
    .Q(\core_pipeline.pipeline_registers.registers[20][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14529_ (.CLK(clknet_leaf_249_clk),
    .D(_01154_),
    .Q(\core_pipeline.pipeline_registers.registers[20][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14530_ (.CLK(clknet_leaf_231_clk),
    .D(_01155_),
    .Q(\core_pipeline.pipeline_registers.registers[20][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14531_ (.CLK(clknet_leaf_9_clk),
    .D(_01156_),
    .Q(\core_pipeline.pipeline_registers.registers[20][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14532_ (.CLK(clknet_leaf_10_clk),
    .D(_01157_),
    .Q(\core_pipeline.pipeline_registers.registers[20][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14533_ (.CLK(clknet_leaf_21_clk),
    .D(_01158_),
    .Q(\core_pipeline.pipeline_registers.registers[20][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14534_ (.CLK(clknet_leaf_246_clk),
    .D(_01159_),
    .Q(\core_pipeline.pipeline_registers.registers[20][16] ));
 sky130_fd_sc_hd__dfxtp_1 _14535_ (.CLK(clknet_leaf_163_clk),
    .D(_01160_),
    .Q(\core_pipeline.pipeline_registers.registers[20][17] ));
 sky130_fd_sc_hd__dfxtp_1 _14536_ (.CLK(clknet_leaf_179_clk),
    .D(_01161_),
    .Q(\core_pipeline.pipeline_registers.registers[20][18] ));
 sky130_fd_sc_hd__dfxtp_1 _14537_ (.CLK(clknet_leaf_193_clk),
    .D(_01162_),
    .Q(\core_pipeline.pipeline_registers.registers[20][19] ));
 sky130_fd_sc_hd__dfxtp_1 _14538_ (.CLK(clknet_leaf_187_clk),
    .D(_01163_),
    .Q(\core_pipeline.pipeline_registers.registers[20][20] ));
 sky130_fd_sc_hd__dfxtp_1 _14539_ (.CLK(clknet_leaf_169_clk),
    .D(_01164_),
    .Q(\core_pipeline.pipeline_registers.registers[20][21] ));
 sky130_fd_sc_hd__dfxtp_1 _14540_ (.CLK(clknet_leaf_202_clk),
    .D(_01165_),
    .Q(\core_pipeline.pipeline_registers.registers[20][22] ));
 sky130_fd_sc_hd__dfxtp_1 _14541_ (.CLK(clknet_leaf_209_clk),
    .D(_01166_),
    .Q(\core_pipeline.pipeline_registers.registers[20][23] ));
 sky130_fd_sc_hd__dfxtp_1 _14542_ (.CLK(clknet_leaf_226_clk),
    .D(_01167_),
    .Q(\core_pipeline.pipeline_registers.registers[20][24] ));
 sky130_fd_sc_hd__dfxtp_1 _14543_ (.CLK(clknet_leaf_10_clk),
    .D(_01168_),
    .Q(\core_pipeline.pipeline_registers.registers[20][25] ));
 sky130_fd_sc_hd__dfxtp_1 _14544_ (.CLK(clknet_leaf_22_clk),
    .D(_01169_),
    .Q(\core_pipeline.pipeline_registers.registers[20][26] ));
 sky130_fd_sc_hd__dfxtp_1 _14545_ (.CLK(clknet_leaf_169_clk),
    .D(_01170_),
    .Q(\core_pipeline.pipeline_registers.registers[20][27] ));
 sky130_fd_sc_hd__dfxtp_1 _14546_ (.CLK(clknet_leaf_183_clk),
    .D(_01171_),
    .Q(\core_pipeline.pipeline_registers.registers[20][28] ));
 sky130_fd_sc_hd__dfxtp_1 _14547_ (.CLK(clknet_leaf_212_clk),
    .D(_01172_),
    .Q(\core_pipeline.pipeline_registers.registers[20][29] ));
 sky130_fd_sc_hd__dfxtp_1 _14548_ (.CLK(clknet_leaf_209_clk),
    .D(_01173_),
    .Q(\core_pipeline.pipeline_registers.registers[20][30] ));
 sky130_fd_sc_hd__dfxtp_1 _14549_ (.CLK(clknet_leaf_177_clk),
    .D(_01174_),
    .Q(\core_pipeline.pipeline_registers.registers[20][31] ));
 sky130_fd_sc_hd__dfxtp_1 _14550_ (.CLK(clknet_leaf_255_clk),
    .D(_01175_),
    .Q(\core_pipeline.pipeline_registers.registers[11][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14551_ (.CLK(clknet_leaf_159_clk),
    .D(_01176_),
    .Q(\core_pipeline.pipeline_registers.registers[11][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14552_ (.CLK(clknet_leaf_192_clk),
    .D(_01177_),
    .Q(\core_pipeline.pipeline_registers.registers[11][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14553_ (.CLK(clknet_leaf_246_clk),
    .D(_01178_),
    .Q(\core_pipeline.pipeline_registers.registers[11][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14554_ (.CLK(clknet_leaf_256_clk),
    .D(_01179_),
    .Q(\core_pipeline.pipeline_registers.registers[11][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14555_ (.CLK(clknet_leaf_201_clk),
    .D(_01180_),
    .Q(\core_pipeline.pipeline_registers.registers[11][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14556_ (.CLK(clknet_leaf_240_clk),
    .D(_01181_),
    .Q(\core_pipeline.pipeline_registers.registers[11][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14557_ (.CLK(clknet_leaf_2_clk),
    .D(_01182_),
    .Q(\core_pipeline.pipeline_registers.registers[11][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14558_ (.CLK(clknet_leaf_240_clk),
    .D(_01183_),
    .Q(\core_pipeline.pipeline_registers.registers[11][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14559_ (.CLK(clknet_leaf_11_clk),
    .D(_01184_),
    .Q(\core_pipeline.pipeline_registers.registers[11][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14560_ (.CLK(clknet_leaf_14_clk),
    .D(_01185_),
    .Q(\core_pipeline.pipeline_registers.registers[11][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14561_ (.CLK(clknet_leaf_2_clk),
    .D(_01186_),
    .Q(\core_pipeline.pipeline_registers.registers[11][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14562_ (.CLK(clknet_leaf_248_clk),
    .D(_01187_),
    .Q(\core_pipeline.pipeline_registers.registers[11][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14563_ (.CLK(clknet_leaf_11_clk),
    .D(_01188_),
    .Q(\core_pipeline.pipeline_registers.registers[11][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14564_ (.CLK(clknet_leaf_15_clk),
    .D(_01189_),
    .Q(\core_pipeline.pipeline_registers.registers[11][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14565_ (.CLK(clknet_leaf_20_clk),
    .D(_01190_),
    .Q(\core_pipeline.pipeline_registers.registers[11][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14566_ (.CLK(clknet_leaf_252_clk),
    .D(_01191_),
    .Q(\core_pipeline.pipeline_registers.registers[11][16] ));
 sky130_fd_sc_hd__dfxtp_1 _14567_ (.CLK(clknet_leaf_213_clk),
    .D(_01192_),
    .Q(\core_pipeline.pipeline_registers.registers[11][17] ));
 sky130_fd_sc_hd__dfxtp_1 _14568_ (.CLK(clknet_leaf_186_clk),
    .D(_01193_),
    .Q(\core_pipeline.pipeline_registers.registers[11][18] ));
 sky130_fd_sc_hd__dfxtp_1 _14569_ (.CLK(clknet_leaf_191_clk),
    .D(_01194_),
    .Q(\core_pipeline.pipeline_registers.registers[11][19] ));
 sky130_fd_sc_hd__dfxtp_1 _14570_ (.CLK(clknet_leaf_189_clk),
    .D(_01195_),
    .Q(\core_pipeline.pipeline_registers.registers[11][20] ));
 sky130_fd_sc_hd__dfxtp_1 _14571_ (.CLK(clknet_leaf_173_clk),
    .D(_01196_),
    .Q(\core_pipeline.pipeline_registers.registers[11][21] ));
 sky130_fd_sc_hd__dfxtp_1 _14572_ (.CLK(clknet_leaf_204_clk),
    .D(_01197_),
    .Q(\core_pipeline.pipeline_registers.registers[11][22] ));
 sky130_fd_sc_hd__dfxtp_1 _14573_ (.CLK(clknet_leaf_218_clk),
    .D(_01198_),
    .Q(\core_pipeline.pipeline_registers.registers[11][23] ));
 sky130_fd_sc_hd__dfxtp_1 _14574_ (.CLK(clknet_leaf_235_clk),
    .D(_01199_),
    .Q(\core_pipeline.pipeline_registers.registers[11][24] ));
 sky130_fd_sc_hd__dfxtp_1 _14575_ (.CLK(clknet_leaf_12_clk),
    .D(_01200_),
    .Q(\core_pipeline.pipeline_registers.registers[11][25] ));
 sky130_fd_sc_hd__dfxtp_1 _14576_ (.CLK(clknet_leaf_17_clk),
    .D(_01201_),
    .Q(\core_pipeline.pipeline_registers.registers[11][26] ));
 sky130_fd_sc_hd__dfxtp_1 _14577_ (.CLK(clknet_leaf_139_clk),
    .D(_01202_),
    .Q(\core_pipeline.pipeline_registers.registers[11][27] ));
 sky130_fd_sc_hd__dfxtp_1 _14578_ (.CLK(clknet_leaf_184_clk),
    .D(_01203_),
    .Q(\core_pipeline.pipeline_registers.registers[11][28] ));
 sky130_fd_sc_hd__dfxtp_1 _14579_ (.CLK(clknet_leaf_214_clk),
    .D(_01204_),
    .Q(\core_pipeline.pipeline_registers.registers[11][29] ));
 sky130_fd_sc_hd__dfxtp_1 _14580_ (.CLK(clknet_leaf_236_clk),
    .D(_01205_),
    .Q(\core_pipeline.pipeline_registers.registers[11][30] ));
 sky130_fd_sc_hd__dfxtp_1 _14581_ (.CLK(clknet_leaf_177_clk),
    .D(_01206_),
    .Q(\core_pipeline.pipeline_registers.registers[11][31] ));
 sky130_fd_sc_hd__dfxtp_2 _14582_ (.CLK(clknet_leaf_35_clk),
    .D(_00000_),
    .Q(\core_pipeline.pipeline_decode.alu_select_a_out[2] ));
 sky130_fd_sc_hd__dfxtp_1 _14583_ (.CLK(clknet_leaf_92_clk),
    .D(_01207_),
    .Q(\core_pipeline.fetch_to_decode_instruction[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14584_ (.CLK(clknet_leaf_222_clk),
    .D(_01208_),
    .Q(\core_pipeline.fetch_to_decode_instruction[1] ));
 sky130_fd_sc_hd__dfxtp_1 _14585_ (.CLK(clknet_leaf_34_clk),
    .D(_01209_),
    .Q(\core_pipeline.fetch_to_decode_instruction[2] ));
 sky130_fd_sc_hd__dfxtp_2 _14586_ (.CLK(clknet_leaf_34_clk),
    .D(_01210_),
    .Q(\core_pipeline.fetch_to_decode_instruction[3] ));
 sky130_fd_sc_hd__dfxtp_4 _14587_ (.CLK(clknet_leaf_89_clk),
    .D(_01211_),
    .Q(\core_pipeline.fetch_to_decode_instruction[4] ));
 sky130_fd_sc_hd__dfxtp_2 _14588_ (.CLK(clknet_leaf_33_clk),
    .D(_01212_),
    .Q(\core_pipeline.fetch_to_decode_instruction[5] ));
 sky130_fd_sc_hd__dfxtp_2 _14589_ (.CLK(clknet_leaf_33_clk),
    .D(_01213_),
    .Q(\core_pipeline.fetch_to_decode_instruction[6] ));
 sky130_fd_sc_hd__dfxtp_2 _14590_ (.CLK(clknet_leaf_33_clk),
    .D(_01214_),
    .Q(\core_pipeline.fetch_to_decode_instruction[7] ));
 sky130_fd_sc_hd__dfxtp_2 _14591_ (.CLK(clknet_leaf_222_clk),
    .D(_01215_),
    .Q(\core_pipeline.fetch_to_decode_instruction[8] ));
 sky130_fd_sc_hd__dfxtp_2 _14592_ (.CLK(clknet_leaf_153_clk),
    .D(_01216_),
    .Q(\core_pipeline.fetch_to_decode_instruction[9] ));
 sky130_fd_sc_hd__dfxtp_2 _14593_ (.CLK(clknet_leaf_92_clk),
    .D(_01217_),
    .Q(\core_pipeline.fetch_to_decode_instruction[10] ));
 sky130_fd_sc_hd__dfxtp_2 _14594_ (.CLK(clknet_leaf_93_clk),
    .D(_01218_),
    .Q(\core_pipeline.fetch_to_decode_instruction[11] ));
 sky130_fd_sc_hd__dfxtp_4 _14595_ (.CLK(clknet_leaf_223_clk),
    .D(_01219_),
    .Q(\core_pipeline.fetch_to_decode_instruction[12] ));
 sky130_fd_sc_hd__dfxtp_4 _14596_ (.CLK(clknet_leaf_223_clk),
    .D(_01220_),
    .Q(\core_pipeline.fetch_to_decode_instruction[13] ));
 sky130_fd_sc_hd__dfxtp_4 _14597_ (.CLK(clknet_leaf_88_clk),
    .D(_01221_),
    .Q(\core_pipeline.fetch_to_decode_instruction[14] ));
 sky130_fd_sc_hd__dfxtp_4 _14598_ (.CLK(clknet_leaf_36_clk),
    .D(_01222_),
    .Q(\core_pipeline.decode_to_regfile_rs1_address[0] ));
 sky130_fd_sc_hd__dfxtp_4 _14599_ (.CLK(clknet_leaf_100_clk),
    .D(_01223_),
    .Q(\core_pipeline.decode_to_regfile_rs1_address[1] ));
 sky130_fd_sc_hd__dfxtp_4 _14600_ (.CLK(clknet_leaf_87_clk),
    .D(_01224_),
    .Q(\core_pipeline.decode_to_regfile_rs1_address[2] ));
 sky130_fd_sc_hd__dfxtp_4 _14601_ (.CLK(clknet_leaf_223_clk),
    .D(_01225_),
    .Q(\core_pipeline.decode_to_regfile_rs1_address[3] ));
 sky130_fd_sc_hd__dfxtp_1 _14602_ (.CLK(clknet_leaf_88_clk),
    .D(_01226_),
    .Q(\core_pipeline.decode_to_regfile_rs1_address[4] ));
 sky130_fd_sc_hd__dfxtp_1 _14603_ (.CLK(clknet_leaf_95_clk),
    .D(_01227_),
    .Q(\core_pipeline.decode_to_csr_read_address[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14604_ (.CLK(clknet_leaf_39_clk),
    .D(_01228_),
    .Q(\core_pipeline.decode_to_csr_read_address[1] ));
 sky130_fd_sc_hd__dfxtp_4 _14605_ (.CLK(clknet_leaf_41_clk),
    .D(_01229_),
    .Q(\core_pipeline.decode_to_csr_read_address[2] ));
 sky130_fd_sc_hd__dfxtp_4 _14606_ (.CLK(clknet_leaf_159_clk),
    .D(_01230_),
    .Q(\core_pipeline.decode_to_csr_read_address[3] ));
 sky130_fd_sc_hd__dfxtp_4 _14607_ (.CLK(clknet_leaf_100_clk),
    .D(_01231_),
    .Q(\core_pipeline.decode_to_csr_read_address[4] ));
 sky130_fd_sc_hd__dfxtp_4 _14608_ (.CLK(clknet_leaf_146_clk),
    .D(_01232_),
    .Q(\core_pipeline.decode_to_csr_read_address[5] ));
 sky130_fd_sc_hd__dfxtp_4 _14609_ (.CLK(clknet_leaf_158_clk),
    .D(_01233_),
    .Q(\core_pipeline.decode_to_csr_read_address[6] ));
 sky130_fd_sc_hd__dfxtp_4 _14610_ (.CLK(clknet_leaf_30_clk),
    .D(_01234_),
    .Q(\core_pipeline.decode_to_csr_read_address[7] ));
 sky130_fd_sc_hd__dfxtp_4 _14611_ (.CLK(clknet_leaf_158_clk),
    .D(_01235_),
    .Q(\core_pipeline.decode_to_csr_read_address[8] ));
 sky130_fd_sc_hd__dfxtp_4 _14612_ (.CLK(clknet_leaf_33_clk),
    .D(_01236_),
    .Q(\core_pipeline.decode_to_csr_read_address[9] ));
 sky130_fd_sc_hd__dfxtp_4 _14613_ (.CLK(clknet_leaf_158_clk),
    .D(_01237_),
    .Q(\core_pipeline.decode_to_csr_read_address[10] ));
 sky130_fd_sc_hd__dfxtp_4 _14614_ (.CLK(clknet_leaf_89_clk),
    .D(_01238_),
    .Q(\core_pipeline.decode_to_csr_read_address[11] ));
 sky130_fd_sc_hd__dfxtp_1 _14615_ (.CLK(clknet_leaf_151_clk),
    .D(_01239_),
    .Q(\core_pipeline.memory_to_writeback_pc[2] ));
 sky130_fd_sc_hd__dfxtp_1 _14616_ (.CLK(clknet_leaf_93_clk),
    .D(_01240_),
    .Q(\core_pipeline.memory_to_writeback_pc[3] ));
 sky130_fd_sc_hd__dfxtp_1 _14617_ (.CLK(clknet_leaf_40_clk),
    .D(_01241_),
    .Q(\core_pipeline.memory_to_writeback_pc[4] ));
 sky130_fd_sc_hd__dfxtp_1 _14618_ (.CLK(clknet_leaf_35_clk),
    .D(_01242_),
    .Q(\core_pipeline.memory_to_writeback_pc[5] ));
 sky130_fd_sc_hd__dfxtp_1 _14619_ (.CLK(clknet_leaf_88_clk),
    .D(_01243_),
    .Q(\core_pipeline.memory_to_writeback_pc[6] ));
 sky130_fd_sc_hd__dfxtp_1 _14620_ (.CLK(clknet_leaf_97_clk),
    .D(_01244_),
    .Q(\core_pipeline.memory_to_writeback_pc[7] ));
 sky130_fd_sc_hd__dfxtp_1 _14621_ (.CLK(clknet_leaf_80_clk),
    .D(_01245_),
    .Q(\core_pipeline.memory_to_writeback_pc[8] ));
 sky130_fd_sc_hd__dfxtp_1 _14622_ (.CLK(clknet_leaf_74_clk),
    .D(_01246_),
    .Q(\core_pipeline.memory_to_writeback_pc[9] ));
 sky130_fd_sc_hd__dfxtp_1 _14623_ (.CLK(clknet_leaf_77_clk),
    .D(_01247_),
    .Q(\core_pipeline.memory_to_writeback_pc[10] ));
 sky130_fd_sc_hd__dfxtp_1 _14624_ (.CLK(clknet_leaf_72_clk),
    .D(_01248_),
    .Q(\core_pipeline.memory_to_writeback_pc[11] ));
 sky130_fd_sc_hd__dfxtp_1 _14625_ (.CLK(clknet_leaf_72_clk),
    .D(_01249_),
    .Q(\core_pipeline.memory_to_writeback_pc[12] ));
 sky130_fd_sc_hd__dfxtp_1 _14626_ (.CLK(clknet_leaf_72_clk),
    .D(_01250_),
    .Q(\core_pipeline.memory_to_writeback_pc[13] ));
 sky130_fd_sc_hd__dfxtp_1 _14627_ (.CLK(clknet_leaf_76_clk),
    .D(_01251_),
    .Q(\core_pipeline.memory_to_writeback_pc[14] ));
 sky130_fd_sc_hd__dfxtp_1 _14628_ (.CLK(clknet_leaf_71_clk),
    .D(_01252_),
    .Q(\core_pipeline.memory_to_writeback_pc[15] ));
 sky130_fd_sc_hd__dfxtp_1 _14629_ (.CLK(clknet_leaf_72_clk),
    .D(_01253_),
    .Q(\core_pipeline.memory_to_writeback_pc[16] ));
 sky130_fd_sc_hd__dfxtp_1 _14630_ (.CLK(clknet_leaf_109_clk),
    .D(_01254_),
    .Q(\core_pipeline.memory_to_writeback_pc[17] ));
 sky130_fd_sc_hd__dfxtp_1 _14631_ (.CLK(clknet_leaf_111_clk),
    .D(_01255_),
    .Q(\core_pipeline.memory_to_writeback_pc[18] ));
 sky130_fd_sc_hd__dfxtp_1 _14632_ (.CLK(clknet_leaf_107_clk),
    .D(_01256_),
    .Q(\core_pipeline.memory_to_writeback_pc[19] ));
 sky130_fd_sc_hd__dfxtp_1 _14633_ (.CLK(clknet_leaf_115_clk),
    .D(_01257_),
    .Q(\core_pipeline.memory_to_writeback_pc[20] ));
 sky130_fd_sc_hd__dfxtp_1 _14634_ (.CLK(clknet_leaf_101_clk),
    .D(_01258_),
    .Q(\core_pipeline.memory_to_writeback_pc[21] ));
 sky130_fd_sc_hd__dfxtp_1 _14635_ (.CLK(clknet_leaf_101_clk),
    .D(_01259_),
    .Q(\core_pipeline.memory_to_writeback_pc[22] ));
 sky130_fd_sc_hd__dfxtp_1 _14636_ (.CLK(clknet_leaf_105_clk),
    .D(_01260_),
    .Q(\core_pipeline.memory_to_writeback_pc[23] ));
 sky130_fd_sc_hd__dfxtp_1 _14637_ (.CLK(clknet_leaf_82_clk),
    .D(_01261_),
    .Q(\core_pipeline.memory_to_writeback_pc[24] ));
 sky130_fd_sc_hd__dfxtp_1 _14638_ (.CLK(clknet_leaf_79_clk),
    .D(_01262_),
    .Q(\core_pipeline.memory_to_writeback_pc[25] ));
 sky130_fd_sc_hd__dfxtp_1 _14639_ (.CLK(clknet_leaf_96_clk),
    .D(_01263_),
    .Q(\core_pipeline.memory_to_writeback_pc[26] ));
 sky130_fd_sc_hd__dfxtp_1 _14640_ (.CLK(clknet_leaf_99_clk),
    .D(_01264_),
    .Q(\core_pipeline.memory_to_writeback_pc[27] ));
 sky130_fd_sc_hd__dfxtp_1 _14641_ (.CLK(clknet_leaf_98_clk),
    .D(_01265_),
    .Q(\core_pipeline.memory_to_writeback_pc[28] ));
 sky130_fd_sc_hd__dfxtp_1 _14642_ (.CLK(clknet_leaf_96_clk),
    .D(_01266_),
    .Q(\core_pipeline.memory_to_writeback_pc[29] ));
 sky130_fd_sc_hd__dfxtp_1 _14643_ (.CLK(clknet_leaf_89_clk),
    .D(_01267_),
    .Q(\core_pipeline.memory_to_writeback_pc[30] ));
 sky130_fd_sc_hd__dfxtp_1 _14644_ (.CLK(clknet_leaf_147_clk),
    .D(_01268_),
    .Q(\core_pipeline.memory_to_writeback_pc[31] ));
 sky130_fd_sc_hd__dfxtp_1 _14645_ (.CLK(clknet_leaf_90_clk),
    .D(_01269_),
    .Q(\core_pipeline.memory_to_writeback_next_pc[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14646_ (.CLK(clknet_leaf_153_clk),
    .D(_01270_),
    .Q(\core_pipeline.memory_to_writeback_next_pc[1] ));
 sky130_fd_sc_hd__dfxtp_1 _14647_ (.CLK(clknet_leaf_150_clk),
    .D(_01271_),
    .Q(\core_pipeline.memory_to_writeback_next_pc[2] ));
 sky130_fd_sc_hd__dfxtp_1 _14648_ (.CLK(clknet_leaf_151_clk),
    .D(_01272_),
    .Q(\core_pipeline.memory_to_writeback_next_pc[3] ));
 sky130_fd_sc_hd__dfxtp_1 _14649_ (.CLK(clknet_leaf_89_clk),
    .D(_01273_),
    .Q(\core_pipeline.memory_to_writeback_next_pc[4] ));
 sky130_fd_sc_hd__dfxtp_1 _14650_ (.CLK(clknet_leaf_93_clk),
    .D(_01274_),
    .Q(\core_pipeline.memory_to_writeback_next_pc[5] ));
 sky130_fd_sc_hd__dfxtp_1 _14651_ (.CLK(clknet_leaf_87_clk),
    .D(_01275_),
    .Q(\core_pipeline.memory_to_writeback_next_pc[6] ));
 sky130_fd_sc_hd__dfxtp_1 _14652_ (.CLK(clknet_leaf_97_clk),
    .D(_01276_),
    .Q(\core_pipeline.memory_to_writeback_next_pc[7] ));
 sky130_fd_sc_hd__dfxtp_1 _14653_ (.CLK(clknet_leaf_80_clk),
    .D(_01277_),
    .Q(\core_pipeline.memory_to_writeback_next_pc[8] ));
 sky130_fd_sc_hd__dfxtp_1 _14654_ (.CLK(clknet_leaf_77_clk),
    .D(_01278_),
    .Q(\core_pipeline.memory_to_writeback_next_pc[9] ));
 sky130_fd_sc_hd__dfxtp_1 _14655_ (.CLK(clknet_leaf_77_clk),
    .D(_01279_),
    .Q(\core_pipeline.memory_to_writeback_next_pc[10] ));
 sky130_fd_sc_hd__dfxtp_1 _14656_ (.CLK(clknet_leaf_74_clk),
    .D(_01280_),
    .Q(\core_pipeline.memory_to_writeback_next_pc[11] ));
 sky130_fd_sc_hd__dfxtp_1 _14657_ (.CLK(clknet_leaf_74_clk),
    .D(_01281_),
    .Q(\core_pipeline.memory_to_writeback_next_pc[12] ));
 sky130_fd_sc_hd__dfxtp_1 _14658_ (.CLK(clknet_leaf_75_clk),
    .D(_01282_),
    .Q(\core_pipeline.memory_to_writeback_next_pc[13] ));
 sky130_fd_sc_hd__dfxtp_1 _14659_ (.CLK(clknet_leaf_108_clk),
    .D(_01283_),
    .Q(\core_pipeline.memory_to_writeback_next_pc[14] ));
 sky130_fd_sc_hd__dfxtp_1 _14660_ (.CLK(clknet_leaf_75_clk),
    .D(_01284_),
    .Q(\core_pipeline.memory_to_writeback_next_pc[15] ));
 sky130_fd_sc_hd__dfxtp_1 _14661_ (.CLK(clknet_leaf_74_clk),
    .D(_01285_),
    .Q(\core_pipeline.memory_to_writeback_next_pc[16] ));
 sky130_fd_sc_hd__dfxtp_1 _14662_ (.CLK(clknet_leaf_109_clk),
    .D(_01286_),
    .Q(\core_pipeline.memory_to_writeback_next_pc[17] ));
 sky130_fd_sc_hd__dfxtp_1 _14663_ (.CLK(clknet_leaf_109_clk),
    .D(_01287_),
    .Q(\core_pipeline.memory_to_writeback_next_pc[18] ));
 sky130_fd_sc_hd__dfxtp_1 _14664_ (.CLK(clknet_leaf_110_clk),
    .D(_01288_),
    .Q(\core_pipeline.memory_to_writeback_next_pc[19] ));
 sky130_fd_sc_hd__dfxtp_1 _14665_ (.CLK(clknet_leaf_115_clk),
    .D(_01289_),
    .Q(\core_pipeline.memory_to_writeback_next_pc[20] ));
 sky130_fd_sc_hd__dfxtp_1 _14666_ (.CLK(clknet_leaf_100_clk),
    .D(_01290_),
    .Q(\core_pipeline.memory_to_writeback_next_pc[21] ));
 sky130_fd_sc_hd__dfxtp_1 _14667_ (.CLK(clknet_leaf_102_clk),
    .D(_01291_),
    .Q(\core_pipeline.memory_to_writeback_next_pc[22] ));
 sky130_fd_sc_hd__dfxtp_1 _14668_ (.CLK(clknet_leaf_105_clk),
    .D(_01292_),
    .Q(\core_pipeline.memory_to_writeback_next_pc[23] ));
 sky130_fd_sc_hd__dfxtp_1 _14669_ (.CLK(clknet_leaf_79_clk),
    .D(_01293_),
    .Q(\core_pipeline.memory_to_writeback_next_pc[24] ));
 sky130_fd_sc_hd__dfxtp_1 _14670_ (.CLK(clknet_leaf_79_clk),
    .D(_01294_),
    .Q(\core_pipeline.memory_to_writeback_next_pc[25] ));
 sky130_fd_sc_hd__dfxtp_1 _14671_ (.CLK(clknet_leaf_107_clk),
    .D(_01295_),
    .Q(\core_pipeline.memory_to_writeback_next_pc[26] ));
 sky130_fd_sc_hd__dfxtp_1 _14672_ (.CLK(clknet_leaf_102_clk),
    .D(_01296_),
    .Q(\core_pipeline.memory_to_writeback_next_pc[27] ));
 sky130_fd_sc_hd__dfxtp_1 _14673_ (.CLK(clknet_leaf_99_clk),
    .D(_01297_),
    .Q(\core_pipeline.memory_to_writeback_next_pc[28] ));
 sky130_fd_sc_hd__dfxtp_1 _14674_ (.CLK(clknet_leaf_96_clk),
    .D(_01298_),
    .Q(\core_pipeline.memory_to_writeback_next_pc[29] ));
 sky130_fd_sc_hd__dfxtp_1 _14675_ (.CLK(clknet_leaf_95_clk),
    .D(_01299_),
    .Q(\core_pipeline.memory_to_writeback_next_pc[30] ));
 sky130_fd_sc_hd__dfxtp_1 _14676_ (.CLK(clknet_leaf_98_clk),
    .D(_01300_),
    .Q(\core_pipeline.memory_to_writeback_next_pc[31] ));
 sky130_fd_sc_hd__dfxtp_1 _14677_ (.CLK(clknet_leaf_38_clk),
    .D(_01301_),
    .Q(\core_pipeline.memory_to_writeback_csr_data[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14678_ (.CLK(clknet_leaf_92_clk),
    .D(_01302_),
    .Q(\core_pipeline.memory_to_writeback_csr_data[1] ));
 sky130_fd_sc_hd__dfxtp_1 _14679_ (.CLK(clknet_leaf_151_clk),
    .D(_01303_),
    .Q(\core_pipeline.memory_to_writeback_csr_data[2] ));
 sky130_fd_sc_hd__dfxtp_1 _14680_ (.CLK(clknet_leaf_36_clk),
    .D(_01304_),
    .Q(\core_pipeline.memory_to_writeback_csr_data[3] ));
 sky130_fd_sc_hd__dfxtp_1 _14681_ (.CLK(clknet_leaf_40_clk),
    .D(_01305_),
    .Q(\core_pipeline.memory_to_writeback_csr_data[4] ));
 sky130_fd_sc_hd__dfxtp_1 _14682_ (.CLK(clknet_leaf_93_clk),
    .D(_01306_),
    .Q(\core_pipeline.memory_to_writeback_csr_data[5] ));
 sky130_fd_sc_hd__dfxtp_1 _14683_ (.CLK(clknet_leaf_88_clk),
    .D(_01307_),
    .Q(\core_pipeline.memory_to_writeback_csr_data[6] ));
 sky130_fd_sc_hd__dfxtp_1 _14684_ (.CLK(clknet_leaf_40_clk),
    .D(_01308_),
    .Q(\core_pipeline.memory_to_writeback_csr_data[7] ));
 sky130_fd_sc_hd__dfxtp_1 _14685_ (.CLK(clknet_leaf_81_clk),
    .D(_01309_),
    .Q(\core_pipeline.memory_to_writeback_csr_data[8] ));
 sky130_fd_sc_hd__dfxtp_1 _14686_ (.CLK(clknet_leaf_81_clk),
    .D(_01310_),
    .Q(\core_pipeline.memory_to_writeback_csr_data[9] ));
 sky130_fd_sc_hd__dfxtp_1 _14687_ (.CLK(clknet_leaf_82_clk),
    .D(_01311_),
    .Q(\core_pipeline.memory_to_writeback_csr_data[10] ));
 sky130_fd_sc_hd__dfxtp_1 _14688_ (.CLK(clknet_leaf_86_clk),
    .D(_01312_),
    .Q(\core_pipeline.memory_to_writeback_csr_data[11] ));
 sky130_fd_sc_hd__dfxtp_1 _14689_ (.CLK(clknet_leaf_73_clk),
    .D(_01313_),
    .Q(\core_pipeline.memory_to_writeback_csr_data[12] ));
 sky130_fd_sc_hd__dfxtp_1 _14690_ (.CLK(clknet_leaf_78_clk),
    .D(_01314_),
    .Q(\core_pipeline.memory_to_writeback_csr_data[13] ));
 sky130_fd_sc_hd__dfxtp_1 _14691_ (.CLK(clknet_leaf_73_clk),
    .D(_01315_),
    .Q(\core_pipeline.memory_to_writeback_csr_data[14] ));
 sky130_fd_sc_hd__dfxtp_1 _14692_ (.CLK(clknet_leaf_78_clk),
    .D(_01316_),
    .Q(\core_pipeline.memory_to_writeback_csr_data[15] ));
 sky130_fd_sc_hd__dfxtp_1 _14693_ (.CLK(clknet_leaf_78_clk),
    .D(_01317_),
    .Q(\core_pipeline.memory_to_writeback_csr_data[16] ));
 sky130_fd_sc_hd__dfxtp_1 _14694_ (.CLK(clknet_leaf_106_clk),
    .D(_01318_),
    .Q(\core_pipeline.memory_to_writeback_csr_data[17] ));
 sky130_fd_sc_hd__dfxtp_1 _14695_ (.CLK(clknet_leaf_102_clk),
    .D(_01319_),
    .Q(\core_pipeline.memory_to_writeback_csr_data[18] ));
 sky130_fd_sc_hd__dfxtp_1 _14696_ (.CLK(clknet_leaf_106_clk),
    .D(_01320_),
    .Q(\core_pipeline.memory_to_writeback_csr_data[19] ));
 sky130_fd_sc_hd__dfxtp_1 _14697_ (.CLK(clknet_leaf_102_clk),
    .D(_01321_),
    .Q(\core_pipeline.memory_to_writeback_csr_data[20] ));
 sky130_fd_sc_hd__dfxtp_1 _14698_ (.CLK(clknet_leaf_103_clk),
    .D(_01322_),
    .Q(\core_pipeline.memory_to_writeback_csr_data[21] ));
 sky130_fd_sc_hd__dfxtp_1 _14699_ (.CLK(clknet_leaf_103_clk),
    .D(_01323_),
    .Q(\core_pipeline.memory_to_writeback_csr_data[22] ));
 sky130_fd_sc_hd__dfxtp_1 _14700_ (.CLK(clknet_leaf_104_clk),
    .D(_01324_),
    .Q(\core_pipeline.memory_to_writeback_csr_data[23] ));
 sky130_fd_sc_hd__dfxtp_1 _14701_ (.CLK(clknet_leaf_80_clk),
    .D(_01325_),
    .Q(\core_pipeline.memory_to_writeback_csr_data[24] ));
 sky130_fd_sc_hd__dfxtp_1 _14702_ (.CLK(clknet_leaf_81_clk),
    .D(_01326_),
    .Q(\core_pipeline.memory_to_writeback_csr_data[25] ));
 sky130_fd_sc_hd__dfxtp_1 _14703_ (.CLK(clknet_leaf_86_clk),
    .D(_01327_),
    .Q(\core_pipeline.memory_to_writeback_csr_data[26] ));
 sky130_fd_sc_hd__dfxtp_1 _14704_ (.CLK(clknet_leaf_99_clk),
    .D(_01328_),
    .Q(\core_pipeline.memory_to_writeback_csr_data[27] ));
 sky130_fd_sc_hd__dfxtp_1 _14705_ (.CLK(clknet_leaf_97_clk),
    .D(_01329_),
    .Q(\core_pipeline.memory_to_writeback_csr_data[28] ));
 sky130_fd_sc_hd__dfxtp_1 _14706_ (.CLK(clknet_leaf_95_clk),
    .D(_01330_),
    .Q(\core_pipeline.memory_to_writeback_csr_data[29] ));
 sky130_fd_sc_hd__dfxtp_1 _14707_ (.CLK(clknet_leaf_88_clk),
    .D(_01331_),
    .Q(\core_pipeline.memory_to_writeback_csr_data[30] ));
 sky130_fd_sc_hd__dfxtp_1 _14708_ (.CLK(clknet_leaf_94_clk),
    .D(_01332_),
    .Q(\core_pipeline.memory_to_writeback_csr_data[31] ));
 sky130_fd_sc_hd__dfxtp_2 _14709_ (.CLK(clknet_leaf_149_clk),
    .D(_01333_),
    .Q(\core_pipeline.memory_to_writeback_csr_write ));
 sky130_fd_sc_hd__dfxtp_4 _14710_ (.CLK(clknet_leaf_94_clk),
    .D(_01334_),
    .Q(\core_pipeline.memory_to_writeback_write_select[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14711_ (.CLK(clknet_leaf_222_clk),
    .D(_01335_),
    .Q(\core_pipeline.memory_to_writeback_write_select[1] ));
 sky130_fd_sc_hd__dfxtp_4 _14712_ (.CLK(clknet_leaf_156_clk),
    .D(_01336_),
    .Q(\core_pipeline.memory_to_writeback_rd_address[0] ));
 sky130_fd_sc_hd__dfxtp_4 _14713_ (.CLK(clknet_leaf_156_clk),
    .D(_01337_),
    .Q(\core_pipeline.memory_to_writeback_rd_address[1] ));
 sky130_fd_sc_hd__dfxtp_4 _14714_ (.CLK(clknet_leaf_156_clk),
    .D(_01338_),
    .Q(\core_pipeline.memory_to_writeback_rd_address[2] ));
 sky130_fd_sc_hd__dfxtp_4 _14715_ (.CLK(clknet_leaf_155_clk),
    .D(_01339_),
    .Q(\core_pipeline.memory_to_writeback_rd_address[3] ));
 sky130_fd_sc_hd__dfxtp_4 _14716_ (.CLK(clknet_leaf_155_clk),
    .D(_01340_),
    .Q(\core_pipeline.memory_to_writeback_rd_address[4] ));
 sky130_fd_sc_hd__dfxtp_4 _14717_ (.CLK(clknet_leaf_140_clk),
    .D(_01341_),
    .Q(\core_pipeline.memory_to_writeback_csr_address[0] ));
 sky130_fd_sc_hd__dfxtp_4 _14718_ (.CLK(clknet_leaf_139_clk),
    .D(_01342_),
    .Q(\core_pipeline.memory_to_writeback_csr_address[1] ));
 sky130_fd_sc_hd__dfxtp_1 _14719_ (.CLK(clknet_leaf_141_clk),
    .D(_01343_),
    .Q(\core_pipeline.memory_to_writeback_csr_address[2] ));
 sky130_fd_sc_hd__dfxtp_1 _14720_ (.CLK(clknet_leaf_140_clk),
    .D(_01344_),
    .Q(\core_pipeline.memory_to_writeback_csr_address[3] ));
 sky130_fd_sc_hd__dfxtp_2 _14721_ (.CLK(clknet_leaf_168_clk),
    .D(_01345_),
    .Q(\core_pipeline.memory_to_writeback_csr_address[4] ));
 sky130_fd_sc_hd__dfxtp_2 _14722_ (.CLK(clknet_leaf_167_clk),
    .D(_01346_),
    .Q(\core_pipeline.memory_to_writeback_csr_address[5] ));
 sky130_fd_sc_hd__dfxtp_2 _14723_ (.CLK(clknet_leaf_141_clk),
    .D(_01347_),
    .Q(\core_pipeline.memory_to_writeback_csr_address[6] ));
 sky130_fd_sc_hd__dfxtp_2 _14724_ (.CLK(clknet_leaf_141_clk),
    .D(_01348_),
    .Q(\core_pipeline.memory_to_writeback_csr_address[7] ));
 sky130_fd_sc_hd__dfxtp_1 _14725_ (.CLK(clknet_leaf_167_clk),
    .D(_01349_),
    .Q(\core_pipeline.memory_to_writeback_csr_address[8] ));
 sky130_fd_sc_hd__dfxtp_1 _14726_ (.CLK(clknet_leaf_167_clk),
    .D(_01350_),
    .Q(\core_pipeline.memory_to_writeback_csr_address[9] ));
 sky130_fd_sc_hd__dfxtp_1 _14727_ (.CLK(clknet_leaf_167_clk),
    .D(_01351_),
    .Q(\core_pipeline.memory_to_writeback_csr_address[10] ));
 sky130_fd_sc_hd__dfxtp_1 _14728_ (.CLK(clknet_leaf_167_clk),
    .D(_01352_),
    .Q(\core_pipeline.memory_to_writeback_csr_address[11] ));
 sky130_fd_sc_hd__dfxtp_4 _14729_ (.CLK(clknet_leaf_149_clk),
    .D(_01353_),
    .Q(\core_pipeline.memory_to_writeback_mret ));
 sky130_fd_sc_hd__dfxtp_4 _14730_ (.CLK(clknet_leaf_150_clk),
    .D(_00040_),
    .Q(\core_pipeline.memory_to_writeback_valid ));
 sky130_fd_sc_hd__dfxtp_1 _14731_ (.CLK(clknet_leaf_43_clk),
    .D(_01354_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_sltu[0] ));
 sky130_fd_sc_hd__dfxtp_2 _14732_ (.CLK(clknet_leaf_149_clk),
    .D(_01355_),
    .Q(\core_pipeline.memory_to_writeback_exception ));
 sky130_fd_sc_hd__dfxtp_1 _14733_ (.CLK(clknet_leaf_151_clk),
    .D(_01356_),
    .Q(\core_pipeline.memory_to_writeback_wfi ));
 sky130_fd_sc_hd__dfxtp_4 _14734_ (.CLK(clknet_leaf_38_clk),
    .D(_01357_),
    .Q(\core_pipeline.memory_to_writeback_alu_data[0] ));
 sky130_fd_sc_hd__dfxtp_4 _14735_ (.CLK(clknet_leaf_92_clk),
    .D(_01358_),
    .Q(\core_pipeline.memory_to_writeback_alu_data[1] ));
 sky130_fd_sc_hd__dfxtp_4 _14736_ (.CLK(clknet_leaf_151_clk),
    .D(_01359_),
    .Q(\core_pipeline.memory_to_writeback_alu_data[2] ));
 sky130_fd_sc_hd__dfxtp_4 _14737_ (.CLK(clknet_leaf_40_clk),
    .D(_01360_),
    .Q(\core_pipeline.memory_to_writeback_alu_data[3] ));
 sky130_fd_sc_hd__dfxtp_4 _14738_ (.CLK(clknet_leaf_39_clk),
    .D(_01361_),
    .Q(\core_pipeline.memory_to_writeback_alu_data[4] ));
 sky130_fd_sc_hd__dfxtp_4 _14739_ (.CLK(clknet_leaf_93_clk),
    .D(_01362_),
    .Q(\core_pipeline.memory_to_writeback_alu_data[5] ));
 sky130_fd_sc_hd__dfxtp_4 _14740_ (.CLK(clknet_leaf_88_clk),
    .D(_01363_),
    .Q(\core_pipeline.memory_to_writeback_alu_data[6] ));
 sky130_fd_sc_hd__dfxtp_4 _14741_ (.CLK(clknet_leaf_40_clk),
    .D(_01364_),
    .Q(\core_pipeline.memory_to_writeback_alu_data[7] ));
 sky130_fd_sc_hd__dfxtp_4 _14742_ (.CLK(clknet_leaf_81_clk),
    .D(_01365_),
    .Q(\core_pipeline.memory_to_writeback_alu_data[8] ));
 sky130_fd_sc_hd__dfxtp_4 _14743_ (.CLK(clknet_leaf_73_clk),
    .D(_01366_),
    .Q(\core_pipeline.memory_to_writeback_alu_data[9] ));
 sky130_fd_sc_hd__dfxtp_4 _14744_ (.CLK(clknet_leaf_78_clk),
    .D(_01367_),
    .Q(\core_pipeline.memory_to_writeback_alu_data[10] ));
 sky130_fd_sc_hd__dfxtp_4 _14745_ (.CLK(clknet_leaf_73_clk),
    .D(_01368_),
    .Q(\core_pipeline.memory_to_writeback_alu_data[11] ));
 sky130_fd_sc_hd__dfxtp_4 _14746_ (.CLK(clknet_leaf_73_clk),
    .D(_01369_),
    .Q(\core_pipeline.memory_to_writeback_alu_data[12] ));
 sky130_fd_sc_hd__dfxtp_4 _14747_ (.CLK(clknet_leaf_70_clk),
    .D(_01370_),
    .Q(\core_pipeline.memory_to_writeback_alu_data[13] ));
 sky130_fd_sc_hd__dfxtp_4 _14748_ (.CLK(clknet_leaf_70_clk),
    .D(_01371_),
    .Q(\core_pipeline.memory_to_writeback_alu_data[14] ));
 sky130_fd_sc_hd__dfxtp_4 _14749_ (.CLK(clknet_leaf_78_clk),
    .D(_01372_),
    .Q(\core_pipeline.memory_to_writeback_alu_data[15] ));
 sky130_fd_sc_hd__dfxtp_4 _14750_ (.CLK(clknet_leaf_78_clk),
    .D(_01373_),
    .Q(\core_pipeline.memory_to_writeback_alu_data[16] ));
 sky130_fd_sc_hd__dfxtp_4 _14751_ (.CLK(clknet_leaf_106_clk),
    .D(_01374_),
    .Q(\core_pipeline.memory_to_writeback_alu_data[17] ));
 sky130_fd_sc_hd__dfxtp_4 _14752_ (.CLK(clknet_leaf_102_clk),
    .D(_01375_),
    .Q(\core_pipeline.memory_to_writeback_alu_data[18] ));
 sky130_fd_sc_hd__dfxtp_4 _14753_ (.CLK(clknet_leaf_115_clk),
    .D(_01376_),
    .Q(\core_pipeline.memory_to_writeback_alu_data[19] ));
 sky130_fd_sc_hd__dfxtp_4 _14754_ (.CLK(clknet_leaf_102_clk),
    .D(_01377_),
    .Q(\core_pipeline.memory_to_writeback_alu_data[20] ));
 sky130_fd_sc_hd__dfxtp_4 _14755_ (.CLK(clknet_leaf_103_clk),
    .D(_01378_),
    .Q(\core_pipeline.memory_to_writeback_alu_data[21] ));
 sky130_fd_sc_hd__dfxtp_4 _14756_ (.CLK(clknet_leaf_103_clk),
    .D(_01379_),
    .Q(\core_pipeline.memory_to_writeback_alu_data[22] ));
 sky130_fd_sc_hd__dfxtp_4 _14757_ (.CLK(clknet_leaf_104_clk),
    .D(_01380_),
    .Q(\core_pipeline.memory_to_writeback_alu_data[23] ));
 sky130_fd_sc_hd__dfxtp_4 _14758_ (.CLK(clknet_leaf_81_clk),
    .D(_01381_),
    .Q(\core_pipeline.memory_to_writeback_alu_data[24] ));
 sky130_fd_sc_hd__dfxtp_4 _14759_ (.CLK(clknet_leaf_81_clk),
    .D(_01382_),
    .Q(\core_pipeline.memory_to_writeback_alu_data[25] ));
 sky130_fd_sc_hd__dfxtp_4 _14760_ (.CLK(clknet_leaf_83_clk),
    .D(_01383_),
    .Q(\core_pipeline.memory_to_writeback_alu_data[26] ));
 sky130_fd_sc_hd__dfxtp_4 _14761_ (.CLK(clknet_leaf_101_clk),
    .D(_01384_),
    .Q(\core_pipeline.memory_to_writeback_alu_data[27] ));
 sky130_fd_sc_hd__dfxtp_4 _14762_ (.CLK(clknet_leaf_98_clk),
    .D(_01385_),
    .Q(\core_pipeline.memory_to_writeback_alu_data[28] ));
 sky130_fd_sc_hd__dfxtp_4 _14763_ (.CLK(clknet_leaf_97_clk),
    .D(_01386_),
    .Q(\core_pipeline.memory_to_writeback_alu_data[29] ));
 sky130_fd_sc_hd__dfxtp_4 _14764_ (.CLK(clknet_leaf_88_clk),
    .D(_01387_),
    .Q(\core_pipeline.memory_to_writeback_alu_data[30] ));
 sky130_fd_sc_hd__dfxtp_4 _14765_ (.CLK(clknet_leaf_94_clk),
    .D(_01388_),
    .Q(\core_pipeline.memory_to_writeback_alu_data[31] ));
 sky130_fd_sc_hd__dfxtp_4 _14766_ (.CLK(clknet_leaf_35_clk),
    .D(_00001_),
    .Q(\core_pipeline.pipeline_decode.alu_select_b_out[1] ));
 sky130_fd_sc_hd__dfxtp_4 _14767_ (.CLK(clknet_leaf_35_clk),
    .D(_00002_),
    .Q(\core_pipeline.pipeline_decode.alu_select_b_out[2] ));
 sky130_fd_sc_hd__dfxtp_1 _14768_ (.CLK(clknet_leaf_151_clk),
    .D(_01389_),
    .Q(\core_pipeline.execute_to_memory_pc[2] ));
 sky130_fd_sc_hd__dfxtp_1 _14769_ (.CLK(clknet_leaf_93_clk),
    .D(_01390_),
    .Q(\core_pipeline.execute_to_memory_pc[3] ));
 sky130_fd_sc_hd__dfxtp_1 _14770_ (.CLK(clknet_leaf_39_clk),
    .D(_01391_),
    .Q(\core_pipeline.execute_to_memory_pc[4] ));
 sky130_fd_sc_hd__dfxtp_1 _14771_ (.CLK(clknet_leaf_36_clk),
    .D(_01392_),
    .Q(\core_pipeline.execute_to_memory_pc[5] ));
 sky130_fd_sc_hd__dfxtp_1 _14772_ (.CLK(clknet_leaf_40_clk),
    .D(_01393_),
    .Q(\core_pipeline.execute_to_memory_pc[6] ));
 sky130_fd_sc_hd__dfxtp_1 _14773_ (.CLK(clknet_leaf_94_clk),
    .D(_01394_),
    .Q(\core_pipeline.execute_to_memory_pc[7] ));
 sky130_fd_sc_hd__dfxtp_1 _14774_ (.CLK(clknet_leaf_80_clk),
    .D(_01395_),
    .Q(\core_pipeline.execute_to_memory_pc[8] ));
 sky130_fd_sc_hd__dfxtp_1 _14775_ (.CLK(clknet_leaf_73_clk),
    .D(_01396_),
    .Q(\core_pipeline.execute_to_memory_pc[9] ));
 sky130_fd_sc_hd__dfxtp_1 _14776_ (.CLK(clknet_leaf_77_clk),
    .D(_01397_),
    .Q(\core_pipeline.execute_to_memory_pc[10] ));
 sky130_fd_sc_hd__dfxtp_1 _14777_ (.CLK(clknet_leaf_71_clk),
    .D(_01398_),
    .Q(\core_pipeline.execute_to_memory_pc[11] ));
 sky130_fd_sc_hd__dfxtp_1 _14778_ (.CLK(clknet_leaf_72_clk),
    .D(_01399_),
    .Q(\core_pipeline.execute_to_memory_pc[12] ));
 sky130_fd_sc_hd__dfxtp_1 _14779_ (.CLK(clknet_leaf_72_clk),
    .D(_01400_),
    .Q(\core_pipeline.execute_to_memory_pc[13] ));
 sky130_fd_sc_hd__dfxtp_1 _14780_ (.CLK(clknet_leaf_76_clk),
    .D(_01401_),
    .Q(\core_pipeline.execute_to_memory_pc[14] ));
 sky130_fd_sc_hd__dfxtp_1 _14781_ (.CLK(clknet_leaf_71_clk),
    .D(_01402_),
    .Q(\core_pipeline.execute_to_memory_pc[15] ));
 sky130_fd_sc_hd__dfxtp_1 _14782_ (.CLK(clknet_leaf_72_clk),
    .D(_01403_),
    .Q(\core_pipeline.execute_to_memory_pc[16] ));
 sky130_fd_sc_hd__dfxtp_1 _14783_ (.CLK(clknet_leaf_109_clk),
    .D(_01404_),
    .Q(\core_pipeline.execute_to_memory_pc[17] ));
 sky130_fd_sc_hd__dfxtp_1 _14784_ (.CLK(clknet_leaf_111_clk),
    .D(_01405_),
    .Q(\core_pipeline.execute_to_memory_pc[18] ));
 sky130_fd_sc_hd__dfxtp_1 _14785_ (.CLK(clknet_leaf_107_clk),
    .D(_01406_),
    .Q(\core_pipeline.execute_to_memory_pc[19] ));
 sky130_fd_sc_hd__dfxtp_1 _14786_ (.CLK(clknet_leaf_116_clk),
    .D(_01407_),
    .Q(\core_pipeline.execute_to_memory_pc[20] ));
 sky130_fd_sc_hd__dfxtp_1 _14787_ (.CLK(clknet_leaf_101_clk),
    .D(_01408_),
    .Q(\core_pipeline.execute_to_memory_pc[21] ));
 sky130_fd_sc_hd__dfxtp_1 _14788_ (.CLK(clknet_leaf_101_clk),
    .D(_01409_),
    .Q(\core_pipeline.execute_to_memory_pc[22] ));
 sky130_fd_sc_hd__dfxtp_1 _14789_ (.CLK(clknet_leaf_105_clk),
    .D(_01410_),
    .Q(\core_pipeline.execute_to_memory_pc[23] ));
 sky130_fd_sc_hd__dfxtp_1 _14790_ (.CLK(clknet_leaf_82_clk),
    .D(_01411_),
    .Q(\core_pipeline.execute_to_memory_pc[24] ));
 sky130_fd_sc_hd__dfxtp_1 _14791_ (.CLK(clknet_leaf_79_clk),
    .D(_01412_),
    .Q(\core_pipeline.execute_to_memory_pc[25] ));
 sky130_fd_sc_hd__dfxtp_1 _14792_ (.CLK(clknet_leaf_96_clk),
    .D(_01413_),
    .Q(\core_pipeline.execute_to_memory_pc[26] ));
 sky130_fd_sc_hd__dfxtp_1 _14793_ (.CLK(clknet_leaf_99_clk),
    .D(_01414_),
    .Q(\core_pipeline.execute_to_memory_pc[27] ));
 sky130_fd_sc_hd__dfxtp_1 _14794_ (.CLK(clknet_leaf_98_clk),
    .D(_01415_),
    .Q(\core_pipeline.execute_to_memory_pc[28] ));
 sky130_fd_sc_hd__dfxtp_1 _14795_ (.CLK(clknet_leaf_87_clk),
    .D(_01416_),
    .Q(\core_pipeline.execute_to_memory_pc[29] ));
 sky130_fd_sc_hd__dfxtp_1 _14796_ (.CLK(clknet_leaf_85_clk),
    .D(_01417_),
    .Q(\core_pipeline.execute_to_memory_pc[30] ));
 sky130_fd_sc_hd__dfxtp_1 _14797_ (.CLK(clknet_leaf_147_clk),
    .D(_01418_),
    .Q(\core_pipeline.execute_to_memory_pc[31] ));
 sky130_fd_sc_hd__dfxtp_1 _14798_ (.CLK(clknet_leaf_35_clk),
    .D(_01419_),
    .Q(\core_pipeline.execute_to_memory_next_pc[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14799_ (.CLK(clknet_leaf_153_clk),
    .D(_01420_),
    .Q(\core_pipeline.execute_to_memory_next_pc[1] ));
 sky130_fd_sc_hd__dfxtp_1 _14800_ (.CLK(clknet_leaf_150_clk),
    .D(_01421_),
    .Q(\core_pipeline.execute_to_memory_next_pc[2] ));
 sky130_fd_sc_hd__dfxtp_1 _14801_ (.CLK(clknet_leaf_151_clk),
    .D(_01422_),
    .Q(\core_pipeline.execute_to_memory_next_pc[3] ));
 sky130_fd_sc_hd__dfxtp_1 _14802_ (.CLK(clknet_leaf_91_clk),
    .D(_01423_),
    .Q(\core_pipeline.execute_to_memory_next_pc[4] ));
 sky130_fd_sc_hd__dfxtp_1 _14803_ (.CLK(clknet_leaf_94_clk),
    .D(_01424_),
    .Q(\core_pipeline.execute_to_memory_next_pc[5] ));
 sky130_fd_sc_hd__dfxtp_1 _14804_ (.CLK(clknet_leaf_87_clk),
    .D(_01425_),
    .Q(\core_pipeline.execute_to_memory_next_pc[6] ));
 sky130_fd_sc_hd__dfxtp_1 _14805_ (.CLK(clknet_leaf_97_clk),
    .D(_01426_),
    .Q(\core_pipeline.execute_to_memory_next_pc[7] ));
 sky130_fd_sc_hd__dfxtp_1 _14806_ (.CLK(clknet_leaf_104_clk),
    .D(_01427_),
    .Q(\core_pipeline.execute_to_memory_next_pc[8] ));
 sky130_fd_sc_hd__dfxtp_1 _14807_ (.CLK(clknet_leaf_77_clk),
    .D(_01428_),
    .Q(\core_pipeline.execute_to_memory_next_pc[9] ));
 sky130_fd_sc_hd__dfxtp_1 _14808_ (.CLK(clknet_leaf_77_clk),
    .D(_01429_),
    .Q(\core_pipeline.execute_to_memory_next_pc[10] ));
 sky130_fd_sc_hd__dfxtp_1 _14809_ (.CLK(clknet_leaf_74_clk),
    .D(_01430_),
    .Q(\core_pipeline.execute_to_memory_next_pc[11] ));
 sky130_fd_sc_hd__dfxtp_1 _14810_ (.CLK(clknet_leaf_74_clk),
    .D(_01431_),
    .Q(\core_pipeline.execute_to_memory_next_pc[12] ));
 sky130_fd_sc_hd__dfxtp_1 _14811_ (.CLK(clknet_leaf_75_clk),
    .D(_01432_),
    .Q(\core_pipeline.execute_to_memory_next_pc[13] ));
 sky130_fd_sc_hd__dfxtp_1 _14812_ (.CLK(clknet_leaf_108_clk),
    .D(_01433_),
    .Q(\core_pipeline.execute_to_memory_next_pc[14] ));
 sky130_fd_sc_hd__dfxtp_1 _14813_ (.CLK(clknet_leaf_75_clk),
    .D(_01434_),
    .Q(\core_pipeline.execute_to_memory_next_pc[15] ));
 sky130_fd_sc_hd__dfxtp_1 _14814_ (.CLK(clknet_leaf_75_clk),
    .D(_01435_),
    .Q(\core_pipeline.execute_to_memory_next_pc[16] ));
 sky130_fd_sc_hd__dfxtp_1 _14815_ (.CLK(clknet_leaf_109_clk),
    .D(_01436_),
    .Q(\core_pipeline.execute_to_memory_next_pc[17] ));
 sky130_fd_sc_hd__dfxtp_1 _14816_ (.CLK(clknet_leaf_109_clk),
    .D(_01437_),
    .Q(\core_pipeline.execute_to_memory_next_pc[18] ));
 sky130_fd_sc_hd__dfxtp_1 _14817_ (.CLK(clknet_leaf_106_clk),
    .D(_01438_),
    .Q(\core_pipeline.execute_to_memory_next_pc[19] ));
 sky130_fd_sc_hd__dfxtp_1 _14818_ (.CLK(clknet_leaf_115_clk),
    .D(_01439_),
    .Q(\core_pipeline.execute_to_memory_next_pc[20] ));
 sky130_fd_sc_hd__dfxtp_1 _14819_ (.CLK(clknet_leaf_101_clk),
    .D(_01440_),
    .Q(\core_pipeline.execute_to_memory_next_pc[21] ));
 sky130_fd_sc_hd__dfxtp_1 _14820_ (.CLK(clknet_leaf_102_clk),
    .D(_01441_),
    .Q(\core_pipeline.execute_to_memory_next_pc[22] ));
 sky130_fd_sc_hd__dfxtp_1 _14821_ (.CLK(clknet_leaf_105_clk),
    .D(_01442_),
    .Q(\core_pipeline.execute_to_memory_next_pc[23] ));
 sky130_fd_sc_hd__dfxtp_1 _14822_ (.CLK(clknet_leaf_79_clk),
    .D(_01443_),
    .Q(\core_pipeline.execute_to_memory_next_pc[24] ));
 sky130_fd_sc_hd__dfxtp_1 _14823_ (.CLK(clknet_leaf_79_clk),
    .D(_01444_),
    .Q(\core_pipeline.execute_to_memory_next_pc[25] ));
 sky130_fd_sc_hd__dfxtp_1 _14824_ (.CLK(clknet_leaf_106_clk),
    .D(_01445_),
    .Q(\core_pipeline.execute_to_memory_next_pc[26] ));
 sky130_fd_sc_hd__dfxtp_1 _14825_ (.CLK(clknet_leaf_106_clk),
    .D(_01446_),
    .Q(\core_pipeline.execute_to_memory_next_pc[27] ));
 sky130_fd_sc_hd__dfxtp_1 _14826_ (.CLK(clknet_leaf_99_clk),
    .D(_01447_),
    .Q(\core_pipeline.execute_to_memory_next_pc[28] ));
 sky130_fd_sc_hd__dfxtp_1 _14827_ (.CLK(clknet_leaf_96_clk),
    .D(_01448_),
    .Q(\core_pipeline.execute_to_memory_next_pc[29] ));
 sky130_fd_sc_hd__dfxtp_1 _14828_ (.CLK(clknet_leaf_95_clk),
    .D(_01449_),
    .Q(\core_pipeline.execute_to_memory_next_pc[30] ));
 sky130_fd_sc_hd__dfxtp_1 _14829_ (.CLK(clknet_leaf_98_clk),
    .D(_01450_),
    .Q(\core_pipeline.execute_to_memory_next_pc[31] ));
 sky130_fd_sc_hd__dfxtp_4 _14830_ (.CLK(clknet_leaf_38_clk),
    .D(_01451_),
    .Q(\core_busio.mem_store_data[0] ));
 sky130_fd_sc_hd__dfxtp_2 _14831_ (.CLK(clknet_leaf_223_clk),
    .D(_01452_),
    .Q(\core_busio.mem_store_data[1] ));
 sky130_fd_sc_hd__dfxtp_2 _14832_ (.CLK(clknet_leaf_223_clk),
    .D(_01453_),
    .Q(\core_busio.mem_store_data[2] ));
 sky130_fd_sc_hd__dfxtp_2 _14833_ (.CLK(clknet_leaf_26_clk),
    .D(_01454_),
    .Q(\core_busio.mem_store_data[3] ));
 sky130_fd_sc_hd__dfxtp_2 _14834_ (.CLK(clknet_leaf_27_clk),
    .D(_01455_),
    .Q(\core_busio.mem_store_data[4] ));
 sky130_fd_sc_hd__dfxtp_2 _14835_ (.CLK(clknet_leaf_223_clk),
    .D(_01456_),
    .Q(\core_busio.mem_store_data[5] ));
 sky130_fd_sc_hd__dfxtp_2 _14836_ (.CLK(clknet_leaf_223_clk),
    .D(_01457_),
    .Q(\core_busio.mem_store_data[6] ));
 sky130_fd_sc_hd__dfxtp_4 _14837_ (.CLK(clknet_leaf_30_clk),
    .D(_01458_),
    .Q(\core_busio.mem_store_data[7] ));
 sky130_fd_sc_hd__dfxtp_1 _14838_ (.CLK(clknet_leaf_26_clk),
    .D(_01459_),
    .Q(\core_busio.mem_store_data[8] ));
 sky130_fd_sc_hd__dfxtp_1 _14839_ (.CLK(clknet_leaf_27_clk),
    .D(_01460_),
    .Q(\core_busio.mem_store_data[9] ));
 sky130_fd_sc_hd__dfxtp_1 _14840_ (.CLK(clknet_leaf_28_clk),
    .D(_01461_),
    .Q(\core_busio.mem_store_data[10] ));
 sky130_fd_sc_hd__dfxtp_1 _14841_ (.CLK(clknet_leaf_27_clk),
    .D(_01462_),
    .Q(\core_busio.mem_store_data[11] ));
 sky130_fd_sc_hd__dfxtp_1 _14842_ (.CLK(clknet_leaf_27_clk),
    .D(_01463_),
    .Q(\core_busio.mem_store_data[12] ));
 sky130_fd_sc_hd__dfxtp_2 _14843_ (.CLK(clknet_leaf_39_clk),
    .D(_01464_),
    .Q(\core_busio.mem_store_data[13] ));
 sky130_fd_sc_hd__dfxtp_1 _14844_ (.CLK(clknet_leaf_26_clk),
    .D(_01465_),
    .Q(\core_busio.mem_store_data[14] ));
 sky130_fd_sc_hd__dfxtp_1 _14845_ (.CLK(clknet_leaf_39_clk),
    .D(_01466_),
    .Q(\core_busio.mem_store_data[15] ));
 sky130_fd_sc_hd__dfxtp_1 _14846_ (.CLK(clknet_leaf_228_clk),
    .D(_01467_),
    .Q(\core_busio.mem_store_data[16] ));
 sky130_fd_sc_hd__dfxtp_1 _14847_ (.CLK(clknet_leaf_223_clk),
    .D(_01468_),
    .Q(\core_busio.mem_store_data[17] ));
 sky130_fd_sc_hd__dfxtp_1 _14848_ (.CLK(clknet_leaf_30_clk),
    .D(_01469_),
    .Q(\core_busio.mem_store_data[18] ));
 sky130_fd_sc_hd__dfxtp_1 _14849_ (.CLK(clknet_leaf_31_clk),
    .D(_01470_),
    .Q(\core_busio.mem_store_data[19] ));
 sky130_fd_sc_hd__dfxtp_1 _14850_ (.CLK(clknet_leaf_224_clk),
    .D(_01471_),
    .Q(\core_busio.mem_store_data[20] ));
 sky130_fd_sc_hd__dfxtp_1 _14851_ (.CLK(clknet_leaf_90_clk),
    .D(_01472_),
    .Q(\core_busio.mem_store_data[21] ));
 sky130_fd_sc_hd__dfxtp_1 _14852_ (.CLK(clknet_leaf_224_clk),
    .D(_01473_),
    .Q(\core_busio.mem_store_data[22] ));
 sky130_fd_sc_hd__dfxtp_1 _14853_ (.CLK(clknet_leaf_35_clk),
    .D(_01474_),
    .Q(\core_busio.mem_store_data[23] ));
 sky130_fd_sc_hd__dfxtp_1 _14854_ (.CLK(clknet_leaf_227_clk),
    .D(_01475_),
    .Q(\core_busio.mem_store_data[24] ));
 sky130_fd_sc_hd__dfxtp_1 _14855_ (.CLK(clknet_leaf_31_clk),
    .D(_01476_),
    .Q(\core_busio.mem_store_data[25] ));
 sky130_fd_sc_hd__dfxtp_1 _14856_ (.CLK(clknet_leaf_31_clk),
    .D(_01477_),
    .Q(\core_busio.mem_store_data[26] ));
 sky130_fd_sc_hd__dfxtp_1 _14857_ (.CLK(clknet_leaf_31_clk),
    .D(_01478_),
    .Q(\core_busio.mem_store_data[27] ));
 sky130_fd_sc_hd__dfxtp_1 _14858_ (.CLK(clknet_leaf_224_clk),
    .D(_01479_),
    .Q(\core_busio.mem_store_data[28] ));
 sky130_fd_sc_hd__dfxtp_1 _14859_ (.CLK(clknet_leaf_91_clk),
    .D(_01480_),
    .Q(\core_busio.mem_store_data[29] ));
 sky130_fd_sc_hd__dfxtp_1 _14860_ (.CLK(clknet_leaf_224_clk),
    .D(_01481_),
    .Q(\core_busio.mem_store_data[30] ));
 sky130_fd_sc_hd__dfxtp_1 _14861_ (.CLK(clknet_leaf_35_clk),
    .D(_01482_),
    .Q(\core_busio.mem_store_data[31] ));
 sky130_fd_sc_hd__dfxtp_1 _14862_ (.CLK(clknet_leaf_38_clk),
    .D(_01483_),
    .Q(\core_pipeline.execute_to_memory_csr_data[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14863_ (.CLK(clknet_leaf_37_clk),
    .D(_01484_),
    .Q(\core_pipeline.execute_to_memory_csr_data[1] ));
 sky130_fd_sc_hd__dfxtp_1 _14864_ (.CLK(clknet_leaf_151_clk),
    .D(_01485_),
    .Q(\core_pipeline.execute_to_memory_csr_data[2] ));
 sky130_fd_sc_hd__dfxtp_1 _14865_ (.CLK(clknet_leaf_36_clk),
    .D(_01486_),
    .Q(\core_pipeline.execute_to_memory_csr_data[3] ));
 sky130_fd_sc_hd__dfxtp_1 _14866_ (.CLK(clknet_leaf_39_clk),
    .D(_01487_),
    .Q(\core_pipeline.execute_to_memory_csr_data[4] ));
 sky130_fd_sc_hd__dfxtp_1 _14867_ (.CLK(clknet_leaf_93_clk),
    .D(_01488_),
    .Q(\core_pipeline.execute_to_memory_csr_data[5] ));
 sky130_fd_sc_hd__dfxtp_1 _14868_ (.CLK(clknet_leaf_85_clk),
    .D(_01489_),
    .Q(\core_pipeline.execute_to_memory_csr_data[6] ));
 sky130_fd_sc_hd__dfxtp_1 _14869_ (.CLK(clknet_leaf_40_clk),
    .D(_01490_),
    .Q(\core_pipeline.execute_to_memory_csr_data[7] ));
 sky130_fd_sc_hd__dfxtp_1 _14870_ (.CLK(clknet_leaf_81_clk),
    .D(_01491_),
    .Q(\core_pipeline.execute_to_memory_csr_data[8] ));
 sky130_fd_sc_hd__dfxtp_1 _14871_ (.CLK(clknet_leaf_82_clk),
    .D(_01492_),
    .Q(\core_pipeline.execute_to_memory_csr_data[9] ));
 sky130_fd_sc_hd__dfxtp_1 _14872_ (.CLK(clknet_leaf_82_clk),
    .D(_01493_),
    .Q(\core_pipeline.execute_to_memory_csr_data[10] ));
 sky130_fd_sc_hd__dfxtp_1 _14873_ (.CLK(clknet_leaf_83_clk),
    .D(_01494_),
    .Q(\core_pipeline.execute_to_memory_csr_data[11] ));
 sky130_fd_sc_hd__dfxtp_1 _14874_ (.CLK(clknet_leaf_73_clk),
    .D(_01495_),
    .Q(\core_pipeline.execute_to_memory_csr_data[12] ));
 sky130_fd_sc_hd__dfxtp_2 _14875_ (.CLK(clknet_leaf_72_clk),
    .D(_01496_),
    .Q(\core_pipeline.execute_to_memory_csr_data[13] ));
 sky130_fd_sc_hd__dfxtp_1 _14876_ (.CLK(clknet_leaf_73_clk),
    .D(_01497_),
    .Q(\core_pipeline.execute_to_memory_csr_data[14] ));
 sky130_fd_sc_hd__dfxtp_1 _14877_ (.CLK(clknet_leaf_82_clk),
    .D(_01498_),
    .Q(\core_pipeline.execute_to_memory_csr_data[15] ));
 sky130_fd_sc_hd__dfxtp_1 _14878_ (.CLK(clknet_leaf_73_clk),
    .D(_01499_),
    .Q(\core_pipeline.execute_to_memory_csr_data[16] ));
 sky130_fd_sc_hd__dfxtp_1 _14879_ (.CLK(clknet_leaf_106_clk),
    .D(_01500_),
    .Q(\core_pipeline.execute_to_memory_csr_data[17] ));
 sky130_fd_sc_hd__dfxtp_1 _14880_ (.CLK(clknet_leaf_102_clk),
    .D(_01501_),
    .Q(\core_pipeline.execute_to_memory_csr_data[18] ));
 sky130_fd_sc_hd__dfxtp_1 _14881_ (.CLK(clknet_leaf_102_clk),
    .D(_01502_),
    .Q(\core_pipeline.execute_to_memory_csr_data[19] ));
 sky130_fd_sc_hd__dfxtp_1 _14882_ (.CLK(clknet_leaf_103_clk),
    .D(_01503_),
    .Q(\core_pipeline.execute_to_memory_csr_data[20] ));
 sky130_fd_sc_hd__dfxtp_1 _14883_ (.CLK(clknet_leaf_103_clk),
    .D(_01504_),
    .Q(\core_pipeline.execute_to_memory_csr_data[21] ));
 sky130_fd_sc_hd__dfxtp_1 _14884_ (.CLK(clknet_leaf_103_clk),
    .D(_01505_),
    .Q(\core_pipeline.execute_to_memory_csr_data[22] ));
 sky130_fd_sc_hd__dfxtp_1 _14885_ (.CLK(clknet_leaf_104_clk),
    .D(_01506_),
    .Q(\core_pipeline.execute_to_memory_csr_data[23] ));
 sky130_fd_sc_hd__dfxtp_1 _14886_ (.CLK(clknet_leaf_81_clk),
    .D(_01507_),
    .Q(\core_pipeline.execute_to_memory_csr_data[24] ));
 sky130_fd_sc_hd__dfxtp_1 _14887_ (.CLK(clknet_leaf_81_clk),
    .D(_01508_),
    .Q(\core_pipeline.execute_to_memory_csr_data[25] ));
 sky130_fd_sc_hd__dfxtp_1 _14888_ (.CLK(clknet_leaf_84_clk),
    .D(_01509_),
    .Q(\core_pipeline.execute_to_memory_csr_data[26] ));
 sky130_fd_sc_hd__dfxtp_1 _14889_ (.CLK(clknet_leaf_99_clk),
    .D(_01510_),
    .Q(\core_pipeline.execute_to_memory_csr_data[27] ));
 sky130_fd_sc_hd__dfxtp_1 _14890_ (.CLK(clknet_leaf_97_clk),
    .D(_01511_),
    .Q(\core_pipeline.execute_to_memory_csr_data[28] ));
 sky130_fd_sc_hd__dfxtp_1 _14891_ (.CLK(clknet_leaf_95_clk),
    .D(_01512_),
    .Q(\core_pipeline.execute_to_memory_csr_data[29] ));
 sky130_fd_sc_hd__dfxtp_1 _14892_ (.CLK(clknet_leaf_88_clk),
    .D(_01513_),
    .Q(\core_pipeline.execute_to_memory_csr_data[30] ));
 sky130_fd_sc_hd__dfxtp_1 _14893_ (.CLK(clknet_leaf_94_clk),
    .D(_01514_),
    .Q(\core_pipeline.execute_to_memory_csr_data[31] ));
 sky130_fd_sc_hd__dfxtp_1 _14894_ (.CLK(clknet_leaf_222_clk),
    .D(_01515_),
    .Q(\core_pipeline.execute_to_memory_jump ));
 sky130_fd_sc_hd__dfxtp_1 _14895_ (.CLK(clknet_leaf_222_clk),
    .D(_01516_),
    .Q(\core_pipeline.execute_to_memory_branch ));
 sky130_fd_sc_hd__dfxtp_1 _14896_ (.CLK(clknet_leaf_157_clk),
    .D(_01517_),
    .Q(\core_pipeline.execute_to_memory_csr_write ));
 sky130_fd_sc_hd__dfxtp_1 _14897_ (.CLK(clknet_leaf_92_clk),
    .D(_01518_),
    .Q(\core_pipeline.execute_to_memory_load ));
 sky130_fd_sc_hd__dfxtp_1 _14898_ (.CLK(clknet_leaf_92_clk),
    .D(_01519_),
    .Q(\core_pipeline.execute_to_memory_store ));
 sky130_fd_sc_hd__dfxtp_2 _14899_ (.CLK(clknet_leaf_223_clk),
    .D(_01520_),
    .Q(\core_busio.mem_size[0] ));
 sky130_fd_sc_hd__dfxtp_4 _14900_ (.CLK(clknet_leaf_223_clk),
    .D(_01521_),
    .Q(\core_busio.mem_size[1] ));
 sky130_fd_sc_hd__dfxtp_1 _14901_ (.CLK(clknet_leaf_92_clk),
    .D(_01522_),
    .Q(\core_busio.mem_signed ));
 sky130_fd_sc_hd__dfxtp_1 _14902_ (.CLK(clknet_leaf_154_clk),
    .D(_01523_),
    .Q(\core_pipeline.execute_to_memory_bypass_memory ));
 sky130_fd_sc_hd__dfxtp_4 _14903_ (.CLK(clknet_leaf_34_clk),
    .D(_01524_),
    .Q(\core_pipeline.execute_to_memory_write_select[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14904_ (.CLK(clknet_leaf_222_clk),
    .D(_01525_),
    .Q(\core_pipeline.execute_to_memory_write_select[1] ));
 sky130_fd_sc_hd__dfxtp_2 _14905_ (.CLK(clknet_leaf_221_clk),
    .D(_01526_),
    .Q(\core_pipeline.execute_to_memory_rd_address[0] ));
 sky130_fd_sc_hd__dfxtp_2 _14906_ (.CLK(clknet_leaf_154_clk),
    .D(_01527_),
    .Q(\core_pipeline.execute_to_memory_rd_address[1] ));
 sky130_fd_sc_hd__dfxtp_2 _14907_ (.CLK(clknet_leaf_221_clk),
    .D(_01528_),
    .Q(\core_pipeline.execute_to_memory_rd_address[2] ));
 sky130_fd_sc_hd__dfxtp_2 _14908_ (.CLK(clknet_leaf_221_clk),
    .D(_01529_),
    .Q(\core_pipeline.execute_to_memory_rd_address[3] ));
 sky130_fd_sc_hd__dfxtp_2 _14909_ (.CLK(clknet_leaf_221_clk),
    .D(_01530_),
    .Q(\core_pipeline.execute_to_memory_rd_address[4] ));
 sky130_fd_sc_hd__dfxtp_1 _14910_ (.CLK(clknet_leaf_138_clk),
    .D(_01531_),
    .Q(\core_pipeline.execute_to_memory_csr_address[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14911_ (.CLK(clknet_leaf_139_clk),
    .D(_01532_),
    .Q(\core_pipeline.execute_to_memory_csr_address[1] ));
 sky130_fd_sc_hd__dfxtp_1 _14912_ (.CLK(clknet_leaf_139_clk),
    .D(_01533_),
    .Q(\core_pipeline.execute_to_memory_csr_address[2] ));
 sky130_fd_sc_hd__dfxtp_1 _14913_ (.CLK(clknet_leaf_170_clk),
    .D(_01534_),
    .Q(\core_pipeline.execute_to_memory_csr_address[3] ));
 sky130_fd_sc_hd__dfxtp_1 _14914_ (.CLK(clknet_leaf_168_clk),
    .D(_01535_),
    .Q(\core_pipeline.execute_to_memory_csr_address[4] ));
 sky130_fd_sc_hd__dfxtp_1 _14915_ (.CLK(clknet_leaf_167_clk),
    .D(_01536_),
    .Q(\core_pipeline.execute_to_memory_csr_address[5] ));
 sky130_fd_sc_hd__dfxtp_1 _14916_ (.CLK(clknet_leaf_168_clk),
    .D(_01537_),
    .Q(\core_pipeline.execute_to_memory_csr_address[6] ));
 sky130_fd_sc_hd__dfxtp_1 _14917_ (.CLK(clknet_leaf_141_clk),
    .D(_01538_),
    .Q(\core_pipeline.execute_to_memory_csr_address[7] ));
 sky130_fd_sc_hd__dfxtp_1 _14918_ (.CLK(clknet_leaf_166_clk),
    .D(_01539_),
    .Q(\core_pipeline.execute_to_memory_csr_address[8] ));
 sky130_fd_sc_hd__dfxtp_1 _14919_ (.CLK(clknet_leaf_167_clk),
    .D(_01540_),
    .Q(\core_pipeline.execute_to_memory_csr_address[9] ));
 sky130_fd_sc_hd__dfxtp_1 _14920_ (.CLK(clknet_leaf_166_clk),
    .D(_01541_),
    .Q(\core_pipeline.execute_to_memory_csr_address[10] ));
 sky130_fd_sc_hd__dfxtp_1 _14921_ (.CLK(clknet_leaf_167_clk),
    .D(_01542_),
    .Q(\core_pipeline.execute_to_memory_csr_address[11] ));
 sky130_fd_sc_hd__dfxtp_1 _14922_ (.CLK(clknet_leaf_150_clk),
    .D(_01543_),
    .Q(\core_pipeline.execute_to_memory_mret ));
 sky130_fd_sc_hd__dfxtp_4 _14923_ (.CLK(clknet_leaf_157_clk),
    .D(_00038_),
    .Q(\core_pipeline.execute_to_memory_valid ));
 sky130_fd_sc_hd__dfxtp_4 _14924_ (.CLK(clknet_leaf_158_clk),
    .D(_01544_),
    .Q(\core_pipeline.execute_to_memory_exception ));
 sky130_fd_sc_hd__dfxtp_1 _14925_ (.CLK(clknet_leaf_32_clk),
    .D(_00039_),
    .Q(\core_pipeline.pipeline_execute.ex_cmp.quasi_result ));
 sky130_fd_sc_hd__dfxtp_1 _14926_ (.CLK(clknet_leaf_223_clk),
    .D(\core_pipeline.decode_to_execute_cmp_function[0] ),
    .Q(\core_pipeline.pipeline_execute.ex_cmp.negate ));
 sky130_fd_sc_hd__dfxtp_2 _14927_ (.CLK(clknet_leaf_41_clk),
    .D(\core_pipeline.decode_to_execute_alu_function[0] ),
    .Q(\core_pipeline.pipeline_execute.ex_alu.old_function[0] ));
 sky130_fd_sc_hd__dfxtp_2 _14928_ (.CLK(clknet_leaf_44_clk),
    .D(\core_pipeline.decode_to_execute_alu_function[1] ),
    .Q(\core_pipeline.pipeline_execute.ex_alu.old_function[1] ));
 sky130_fd_sc_hd__dfxtp_2 _14929_ (.CLK(clknet_leaf_44_clk),
    .D(\core_pipeline.decode_to_execute_alu_function[2] ),
    .Q(\core_pipeline.pipeline_execute.ex_alu.old_function[2] ));
 sky130_fd_sc_hd__dfxtp_1 _14930_ (.CLK(clknet_leaf_45_clk),
    .D(_01545_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_or[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14931_ (.CLK(clknet_leaf_48_clk),
    .D(_01546_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_or[1] ));
 sky130_fd_sc_hd__dfxtp_1 _14932_ (.CLK(clknet_leaf_48_clk),
    .D(_01547_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_or[2] ));
 sky130_fd_sc_hd__dfxtp_1 _14933_ (.CLK(clknet_leaf_50_clk),
    .D(_01548_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_or[3] ));
 sky130_fd_sc_hd__dfxtp_1 _14934_ (.CLK(clknet_leaf_47_clk),
    .D(_01549_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_or[4] ));
 sky130_fd_sc_hd__dfxtp_1 _14935_ (.CLK(clknet_leaf_47_clk),
    .D(_01550_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_or[5] ));
 sky130_fd_sc_hd__dfxtp_1 _14936_ (.CLK(clknet_leaf_54_clk),
    .D(_01551_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_or[6] ));
 sky130_fd_sc_hd__dfxtp_1 _14937_ (.CLK(clknet_leaf_44_clk),
    .D(_01552_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_or[7] ));
 sky130_fd_sc_hd__dfxtp_1 _14938_ (.CLK(clknet_leaf_61_clk),
    .D(_01553_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_or[8] ));
 sky130_fd_sc_hd__dfxtp_1 _14939_ (.CLK(clknet_leaf_62_clk),
    .D(_01554_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_or[9] ));
 sky130_fd_sc_hd__dfxtp_1 _14940_ (.CLK(clknet_leaf_61_clk),
    .D(_01555_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_or[10] ));
 sky130_fd_sc_hd__dfxtp_1 _14941_ (.CLK(clknet_leaf_62_clk),
    .D(_01556_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_or[11] ));
 sky130_fd_sc_hd__dfxtp_1 _14942_ (.CLK(clknet_leaf_61_clk),
    .D(_01557_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_or[12] ));
 sky130_fd_sc_hd__dfxtp_1 _14943_ (.CLK(clknet_leaf_62_clk),
    .D(_01558_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_or[13] ));
 sky130_fd_sc_hd__dfxtp_1 _14944_ (.CLK(clknet_leaf_60_clk),
    .D(_01559_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_or[14] ));
 sky130_fd_sc_hd__dfxtp_1 _14945_ (.CLK(clknet_leaf_64_clk),
    .D(_01560_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_or[15] ));
 sky130_fd_sc_hd__dfxtp_1 _14946_ (.CLK(clknet_leaf_64_clk),
    .D(_01561_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_or[16] ));
 sky130_fd_sc_hd__dfxtp_1 _14947_ (.CLK(clknet_leaf_64_clk),
    .D(_01562_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_or[17] ));
 sky130_fd_sc_hd__dfxtp_1 _14948_ (.CLK(clknet_leaf_65_clk),
    .D(_01563_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_or[18] ));
 sky130_fd_sc_hd__dfxtp_1 _14949_ (.CLK(clknet_leaf_66_clk),
    .D(_01564_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_or[19] ));
 sky130_fd_sc_hd__dfxtp_1 _14950_ (.CLK(clknet_leaf_56_clk),
    .D(_01565_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_or[20] ));
 sky130_fd_sc_hd__dfxtp_1 _14951_ (.CLK(clknet_leaf_42_clk),
    .D(_01566_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_or[21] ));
 sky130_fd_sc_hd__dfxtp_1 _14952_ (.CLK(clknet_leaf_67_clk),
    .D(_01567_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_or[22] ));
 sky130_fd_sc_hd__dfxtp_1 _14953_ (.CLK(clknet_leaf_42_clk),
    .D(_01568_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_or[23] ));
 sky130_fd_sc_hd__dfxtp_1 _14954_ (.CLK(clknet_leaf_58_clk),
    .D(_01569_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_or[24] ));
 sky130_fd_sc_hd__dfxtp_1 _14955_ (.CLK(clknet_leaf_57_clk),
    .D(_01570_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_or[25] ));
 sky130_fd_sc_hd__dfxtp_1 _14956_ (.CLK(clknet_leaf_57_clk),
    .D(_01571_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_or[26] ));
 sky130_fd_sc_hd__dfxtp_1 _14957_ (.CLK(clknet_leaf_62_clk),
    .D(_01572_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_or[27] ));
 sky130_fd_sc_hd__dfxtp_1 _14958_ (.CLK(clknet_leaf_57_clk),
    .D(_01573_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_or[28] ));
 sky130_fd_sc_hd__dfxtp_1 _14959_ (.CLK(clknet_leaf_55_clk),
    .D(_01574_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_or[29] ));
 sky130_fd_sc_hd__dfxtp_1 _14960_ (.CLK(clknet_leaf_42_clk),
    .D(_01575_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_or[30] ));
 sky130_fd_sc_hd__dfxtp_1 _14961_ (.CLK(clknet_leaf_43_clk),
    .D(_01576_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_or[31] ));
 sky130_fd_sc_hd__dfxtp_1 _14962_ (.CLK(clknet_leaf_51_clk),
    .D(_01577_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_srl_sra[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14963_ (.CLK(clknet_leaf_51_clk),
    .D(_01578_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_srl_sra[1] ));
 sky130_fd_sc_hd__dfxtp_1 _14964_ (.CLK(clknet_leaf_51_clk),
    .D(_01579_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_srl_sra[2] ));
 sky130_fd_sc_hd__dfxtp_1 _14965_ (.CLK(clknet_leaf_54_clk),
    .D(_01580_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_srl_sra[3] ));
 sky130_fd_sc_hd__dfxtp_1 _14966_ (.CLK(clknet_leaf_51_clk),
    .D(_01581_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_srl_sra[4] ));
 sky130_fd_sc_hd__dfxtp_1 _14967_ (.CLK(clknet_leaf_54_clk),
    .D(_01582_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_srl_sra[5] ));
 sky130_fd_sc_hd__dfxtp_1 _14968_ (.CLK(clknet_leaf_54_clk),
    .D(_01583_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_srl_sra[6] ));
 sky130_fd_sc_hd__dfxtp_1 _14969_ (.CLK(clknet_leaf_43_clk),
    .D(_01584_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_srl_sra[7] ));
 sky130_fd_sc_hd__dfxtp_1 _14970_ (.CLK(clknet_leaf_58_clk),
    .D(_01585_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_srl_sra[8] ));
 sky130_fd_sc_hd__dfxtp_1 _14971_ (.CLK(clknet_leaf_58_clk),
    .D(_01586_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_srl_sra[9] ));
 sky130_fd_sc_hd__dfxtp_1 _14972_ (.CLK(clknet_leaf_58_clk),
    .D(_01587_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_srl_sra[10] ));
 sky130_fd_sc_hd__dfxtp_1 _14973_ (.CLK(clknet_leaf_57_clk),
    .D(_01588_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_srl_sra[11] ));
 sky130_fd_sc_hd__dfxtp_1 _14974_ (.CLK(clknet_leaf_58_clk),
    .D(_01589_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_srl_sra[12] ));
 sky130_fd_sc_hd__dfxtp_1 _14975_ (.CLK(clknet_leaf_65_clk),
    .D(_01590_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_srl_sra[13] ));
 sky130_fd_sc_hd__dfxtp_1 _14976_ (.CLK(clknet_leaf_60_clk),
    .D(_01591_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_srl_sra[14] ));
 sky130_fd_sc_hd__dfxtp_1 _14977_ (.CLK(clknet_leaf_65_clk),
    .D(_01592_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_srl_sra[15] ));
 sky130_fd_sc_hd__dfxtp_1 _14978_ (.CLK(clknet_leaf_60_clk),
    .D(_01593_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_srl_sra[16] ));
 sky130_fd_sc_hd__dfxtp_1 _14979_ (.CLK(clknet_leaf_58_clk),
    .D(_01594_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_srl_sra[17] ));
 sky130_fd_sc_hd__dfxtp_1 _14980_ (.CLK(clknet_leaf_58_clk),
    .D(_01595_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_srl_sra[18] ));
 sky130_fd_sc_hd__dfxtp_1 _14981_ (.CLK(clknet_leaf_42_clk),
    .D(_01596_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_srl_sra[19] ));
 sky130_fd_sc_hd__dfxtp_1 _14982_ (.CLK(clknet_leaf_56_clk),
    .D(_01597_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_srl_sra[20] ));
 sky130_fd_sc_hd__dfxtp_1 _14983_ (.CLK(clknet_leaf_55_clk),
    .D(_01598_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_srl_sra[21] ));
 sky130_fd_sc_hd__dfxtp_1 _14984_ (.CLK(clknet_leaf_55_clk),
    .D(_01599_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_srl_sra[22] ));
 sky130_fd_sc_hd__dfxtp_1 _14985_ (.CLK(clknet_leaf_55_clk),
    .D(_01600_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_srl_sra[23] ));
 sky130_fd_sc_hd__dfxtp_1 _14986_ (.CLK(clknet_leaf_58_clk),
    .D(_01601_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_srl_sra[24] ));
 sky130_fd_sc_hd__dfxtp_1 _14987_ (.CLK(clknet_leaf_58_clk),
    .D(_01602_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_srl_sra[25] ));
 sky130_fd_sc_hd__dfxtp_1 _14988_ (.CLK(clknet_leaf_58_clk),
    .D(_01603_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_srl_sra[26] ));
 sky130_fd_sc_hd__dfxtp_1 _14989_ (.CLK(clknet_leaf_57_clk),
    .D(_01604_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_srl_sra[27] ));
 sky130_fd_sc_hd__dfxtp_1 _14990_ (.CLK(clknet_leaf_57_clk),
    .D(_01605_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_srl_sra[28] ));
 sky130_fd_sc_hd__dfxtp_1 _14991_ (.CLK(clknet_leaf_55_clk),
    .D(_01606_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_srl_sra[29] ));
 sky130_fd_sc_hd__dfxtp_1 _14992_ (.CLK(clknet_leaf_55_clk),
    .D(_01607_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_srl_sra[30] ));
 sky130_fd_sc_hd__dfxtp_1 _14993_ (.CLK(clknet_leaf_43_clk),
    .D(_01608_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_srl_sra[31] ));
 sky130_fd_sc_hd__dfxtp_1 _14994_ (.CLK(clknet_leaf_45_clk),
    .D(_01609_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_xor[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14995_ (.CLK(clknet_leaf_48_clk),
    .D(_01610_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_xor[1] ));
 sky130_fd_sc_hd__dfxtp_1 _14996_ (.CLK(clknet_leaf_47_clk),
    .D(_01611_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_xor[2] ));
 sky130_fd_sc_hd__dfxtp_1 _14997_ (.CLK(clknet_leaf_50_clk),
    .D(_01612_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_xor[3] ));
 sky130_fd_sc_hd__dfxtp_1 _14998_ (.CLK(clknet_leaf_48_clk),
    .D(_01613_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_xor[4] ));
 sky130_fd_sc_hd__dfxtp_1 _14999_ (.CLK(clknet_leaf_47_clk),
    .D(_01614_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_xor[5] ));
 sky130_fd_sc_hd__dfxtp_1 _15000_ (.CLK(clknet_leaf_54_clk),
    .D(_01615_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_xor[6] ));
 sky130_fd_sc_hd__dfxtp_1 _15001_ (.CLK(clknet_leaf_43_clk),
    .D(_01616_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_xor[7] ));
 sky130_fd_sc_hd__dfxtp_1 _15002_ (.CLK(clknet_leaf_61_clk),
    .D(_01617_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_xor[8] ));
 sky130_fd_sc_hd__dfxtp_1 _15003_ (.CLK(clknet_leaf_61_clk),
    .D(_01618_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_xor[9] ));
 sky130_fd_sc_hd__dfxtp_1 _15004_ (.CLK(clknet_leaf_61_clk),
    .D(_01619_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_xor[10] ));
 sky130_fd_sc_hd__dfxtp_1 _15005_ (.CLK(clknet_leaf_62_clk),
    .D(_01620_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_xor[11] ));
 sky130_fd_sc_hd__dfxtp_1 _15006_ (.CLK(clknet_leaf_61_clk),
    .D(_01621_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_xor[12] ));
 sky130_fd_sc_hd__dfxtp_1 _15007_ (.CLK(clknet_leaf_65_clk),
    .D(_01622_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_xor[13] ));
 sky130_fd_sc_hd__dfxtp_1 _15008_ (.CLK(clknet_leaf_60_clk),
    .D(_01623_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_xor[14] ));
 sky130_fd_sc_hd__dfxtp_1 _15009_ (.CLK(clknet_leaf_64_clk),
    .D(_01624_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_xor[15] ));
 sky130_fd_sc_hd__dfxtp_1 _15010_ (.CLK(clknet_leaf_65_clk),
    .D(_01625_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_xor[16] ));
 sky130_fd_sc_hd__dfxtp_1 _15011_ (.CLK(clknet_leaf_65_clk),
    .D(_01626_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_xor[17] ));
 sky130_fd_sc_hd__dfxtp_1 _15012_ (.CLK(clknet_leaf_65_clk),
    .D(_01627_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_xor[18] ));
 sky130_fd_sc_hd__dfxtp_1 _15013_ (.CLK(clknet_leaf_66_clk),
    .D(_01628_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_xor[19] ));
 sky130_fd_sc_hd__dfxtp_1 _15014_ (.CLK(clknet_leaf_66_clk),
    .D(_01629_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_xor[20] ));
 sky130_fd_sc_hd__dfxtp_1 _15015_ (.CLK(clknet_leaf_56_clk),
    .D(_01630_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_xor[21] ));
 sky130_fd_sc_hd__dfxtp_1 _15016_ (.CLK(clknet_leaf_56_clk),
    .D(_01631_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_xor[22] ));
 sky130_fd_sc_hd__dfxtp_1 _15017_ (.CLK(clknet_leaf_56_clk),
    .D(_01632_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_xor[23] ));
 sky130_fd_sc_hd__dfxtp_1 _15018_ (.CLK(clknet_leaf_60_clk),
    .D(_01633_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_xor[24] ));
 sky130_fd_sc_hd__dfxtp_1 _15019_ (.CLK(clknet_leaf_60_clk),
    .D(_01634_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_xor[25] ));
 sky130_fd_sc_hd__dfxtp_1 _15020_ (.CLK(clknet_leaf_60_clk),
    .D(_01635_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_xor[26] ));
 sky130_fd_sc_hd__dfxtp_1 _15021_ (.CLK(clknet_leaf_57_clk),
    .D(_01636_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_xor[27] ));
 sky130_fd_sc_hd__dfxtp_1 _15022_ (.CLK(clknet_leaf_59_clk),
    .D(_01637_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_xor[28] ));
 sky130_fd_sc_hd__dfxtp_1 _15023_ (.CLK(clknet_leaf_55_clk),
    .D(_01638_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_xor[29] ));
 sky130_fd_sc_hd__dfxtp_1 _15024_ (.CLK(clknet_leaf_42_clk),
    .D(_01639_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_xor[30] ));
 sky130_fd_sc_hd__dfxtp_1 _15025_ (.CLK(clknet_leaf_42_clk),
    .D(_01640_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_xor[31] ));
 sky130_fd_sc_hd__dfxtp_1 _15026_ (.CLK(clknet_leaf_43_clk),
    .D(_01641_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_slt[0] ));
 sky130_fd_sc_hd__dfxtp_1 _15027_ (.CLK(clknet_leaf_55_clk),
    .D(_01642_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_sll[16] ));
 sky130_fd_sc_hd__dfxtp_2 _15028_ (.CLK(clknet_leaf_59_clk),
    .D(_01643_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_sll[17] ));
 sky130_fd_sc_hd__dfxtp_2 _15029_ (.CLK(clknet_leaf_59_clk),
    .D(_01644_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_sll[18] ));
 sky130_fd_sc_hd__dfxtp_2 _15030_ (.CLK(clknet_leaf_52_clk),
    .D(_01645_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_sll[19] ));
 sky130_fd_sc_hd__dfxtp_2 _15031_ (.CLK(clknet_5_10_0_clk),
    .D(_01646_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_sll[20] ));
 sky130_fd_sc_hd__dfxtp_2 _15032_ (.CLK(clknet_leaf_52_clk),
    .D(_01647_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_sll[21] ));
 sky130_fd_sc_hd__dfxtp_1 _15033_ (.CLK(clknet_leaf_59_clk),
    .D(_01648_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_sll[22] ));
 sky130_fd_sc_hd__dfxtp_2 _15034_ (.CLK(clknet_leaf_52_clk),
    .D(_01649_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_sll[23] ));
 sky130_fd_sc_hd__dfxtp_1 _15035_ (.CLK(clknet_leaf_59_clk),
    .D(_01650_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_sll[24] ));
 sky130_fd_sc_hd__dfxtp_1 _15036_ (.CLK(clknet_leaf_59_clk),
    .D(_01651_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_sll[25] ));
 sky130_fd_sc_hd__dfxtp_1 _15037_ (.CLK(clknet_leaf_59_clk),
    .D(_01652_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_sll[26] ));
 sky130_fd_sc_hd__dfxtp_1 _15038_ (.CLK(clknet_leaf_59_clk),
    .D(_01653_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_sll[27] ));
 sky130_fd_sc_hd__dfxtp_1 _15039_ (.CLK(clknet_leaf_59_clk),
    .D(_01654_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_sll[28] ));
 sky130_fd_sc_hd__dfxtp_1 _15040_ (.CLK(clknet_leaf_52_clk),
    .D(_01655_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_sll[29] ));
 sky130_fd_sc_hd__dfxtp_2 _15041_ (.CLK(clknet_leaf_59_clk),
    .D(_01656_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_sll[30] ));
 sky130_fd_sc_hd__dfxtp_1 _15042_ (.CLK(clknet_leaf_52_clk),
    .D(_01657_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_sll[31] ));
 sky130_fd_sc_hd__dfxtp_4 _15043_ (.CLK(clknet_leaf_45_clk),
    .D(_01658_),
    .Q(\core_busio.mem_address[0] ));
 sky130_fd_sc_hd__dfxtp_1 _15044_ (.CLK(clknet_leaf_46_clk),
    .D(_01659_),
    .Q(\core_busio.mem_address[1] ));
 sky130_fd_sc_hd__dfxtp_4 _15045_ (.CLK(clknet_leaf_46_clk),
    .D(_01660_),
    .Q(\core_busio.mem_address[2] ));
 sky130_fd_sc_hd__dfxtp_4 _15046_ (.CLK(clknet_leaf_45_clk),
    .D(_01661_),
    .Q(\core_busio.mem_address[3] ));
 sky130_fd_sc_hd__dfxtp_4 _15047_ (.CLK(clknet_leaf_44_clk),
    .D(_01662_),
    .Q(\core_busio.mem_address[4] ));
 sky130_fd_sc_hd__dfxtp_4 _15048_ (.CLK(clknet_leaf_44_clk),
    .D(_01663_),
    .Q(\core_busio.mem_address[5] ));
 sky130_fd_sc_hd__dfxtp_4 _15049_ (.CLK(clknet_leaf_41_clk),
    .D(_01664_),
    .Q(\core_busio.mem_address[6] ));
 sky130_fd_sc_hd__dfxtp_4 _15050_ (.CLK(clknet_leaf_39_clk),
    .D(_01665_),
    .Q(\core_busio.mem_address[7] ));
 sky130_fd_sc_hd__dfxtp_4 _15051_ (.CLK(clknet_leaf_63_clk),
    .D(_01666_),
    .Q(\core_busio.mem_address[8] ));
 sky130_fd_sc_hd__dfxtp_4 _15052_ (.CLK(clknet_leaf_63_clk),
    .D(_01667_),
    .Q(\core_busio.mem_address[9] ));
 sky130_fd_sc_hd__dfxtp_4 _15053_ (.CLK(clknet_leaf_63_clk),
    .D(_01668_),
    .Q(\core_busio.mem_address[10] ));
 sky130_fd_sc_hd__dfxtp_4 _15054_ (.CLK(clknet_leaf_63_clk),
    .D(_01669_),
    .Q(\core_busio.mem_address[11] ));
 sky130_fd_sc_hd__dfxtp_2 _15055_ (.CLK(clknet_leaf_70_clk),
    .D(_01670_),
    .Q(\core_busio.mem_address[12] ));
 sky130_fd_sc_hd__dfxtp_4 _15056_ (.CLK(clknet_leaf_71_clk),
    .D(_01671_),
    .Q(\core_busio.mem_address[13] ));
 sky130_fd_sc_hd__dfxtp_4 _15057_ (.CLK(clknet_leaf_71_clk),
    .D(_01672_),
    .Q(\core_busio.mem_address[14] ));
 sky130_fd_sc_hd__dfxtp_4 _15058_ (.CLK(clknet_leaf_71_clk),
    .D(_01673_),
    .Q(\core_busio.mem_address[15] ));
 sky130_fd_sc_hd__dfxtp_2 _15059_ (.CLK(clknet_leaf_70_clk),
    .D(_01674_),
    .Q(\core_busio.mem_address[16] ));
 sky130_fd_sc_hd__dfxtp_4 _15060_ (.CLK(clknet_leaf_69_clk),
    .D(_01675_),
    .Q(\core_busio.mem_address[17] ));
 sky130_fd_sc_hd__dfxtp_4 _15061_ (.CLK(clknet_leaf_69_clk),
    .D(_01676_),
    .Q(\core_busio.mem_address[18] ));
 sky130_fd_sc_hd__dfxtp_4 _15062_ (.CLK(clknet_leaf_69_clk),
    .D(_01677_),
    .Q(\core_busio.mem_address[19] ));
 sky130_fd_sc_hd__dfxtp_4 _15063_ (.CLK(clknet_leaf_82_clk),
    .D(_01678_),
    .Q(\core_busio.mem_address[20] ));
 sky130_fd_sc_hd__dfxtp_4 _15064_ (.CLK(clknet_leaf_82_clk),
    .D(_01679_),
    .Q(\core_busio.mem_address[21] ));
 sky130_fd_sc_hd__dfxtp_4 _15065_ (.CLK(clknet_leaf_82_clk),
    .D(_01680_),
    .Q(\core_busio.mem_address[22] ));
 sky130_fd_sc_hd__dfxtp_2 _15066_ (.CLK(clknet_leaf_82_clk),
    .D(_01681_),
    .Q(\core_busio.mem_address[23] ));
 sky130_fd_sc_hd__dfxtp_4 _15067_ (.CLK(clknet_leaf_69_clk),
    .D(_01682_),
    .Q(\core_busio.mem_address[24] ));
 sky130_fd_sc_hd__dfxtp_2 _15068_ (.CLK(clknet_leaf_68_clk),
    .D(_01683_),
    .Q(\core_busio.mem_address[25] ));
 sky130_fd_sc_hd__dfxtp_4 _15069_ (.CLK(clknet_leaf_68_clk),
    .D(_01684_),
    .Q(\core_busio.mem_address[26] ));
 sky130_fd_sc_hd__dfxtp_4 _15070_ (.CLK(clknet_leaf_67_clk),
    .D(_01685_),
    .Q(\core_busio.mem_address[27] ));
 sky130_fd_sc_hd__dfxtp_4 _15071_ (.CLK(clknet_leaf_83_clk),
    .D(_01686_),
    .Q(\core_busio.mem_address[28] ));
 sky130_fd_sc_hd__dfxtp_4 _15072_ (.CLK(clknet_leaf_42_clk),
    .D(_01687_),
    .Q(\core_busio.mem_address[29] ));
 sky130_fd_sc_hd__dfxtp_4 _15073_ (.CLK(clknet_leaf_41_clk),
    .D(_01688_),
    .Q(\core_busio.mem_address[30] ));
 sky130_fd_sc_hd__dfxtp_4 _15074_ (.CLK(clknet_leaf_41_clk),
    .D(_01689_),
    .Q(\core_busio.mem_address[31] ));
 sky130_fd_sc_hd__dfxtp_1 _15075_ (.CLK(clknet_leaf_152_clk),
    .D(_01690_),
    .Q(\core_pipeline.execute_to_memory_wfi ));
 sky130_fd_sc_hd__dfxtp_1 _15076_ (.CLK(clknet_leaf_251_clk),
    .D(_01691_),
    .Q(\core_pipeline.pipeline_registers.registers[17][0] ));
 sky130_fd_sc_hd__dfxtp_1 _15077_ (.CLK(clknet_leaf_164_clk),
    .D(_01692_),
    .Q(\core_pipeline.pipeline_registers.registers[17][1] ));
 sky130_fd_sc_hd__dfxtp_1 _15078_ (.CLK(clknet_leaf_197_clk),
    .D(_01693_),
    .Q(\core_pipeline.pipeline_registers.registers[17][2] ));
 sky130_fd_sc_hd__dfxtp_1 _15079_ (.CLK(clknet_leaf_235_clk),
    .D(_01694_),
    .Q(\core_pipeline.pipeline_registers.registers[17][3] ));
 sky130_fd_sc_hd__dfxtp_1 _15080_ (.CLK(clknet_leaf_250_clk),
    .D(_01695_),
    .Q(\core_pipeline.pipeline_registers.registers[17][4] ));
 sky130_fd_sc_hd__dfxtp_1 _15081_ (.CLK(clknet_leaf_202_clk),
    .D(_01696_),
    .Q(\core_pipeline.pipeline_registers.registers[17][5] ));
 sky130_fd_sc_hd__dfxtp_1 _15082_ (.CLK(clknet_leaf_207_clk),
    .D(_01697_),
    .Q(\core_pipeline.pipeline_registers.registers[17][6] ));
 sky130_fd_sc_hd__dfxtp_1 _15083_ (.CLK(clknet_leaf_232_clk),
    .D(_01698_),
    .Q(\core_pipeline.pipeline_registers.registers[17][7] ));
 sky130_fd_sc_hd__dfxtp_1 _15084_ (.CLK(clknet_leaf_238_clk),
    .D(_01699_),
    .Q(\core_pipeline.pipeline_registers.registers[17][8] ));
 sky130_fd_sc_hd__dfxtp_1 _15085_ (.CLK(clknet_leaf_6_clk),
    .D(_01700_),
    .Q(\core_pipeline.pipeline_registers.registers[17][9] ));
 sky130_fd_sc_hd__dfxtp_1 _15086_ (.CLK(clknet_leaf_8_clk),
    .D(_01701_),
    .Q(\core_pipeline.pipeline_registers.registers[17][10] ));
 sky130_fd_sc_hd__dfxtp_1 _15087_ (.CLK(clknet_leaf_5_clk),
    .D(_01702_),
    .Q(\core_pipeline.pipeline_registers.registers[17][11] ));
 sky130_fd_sc_hd__dfxtp_1 _15088_ (.CLK(clknet_leaf_25_clk),
    .D(_01703_),
    .Q(\core_pipeline.pipeline_registers.registers[17][12] ));
 sky130_fd_sc_hd__dfxtp_1 _15089_ (.CLK(clknet_leaf_22_clk),
    .D(_01704_),
    .Q(\core_pipeline.pipeline_registers.registers[17][13] ));
 sky130_fd_sc_hd__dfxtp_1 _15090_ (.CLK(clknet_leaf_6_clk),
    .D(_01705_),
    .Q(\core_pipeline.pipeline_registers.registers[17][14] ));
 sky130_fd_sc_hd__dfxtp_1 _15091_ (.CLK(clknet_leaf_20_clk),
    .D(_01706_),
    .Q(\core_pipeline.pipeline_registers.registers[17][15] ));
 sky130_fd_sc_hd__dfxtp_1 _15092_ (.CLK(clknet_leaf_245_clk),
    .D(_01707_),
    .Q(\core_pipeline.pipeline_registers.registers[17][16] ));
 sky130_fd_sc_hd__dfxtp_1 _15093_ (.CLK(clknet_leaf_213_clk),
    .D(_01708_),
    .Q(\core_pipeline.pipeline_registers.registers[17][17] ));
 sky130_fd_sc_hd__dfxtp_1 _15094_ (.CLK(clknet_leaf_181_clk),
    .D(_01709_),
    .Q(\core_pipeline.pipeline_registers.registers[17][18] ));
 sky130_fd_sc_hd__dfxtp_1 _15095_ (.CLK(clknet_leaf_195_clk),
    .D(_01710_),
    .Q(\core_pipeline.pipeline_registers.registers[17][19] ));
 sky130_fd_sc_hd__dfxtp_1 _15096_ (.CLK(clknet_leaf_190_clk),
    .D(_01711_),
    .Q(\core_pipeline.pipeline_registers.registers[17][20] ));
 sky130_fd_sc_hd__dfxtp_1 _15097_ (.CLK(clknet_leaf_170_clk),
    .D(_01712_),
    .Q(\core_pipeline.pipeline_registers.registers[17][21] ));
 sky130_fd_sc_hd__dfxtp_1 _15098_ (.CLK(clknet_leaf_211_clk),
    .D(_01713_),
    .Q(\core_pipeline.pipeline_registers.registers[17][22] ));
 sky130_fd_sc_hd__dfxtp_1 _15099_ (.CLK(clknet_leaf_217_clk),
    .D(_01714_),
    .Q(\core_pipeline.pipeline_registers.registers[17][23] ));
 sky130_fd_sc_hd__dfxtp_1 _15100_ (.CLK(clknet_leaf_225_clk),
    .D(_01715_),
    .Q(\core_pipeline.pipeline_registers.registers[17][24] ));
 sky130_fd_sc_hd__dfxtp_1 _15101_ (.CLK(clknet_leaf_8_clk),
    .D(_01716_),
    .Q(\core_pipeline.pipeline_registers.registers[17][25] ));
 sky130_fd_sc_hd__dfxtp_1 _15102_ (.CLK(clknet_leaf_18_clk),
    .D(_01717_),
    .Q(\core_pipeline.pipeline_registers.registers[17][26] ));
 sky130_fd_sc_hd__dfxtp_1 _15103_ (.CLK(clknet_leaf_168_clk),
    .D(_01718_),
    .Q(\core_pipeline.pipeline_registers.registers[17][27] ));
 sky130_fd_sc_hd__dfxtp_1 _15104_ (.CLK(clknet_leaf_183_clk),
    .D(_01719_),
    .Q(\core_pipeline.pipeline_registers.registers[17][28] ));
 sky130_fd_sc_hd__dfxtp_1 _15105_ (.CLK(clknet_leaf_212_clk),
    .D(_01720_),
    .Q(\core_pipeline.pipeline_registers.registers[17][29] ));
 sky130_fd_sc_hd__dfxtp_1 _15106_ (.CLK(clknet_leaf_210_clk),
    .D(_01721_),
    .Q(\core_pipeline.pipeline_registers.registers[17][30] ));
 sky130_fd_sc_hd__dfxtp_1 _15107_ (.CLK(clknet_leaf_177_clk),
    .D(_01722_),
    .Q(\core_pipeline.pipeline_registers.registers[17][31] ));
 sky130_fd_sc_hd__dfxtp_1 _15108_ (.CLK(clknet_leaf_251_clk),
    .D(_01723_),
    .Q(\core_pipeline.pipeline_registers.registers[16][0] ));
 sky130_fd_sc_hd__dfxtp_1 _15109_ (.CLK(clknet_leaf_161_clk),
    .D(_01724_),
    .Q(\core_pipeline.pipeline_registers.registers[16][1] ));
 sky130_fd_sc_hd__dfxtp_1 _15110_ (.CLK(clknet_leaf_197_clk),
    .D(_01725_),
    .Q(\core_pipeline.pipeline_registers.registers[16][2] ));
 sky130_fd_sc_hd__dfxtp_1 _15111_ (.CLK(clknet_leaf_236_clk),
    .D(_01726_),
    .Q(\core_pipeline.pipeline_registers.registers[16][3] ));
 sky130_fd_sc_hd__dfxtp_1 _15112_ (.CLK(clknet_leaf_250_clk),
    .D(_01727_),
    .Q(\core_pipeline.pipeline_registers.registers[16][4] ));
 sky130_fd_sc_hd__dfxtp_1 _15113_ (.CLK(clknet_leaf_199_clk),
    .D(_01728_),
    .Q(\core_pipeline.pipeline_registers.registers[16][5] ));
 sky130_fd_sc_hd__dfxtp_1 _15114_ (.CLK(clknet_leaf_207_clk),
    .D(_01729_),
    .Q(\core_pipeline.pipeline_registers.registers[16][6] ));
 sky130_fd_sc_hd__dfxtp_1 _15115_ (.CLK(clknet_leaf_232_clk),
    .D(_01730_),
    .Q(\core_pipeline.pipeline_registers.registers[16][7] ));
 sky130_fd_sc_hd__dfxtp_1 _15116_ (.CLK(clknet_leaf_238_clk),
    .D(_01731_),
    .Q(\core_pipeline.pipeline_registers.registers[16][8] ));
 sky130_fd_sc_hd__dfxtp_1 _15117_ (.CLK(clknet_leaf_248_clk),
    .D(_01732_),
    .Q(\core_pipeline.pipeline_registers.registers[16][9] ));
 sky130_fd_sc_hd__dfxtp_1 _15118_ (.CLK(clknet_leaf_8_clk),
    .D(_01733_),
    .Q(\core_pipeline.pipeline_registers.registers[16][10] ));
 sky130_fd_sc_hd__dfxtp_1 _15119_ (.CLK(clknet_leaf_249_clk),
    .D(_01734_),
    .Q(\core_pipeline.pipeline_registers.registers[16][11] ));
 sky130_fd_sc_hd__dfxtp_1 _15120_ (.CLK(clknet_leaf_229_clk),
    .D(_01735_),
    .Q(\core_pipeline.pipeline_registers.registers[16][12] ));
 sky130_fd_sc_hd__dfxtp_1 _15121_ (.CLK(clknet_leaf_9_clk),
    .D(_01736_),
    .Q(\core_pipeline.pipeline_registers.registers[16][13] ));
 sky130_fd_sc_hd__dfxtp_1 _15122_ (.CLK(clknet_leaf_6_clk),
    .D(_01737_),
    .Q(\core_pipeline.pipeline_registers.registers[16][14] ));
 sky130_fd_sc_hd__dfxtp_1 _15123_ (.CLK(clknet_leaf_28_clk),
    .D(_01738_),
    .Q(\core_pipeline.pipeline_registers.registers[16][15] ));
 sky130_fd_sc_hd__dfxtp_1 _15124_ (.CLK(clknet_leaf_245_clk),
    .D(_01739_),
    .Q(\core_pipeline.pipeline_registers.registers[16][16] ));
 sky130_fd_sc_hd__dfxtp_1 _15125_ (.CLK(clknet_leaf_163_clk),
    .D(_01740_),
    .Q(\core_pipeline.pipeline_registers.registers[16][17] ));
 sky130_fd_sc_hd__dfxtp_1 _15126_ (.CLK(clknet_leaf_179_clk),
    .D(_01741_),
    .Q(\core_pipeline.pipeline_registers.registers[16][18] ));
 sky130_fd_sc_hd__dfxtp_1 _15127_ (.CLK(clknet_leaf_194_clk),
    .D(_01742_),
    .Q(\core_pipeline.pipeline_registers.registers[16][19] ));
 sky130_fd_sc_hd__dfxtp_1 _15128_ (.CLK(clknet_leaf_187_clk),
    .D(_01743_),
    .Q(\core_pipeline.pipeline_registers.registers[16][20] ));
 sky130_fd_sc_hd__dfxtp_1 _15129_ (.CLK(clknet_leaf_170_clk),
    .D(_01744_),
    .Q(\core_pipeline.pipeline_registers.registers[16][21] ));
 sky130_fd_sc_hd__dfxtp_1 _15130_ (.CLK(clknet_leaf_211_clk),
    .D(_01745_),
    .Q(\core_pipeline.pipeline_registers.registers[16][22] ));
 sky130_fd_sc_hd__dfxtp_1 _15131_ (.CLK(clknet_leaf_217_clk),
    .D(_01746_),
    .Q(\core_pipeline.pipeline_registers.registers[16][23] ));
 sky130_fd_sc_hd__dfxtp_1 _15132_ (.CLK(clknet_leaf_225_clk),
    .D(_01747_),
    .Q(\core_pipeline.pipeline_registers.registers[16][24] ));
 sky130_fd_sc_hd__dfxtp_1 _15133_ (.CLK(clknet_leaf_8_clk),
    .D(_01748_),
    .Q(\core_pipeline.pipeline_registers.registers[16][25] ));
 sky130_fd_sc_hd__dfxtp_1 _15134_ (.CLK(clknet_leaf_21_clk),
    .D(_01749_),
    .Q(\core_pipeline.pipeline_registers.registers[16][26] ));
 sky130_fd_sc_hd__dfxtp_1 _15135_ (.CLK(clknet_leaf_168_clk),
    .D(_01750_),
    .Q(\core_pipeline.pipeline_registers.registers[16][27] ));
 sky130_fd_sc_hd__dfxtp_1 _15136_ (.CLK(clknet_leaf_183_clk),
    .D(_01751_),
    .Q(\core_pipeline.pipeline_registers.registers[16][28] ));
 sky130_fd_sc_hd__dfxtp_1 _15137_ (.CLK(clknet_leaf_212_clk),
    .D(_01752_),
    .Q(\core_pipeline.pipeline_registers.registers[16][29] ));
 sky130_fd_sc_hd__dfxtp_1 _15138_ (.CLK(clknet_leaf_210_clk),
    .D(_01753_),
    .Q(\core_pipeline.pipeline_registers.registers[16][30] ));
 sky130_fd_sc_hd__dfxtp_1 _15139_ (.CLK(clknet_leaf_176_clk),
    .D(_01754_),
    .Q(\core_pipeline.pipeline_registers.registers[16][31] ));
 sky130_fd_sc_hd__dfxtp_1 _15140_ (.CLK(clknet_leaf_255_clk),
    .D(_01755_),
    .Q(\core_pipeline.pipeline_registers.registers[15][0] ));
 sky130_fd_sc_hd__dfxtp_1 _15141_ (.CLK(clknet_leaf_166_clk),
    .D(_01756_),
    .Q(\core_pipeline.pipeline_registers.registers[15][1] ));
 sky130_fd_sc_hd__dfxtp_1 _15142_ (.CLK(clknet_leaf_200_clk),
    .D(_01757_),
    .Q(\core_pipeline.pipeline_registers.registers[15][2] ));
 sky130_fd_sc_hd__dfxtp_1 _15143_ (.CLK(clknet_leaf_246_clk),
    .D(_01758_),
    .Q(\core_pipeline.pipeline_registers.registers[15][3] ));
 sky130_fd_sc_hd__dfxtp_1 _15144_ (.CLK(clknet_leaf_0_clk),
    .D(_01759_),
    .Q(\core_pipeline.pipeline_registers.registers[15][4] ));
 sky130_fd_sc_hd__dfxtp_1 _15145_ (.CLK(clknet_leaf_201_clk),
    .D(_01760_),
    .Q(\core_pipeline.pipeline_registers.registers[15][5] ));
 sky130_fd_sc_hd__dfxtp_1 _15146_ (.CLK(clknet_leaf_240_clk),
    .D(_01761_),
    .Q(\core_pipeline.pipeline_registers.registers[15][6] ));
 sky130_fd_sc_hd__dfxtp_1 _15147_ (.CLK(clknet_leaf_2_clk),
    .D(_01762_),
    .Q(\core_pipeline.pipeline_registers.registers[15][7] ));
 sky130_fd_sc_hd__dfxtp_1 _15148_ (.CLK(clknet_leaf_241_clk),
    .D(_01763_),
    .Q(\core_pipeline.pipeline_registers.registers[15][8] ));
 sky130_fd_sc_hd__dfxtp_1 _15149_ (.CLK(clknet_leaf_11_clk),
    .D(_01764_),
    .Q(\core_pipeline.pipeline_registers.registers[15][9] ));
 sky130_fd_sc_hd__dfxtp_1 _15150_ (.CLK(clknet_leaf_13_clk),
    .D(_01765_),
    .Q(\core_pipeline.pipeline_registers.registers[15][10] ));
 sky130_fd_sc_hd__dfxtp_1 _15151_ (.CLK(clknet_leaf_2_clk),
    .D(_01766_),
    .Q(\core_pipeline.pipeline_registers.registers[15][11] ));
 sky130_fd_sc_hd__dfxtp_1 _15152_ (.CLK(clknet_leaf_249_clk),
    .D(_01767_),
    .Q(\core_pipeline.pipeline_registers.registers[15][12] ));
 sky130_fd_sc_hd__dfxtp_1 _15153_ (.CLK(clknet_leaf_12_clk),
    .D(_01768_),
    .Q(\core_pipeline.pipeline_registers.registers[15][13] ));
 sky130_fd_sc_hd__dfxtp_1 _15154_ (.CLK(clknet_leaf_15_clk),
    .D(_01769_),
    .Q(\core_pipeline.pipeline_registers.registers[15][14] ));
 sky130_fd_sc_hd__dfxtp_1 _15155_ (.CLK(clknet_leaf_19_clk),
    .D(_01770_),
    .Q(\core_pipeline.pipeline_registers.registers[15][15] ));
 sky130_fd_sc_hd__dfxtp_1 _15156_ (.CLK(clknet_leaf_252_clk),
    .D(_01771_),
    .Q(\core_pipeline.pipeline_registers.registers[15][16] ));
 sky130_fd_sc_hd__dfxtp_1 _15157_ (.CLK(clknet_leaf_213_clk),
    .D(_01772_),
    .Q(\core_pipeline.pipeline_registers.registers[15][17] ));
 sky130_fd_sc_hd__dfxtp_1 _15158_ (.CLK(clknet_leaf_183_clk),
    .D(_01773_),
    .Q(\core_pipeline.pipeline_registers.registers[15][18] ));
 sky130_fd_sc_hd__dfxtp_1 _15159_ (.CLK(clknet_leaf_192_clk),
    .D(_01774_),
    .Q(\core_pipeline.pipeline_registers.registers[15][19] ));
 sky130_fd_sc_hd__dfxtp_1 _15160_ (.CLK(clknet_leaf_191_clk),
    .D(_01775_),
    .Q(\core_pipeline.pipeline_registers.registers[15][20] ));
 sky130_fd_sc_hd__dfxtp_1 _15161_ (.CLK(clknet_leaf_169_clk),
    .D(_01776_),
    .Q(\core_pipeline.pipeline_registers.registers[15][21] ));
 sky130_fd_sc_hd__dfxtp_1 _15162_ (.CLK(clknet_leaf_203_clk),
    .D(_01777_),
    .Q(\core_pipeline.pipeline_registers.registers[15][22] ));
 sky130_fd_sc_hd__dfxtp_1 _15163_ (.CLK(clknet_leaf_218_clk),
    .D(_01778_),
    .Q(\core_pipeline.pipeline_registers.registers[15][23] ));
 sky130_fd_sc_hd__dfxtp_1 _15164_ (.CLK(clknet_leaf_229_clk),
    .D(_01779_),
    .Q(\core_pipeline.pipeline_registers.registers[15][24] ));
 sky130_fd_sc_hd__dfxtp_1 _15165_ (.CLK(clknet_leaf_14_clk),
    .D(_01780_),
    .Q(\core_pipeline.pipeline_registers.registers[15][25] ));
 sky130_fd_sc_hd__dfxtp_1 _15166_ (.CLK(clknet_leaf_16_clk),
    .D(_01781_),
    .Q(\core_pipeline.pipeline_registers.registers[15][26] ));
 sky130_fd_sc_hd__dfxtp_1 _15167_ (.CLK(clknet_leaf_170_clk),
    .D(_01782_),
    .Q(\core_pipeline.pipeline_registers.registers[15][27] ));
 sky130_fd_sc_hd__dfxtp_1 _15168_ (.CLK(clknet_leaf_176_clk),
    .D(_01783_),
    .Q(\core_pipeline.pipeline_registers.registers[15][28] ));
 sky130_fd_sc_hd__dfxtp_1 _15169_ (.CLK(clknet_leaf_214_clk),
    .D(_01784_),
    .Q(\core_pipeline.pipeline_registers.registers[15][29] ));
 sky130_fd_sc_hd__dfxtp_1 _15170_ (.CLK(clknet_leaf_236_clk),
    .D(_01785_),
    .Q(\core_pipeline.pipeline_registers.registers[15][30] ));
 sky130_fd_sc_hd__dfxtp_1 _15171_ (.CLK(clknet_leaf_173_clk),
    .D(_01786_),
    .Q(\core_pipeline.pipeline_registers.registers[15][31] ));
 sky130_fd_sc_hd__dfxtp_1 _15172_ (.CLK(clknet_leaf_253_clk),
    .D(_01787_),
    .Q(\core_pipeline.pipeline_registers.registers[9][0] ));
 sky130_fd_sc_hd__dfxtp_1 _15173_ (.CLK(clknet_leaf_161_clk),
    .D(_01788_),
    .Q(\core_pipeline.pipeline_registers.registers[9][1] ));
 sky130_fd_sc_hd__dfxtp_1 _15174_ (.CLK(clknet_leaf_192_clk),
    .D(_01789_),
    .Q(\core_pipeline.pipeline_registers.registers[9][2] ));
 sky130_fd_sc_hd__dfxtp_1 _15175_ (.CLK(clknet_leaf_246_clk),
    .D(_01790_),
    .Q(\core_pipeline.pipeline_registers.registers[9][3] ));
 sky130_fd_sc_hd__dfxtp_1 _15176_ (.CLK(clknet_leaf_256_clk),
    .D(_01791_),
    .Q(\core_pipeline.pipeline_registers.registers[9][4] ));
 sky130_fd_sc_hd__dfxtp_1 _15177_ (.CLK(clknet_leaf_201_clk),
    .D(_01792_),
    .Q(\core_pipeline.pipeline_registers.registers[9][5] ));
 sky130_fd_sc_hd__dfxtp_1 _15178_ (.CLK(clknet_leaf_205_clk),
    .D(_01793_),
    .Q(\core_pipeline.pipeline_registers.registers[9][6] ));
 sky130_fd_sc_hd__dfxtp_1 _15179_ (.CLK(clknet_leaf_2_clk),
    .D(_01794_),
    .Q(\core_pipeline.pipeline_registers.registers[9][7] ));
 sky130_fd_sc_hd__dfxtp_1 _15180_ (.CLK(clknet_leaf_240_clk),
    .D(_01795_),
    .Q(\core_pipeline.pipeline_registers.registers[9][8] ));
 sky130_fd_sc_hd__dfxtp_1 _15181_ (.CLK(clknet_leaf_3_clk),
    .D(_01796_),
    .Q(\core_pipeline.pipeline_registers.registers[9][9] ));
 sky130_fd_sc_hd__dfxtp_1 _15182_ (.CLK(clknet_leaf_14_clk),
    .D(_01797_),
    .Q(\core_pipeline.pipeline_registers.registers[9][10] ));
 sky130_fd_sc_hd__dfxtp_1 _15183_ (.CLK(clknet_leaf_2_clk),
    .D(_01798_),
    .Q(\core_pipeline.pipeline_registers.registers[9][11] ));
 sky130_fd_sc_hd__dfxtp_1 _15184_ (.CLK(clknet_leaf_248_clk),
    .D(_01799_),
    .Q(\core_pipeline.pipeline_registers.registers[9][12] ));
 sky130_fd_sc_hd__dfxtp_1 _15185_ (.CLK(clknet_leaf_11_clk),
    .D(_01800_),
    .Q(\core_pipeline.pipeline_registers.registers[9][13] ));
 sky130_fd_sc_hd__dfxtp_1 _15186_ (.CLK(clknet_leaf_15_clk),
    .D(_01801_),
    .Q(\core_pipeline.pipeline_registers.registers[9][14] ));
 sky130_fd_sc_hd__dfxtp_1 _15187_ (.CLK(clknet_leaf_46_clk),
    .D(_01802_),
    .Q(\core_pipeline.pipeline_registers.registers[9][15] ));
 sky130_fd_sc_hd__dfxtp_1 _15188_ (.CLK(clknet_leaf_252_clk),
    .D(_01803_),
    .Q(\core_pipeline.pipeline_registers.registers[9][16] ));
 sky130_fd_sc_hd__dfxtp_1 _15189_ (.CLK(clknet_leaf_213_clk),
    .D(_01804_),
    .Q(\core_pipeline.pipeline_registers.registers[9][17] ));
 sky130_fd_sc_hd__dfxtp_1 _15190_ (.CLK(clknet_leaf_186_clk),
    .D(_01805_),
    .Q(\core_pipeline.pipeline_registers.registers[9][18] ));
 sky130_fd_sc_hd__dfxtp_1 _15191_ (.CLK(clknet_leaf_191_clk),
    .D(_01806_),
    .Q(\core_pipeline.pipeline_registers.registers[9][19] ));
 sky130_fd_sc_hd__dfxtp_1 _15192_ (.CLK(clknet_leaf_188_clk),
    .D(_01807_),
    .Q(\core_pipeline.pipeline_registers.registers[9][20] ));
 sky130_fd_sc_hd__dfxtp_1 _15193_ (.CLK(clknet_leaf_173_clk),
    .D(_01808_),
    .Q(\core_pipeline.pipeline_registers.registers[9][21] ));
 sky130_fd_sc_hd__dfxtp_1 _15194_ (.CLK(clknet_leaf_203_clk),
    .D(_01809_),
    .Q(\core_pipeline.pipeline_registers.registers[9][22] ));
 sky130_fd_sc_hd__dfxtp_1 _15195_ (.CLK(clknet_leaf_218_clk),
    .D(_01810_),
    .Q(\core_pipeline.pipeline_registers.registers[9][23] ));
 sky130_fd_sc_hd__dfxtp_1 _15196_ (.CLK(clknet_leaf_235_clk),
    .D(_01811_),
    .Q(\core_pipeline.pipeline_registers.registers[9][24] ));
 sky130_fd_sc_hd__dfxtp_1 _15197_ (.CLK(clknet_leaf_12_clk),
    .D(_01812_),
    .Q(\core_pipeline.pipeline_registers.registers[9][25] ));
 sky130_fd_sc_hd__dfxtp_1 _15198_ (.CLK(clknet_leaf_18_clk),
    .D(_01813_),
    .Q(\core_pipeline.pipeline_registers.registers[9][26] ));
 sky130_fd_sc_hd__dfxtp_1 _15199_ (.CLK(clknet_leaf_138_clk),
    .D(_01814_),
    .Q(\core_pipeline.pipeline_registers.registers[9][27] ));
 sky130_fd_sc_hd__dfxtp_1 _15200_ (.CLK(clknet_leaf_184_clk),
    .D(_01815_),
    .Q(\core_pipeline.pipeline_registers.registers[9][28] ));
 sky130_fd_sc_hd__dfxtp_1 _15201_ (.CLK(clknet_leaf_212_clk),
    .D(_01816_),
    .Q(\core_pipeline.pipeline_registers.registers[9][29] ));
 sky130_fd_sc_hd__dfxtp_1 _15202_ (.CLK(clknet_leaf_237_clk),
    .D(_01817_),
    .Q(\core_pipeline.pipeline_registers.registers[9][30] ));
 sky130_fd_sc_hd__dfxtp_1 _15203_ (.CLK(clknet_leaf_174_clk),
    .D(_01818_),
    .Q(\core_pipeline.pipeline_registers.registers[9][31] ));
 sky130_fd_sc_hd__dfxtp_1 _15204_ (.CLK(clknet_leaf_149_clk),
    .D(_01819_),
    .Q(\core_pipeline.memory_to_writeback_ecause[1] ));
 sky130_fd_sc_hd__dfxtp_1 _15205_ (.CLK(clknet_leaf_149_clk),
    .D(_01820_),
    .Q(\core_pipeline.memory_to_writeback_ecause[2] ));
 sky130_fd_sc_hd__dfxtp_1 _15206_ (.CLK(clknet_leaf_157_clk),
    .D(_01821_),
    .Q(\core_pipeline.execute_to_memory_ecause[0] ));
 sky130_fd_sc_hd__dfxtp_1 _15207_ (.CLK(clknet_leaf_150_clk),
    .D(_01822_),
    .Q(\core_pipeline.execute_to_memory_ecause[1] ));
 sky130_fd_sc_hd__dfxtp_1 _15208_ (.CLK(clknet_leaf_157_clk),
    .D(_01823_),
    .Q(\core_pipeline.execute_to_memory_ecause[3] ));
 sky130_fd_sc_hd__dfxtp_1 _15209_ (.CLK(clknet_leaf_255_clk),
    .D(_01824_),
    .Q(\core_pipeline.pipeline_registers.registers[14][0] ));
 sky130_fd_sc_hd__dfxtp_1 _15210_ (.CLK(clknet_leaf_166_clk),
    .D(_01825_),
    .Q(\core_pipeline.pipeline_registers.registers[14][1] ));
 sky130_fd_sc_hd__dfxtp_1 _15211_ (.CLK(clknet_leaf_199_clk),
    .D(_01826_),
    .Q(\core_pipeline.pipeline_registers.registers[14][2] ));
 sky130_fd_sc_hd__dfxtp_1 _15212_ (.CLK(clknet_leaf_246_clk),
    .D(_01827_),
    .Q(\core_pipeline.pipeline_registers.registers[14][3] ));
 sky130_fd_sc_hd__dfxtp_1 _15213_ (.CLK(clknet_leaf_0_clk),
    .D(_01828_),
    .Q(\core_pipeline.pipeline_registers.registers[14][4] ));
 sky130_fd_sc_hd__dfxtp_1 _15214_ (.CLK(clknet_leaf_201_clk),
    .D(_01829_),
    .Q(\core_pipeline.pipeline_registers.registers[14][5] ));
 sky130_fd_sc_hd__dfxtp_1 _15215_ (.CLK(clknet_leaf_240_clk),
    .D(_01830_),
    .Q(\core_pipeline.pipeline_registers.registers[14][6] ));
 sky130_fd_sc_hd__dfxtp_1 _15216_ (.CLK(clknet_leaf_2_clk),
    .D(_01831_),
    .Q(\core_pipeline.pipeline_registers.registers[14][7] ));
 sky130_fd_sc_hd__dfxtp_1 _15217_ (.CLK(clknet_leaf_241_clk),
    .D(_01832_),
    .Q(\core_pipeline.pipeline_registers.registers[14][8] ));
 sky130_fd_sc_hd__dfxtp_1 _15218_ (.CLK(clknet_leaf_11_clk),
    .D(_01833_),
    .Q(\core_pipeline.pipeline_registers.registers[14][9] ));
 sky130_fd_sc_hd__dfxtp_1 _15219_ (.CLK(clknet_leaf_13_clk),
    .D(_01834_),
    .Q(\core_pipeline.pipeline_registers.registers[14][10] ));
 sky130_fd_sc_hd__dfxtp_1 _15220_ (.CLK(clknet_leaf_2_clk),
    .D(_01835_),
    .Q(\core_pipeline.pipeline_registers.registers[14][11] ));
 sky130_fd_sc_hd__dfxtp_1 _15221_ (.CLK(clknet_leaf_249_clk),
    .D(_01836_),
    .Q(\core_pipeline.pipeline_registers.registers[14][12] ));
 sky130_fd_sc_hd__dfxtp_1 _15222_ (.CLK(clknet_leaf_12_clk),
    .D(_01837_),
    .Q(\core_pipeline.pipeline_registers.registers[14][13] ));
 sky130_fd_sc_hd__dfxtp_1 _15223_ (.CLK(clknet_leaf_15_clk),
    .D(_01838_),
    .Q(\core_pipeline.pipeline_registers.registers[14][14] ));
 sky130_fd_sc_hd__dfxtp_1 _15224_ (.CLK(clknet_leaf_19_clk),
    .D(_01839_),
    .Q(\core_pipeline.pipeline_registers.registers[14][15] ));
 sky130_fd_sc_hd__dfxtp_1 _15225_ (.CLK(clknet_leaf_252_clk),
    .D(_01840_),
    .Q(\core_pipeline.pipeline_registers.registers[14][16] ));
 sky130_fd_sc_hd__dfxtp_1 _15226_ (.CLK(clknet_leaf_212_clk),
    .D(_01841_),
    .Q(\core_pipeline.pipeline_registers.registers[14][17] ));
 sky130_fd_sc_hd__dfxtp_1 _15227_ (.CLK(clknet_leaf_183_clk),
    .D(_01842_),
    .Q(\core_pipeline.pipeline_registers.registers[14][18] ));
 sky130_fd_sc_hd__dfxtp_1 _15228_ (.CLK(clknet_leaf_192_clk),
    .D(_01843_),
    .Q(\core_pipeline.pipeline_registers.registers[14][19] ));
 sky130_fd_sc_hd__dfxtp_1 _15229_ (.CLK(clknet_leaf_191_clk),
    .D(_01844_),
    .Q(\core_pipeline.pipeline_registers.registers[14][20] ));
 sky130_fd_sc_hd__dfxtp_1 _15230_ (.CLK(clknet_leaf_170_clk),
    .D(_01845_),
    .Q(\core_pipeline.pipeline_registers.registers[14][21] ));
 sky130_fd_sc_hd__dfxtp_1 _15231_ (.CLK(clknet_leaf_203_clk),
    .D(_01846_),
    .Q(\core_pipeline.pipeline_registers.registers[14][22] ));
 sky130_fd_sc_hd__dfxtp_1 _15232_ (.CLK(clknet_leaf_218_clk),
    .D(_01847_),
    .Q(\core_pipeline.pipeline_registers.registers[14][23] ));
 sky130_fd_sc_hd__dfxtp_1 _15233_ (.CLK(clknet_leaf_229_clk),
    .D(_01848_),
    .Q(\core_pipeline.pipeline_registers.registers[14][24] ));
 sky130_fd_sc_hd__dfxtp_1 _15234_ (.CLK(clknet_leaf_14_clk),
    .D(_01849_),
    .Q(\core_pipeline.pipeline_registers.registers[14][25] ));
 sky130_fd_sc_hd__dfxtp_1 _15235_ (.CLK(clknet_leaf_16_clk),
    .D(_01850_),
    .Q(\core_pipeline.pipeline_registers.registers[14][26] ));
 sky130_fd_sc_hd__dfxtp_1 _15236_ (.CLK(clknet_leaf_170_clk),
    .D(_01851_),
    .Q(\core_pipeline.pipeline_registers.registers[14][27] ));
 sky130_fd_sc_hd__dfxtp_1 _15237_ (.CLK(clknet_leaf_176_clk),
    .D(_01852_),
    .Q(\core_pipeline.pipeline_registers.registers[14][28] ));
 sky130_fd_sc_hd__dfxtp_1 _15238_ (.CLK(clknet_leaf_214_clk),
    .D(_01853_),
    .Q(\core_pipeline.pipeline_registers.registers[14][29] ));
 sky130_fd_sc_hd__dfxtp_1 _15239_ (.CLK(clknet_leaf_236_clk),
    .D(_01854_),
    .Q(\core_pipeline.pipeline_registers.registers[14][30] ));
 sky130_fd_sc_hd__dfxtp_1 _15240_ (.CLK(clknet_leaf_173_clk),
    .D(_01855_),
    .Q(\core_pipeline.pipeline_registers.registers[14][31] ));
 sky130_fd_sc_hd__dfxtp_1 _15241_ (.CLK(clknet_leaf_254_clk),
    .D(_01856_),
    .Q(\core_pipeline.pipeline_registers.registers[13][0] ));
 sky130_fd_sc_hd__dfxtp_1 _15242_ (.CLK(clknet_leaf_166_clk),
    .D(_01857_),
    .Q(\core_pipeline.pipeline_registers.registers[13][1] ));
 sky130_fd_sc_hd__dfxtp_1 _15243_ (.CLK(clknet_leaf_192_clk),
    .D(_01858_),
    .Q(\core_pipeline.pipeline_registers.registers[13][2] ));
 sky130_fd_sc_hd__dfxtp_1 _15244_ (.CLK(clknet_leaf_238_clk),
    .D(_01859_),
    .Q(\core_pipeline.pipeline_registers.registers[13][3] ));
 sky130_fd_sc_hd__dfxtp_1 _15245_ (.CLK(clknet_leaf_0_clk),
    .D(_01860_),
    .Q(\core_pipeline.pipeline_registers.registers[13][4] ));
 sky130_fd_sc_hd__dfxtp_1 _15246_ (.CLK(clknet_leaf_201_clk),
    .D(_01861_),
    .Q(\core_pipeline.pipeline_registers.registers[13][5] ));
 sky130_fd_sc_hd__dfxtp_1 _15247_ (.CLK(clknet_leaf_240_clk),
    .D(_01862_),
    .Q(\core_pipeline.pipeline_registers.registers[13][6] ));
 sky130_fd_sc_hd__dfxtp_1 _15248_ (.CLK(clknet_leaf_1_clk),
    .D(_01863_),
    .Q(\core_pipeline.pipeline_registers.registers[13][7] ));
 sky130_fd_sc_hd__dfxtp_1 _15249_ (.CLK(clknet_leaf_241_clk),
    .D(_01864_),
    .Q(\core_pipeline.pipeline_registers.registers[13][8] ));
 sky130_fd_sc_hd__dfxtp_1 _15250_ (.CLK(clknet_leaf_10_clk),
    .D(_01865_),
    .Q(\core_pipeline.pipeline_registers.registers[13][9] ));
 sky130_fd_sc_hd__dfxtp_1 _15251_ (.CLK(clknet_leaf_14_clk),
    .D(_01866_),
    .Q(\core_pipeline.pipeline_registers.registers[13][10] ));
 sky130_fd_sc_hd__dfxtp_1 _15252_ (.CLK(clknet_leaf_1_clk),
    .D(_01867_),
    .Q(\core_pipeline.pipeline_registers.registers[13][11] ));
 sky130_fd_sc_hd__dfxtp_1 _15253_ (.CLK(clknet_leaf_249_clk),
    .D(_01868_),
    .Q(\core_pipeline.pipeline_registers.registers[13][12] ));
 sky130_fd_sc_hd__dfxtp_1 _15254_ (.CLK(clknet_leaf_12_clk),
    .D(_01869_),
    .Q(\core_pipeline.pipeline_registers.registers[13][13] ));
 sky130_fd_sc_hd__dfxtp_1 _15255_ (.CLK(clknet_leaf_15_clk),
    .D(_01870_),
    .Q(\core_pipeline.pipeline_registers.registers[13][14] ));
 sky130_fd_sc_hd__dfxtp_1 _15256_ (.CLK(clknet_leaf_19_clk),
    .D(_01871_),
    .Q(\core_pipeline.pipeline_registers.registers[13][15] ));
 sky130_fd_sc_hd__dfxtp_1 _15257_ (.CLK(clknet_leaf_252_clk),
    .D(_01872_),
    .Q(\core_pipeline.pipeline_registers.registers[13][16] ));
 sky130_fd_sc_hd__dfxtp_1 _15258_ (.CLK(clknet_leaf_213_clk),
    .D(_01873_),
    .Q(\core_pipeline.pipeline_registers.registers[13][17] ));
 sky130_fd_sc_hd__dfxtp_1 _15259_ (.CLK(clknet_leaf_183_clk),
    .D(_01874_),
    .Q(\core_pipeline.pipeline_registers.registers[13][18] ));
 sky130_fd_sc_hd__dfxtp_1 _15260_ (.CLK(clknet_leaf_192_clk),
    .D(_01875_),
    .Q(\core_pipeline.pipeline_registers.registers[13][19] ));
 sky130_fd_sc_hd__dfxtp_1 _15261_ (.CLK(clknet_leaf_189_clk),
    .D(_01876_),
    .Q(\core_pipeline.pipeline_registers.registers[13][20] ));
 sky130_fd_sc_hd__dfxtp_1 _15262_ (.CLK(clknet_leaf_170_clk),
    .D(_01877_),
    .Q(\core_pipeline.pipeline_registers.registers[13][21] ));
 sky130_fd_sc_hd__dfxtp_1 _15263_ (.CLK(clknet_leaf_203_clk),
    .D(_01878_),
    .Q(\core_pipeline.pipeline_registers.registers[13][22] ));
 sky130_fd_sc_hd__dfxtp_1 _15264_ (.CLK(clknet_leaf_218_clk),
    .D(_01879_),
    .Q(\core_pipeline.pipeline_registers.registers[13][23] ));
 sky130_fd_sc_hd__dfxtp_1 _15265_ (.CLK(clknet_leaf_227_clk),
    .D(_01880_),
    .Q(\core_pipeline.pipeline_registers.registers[13][24] ));
 sky130_fd_sc_hd__dfxtp_1 _15266_ (.CLK(clknet_leaf_14_clk),
    .D(_01881_),
    .Q(\core_pipeline.pipeline_registers.registers[13][25] ));
 sky130_fd_sc_hd__dfxtp_1 _15267_ (.CLK(clknet_leaf_17_clk),
    .D(_01882_),
    .Q(\core_pipeline.pipeline_registers.registers[13][26] ));
 sky130_fd_sc_hd__dfxtp_1 _15268_ (.CLK(clknet_leaf_170_clk),
    .D(_01883_),
    .Q(\core_pipeline.pipeline_registers.registers[13][27] ));
 sky130_fd_sc_hd__dfxtp_1 _15269_ (.CLK(clknet_leaf_175_clk),
    .D(_01884_),
    .Q(\core_pipeline.pipeline_registers.registers[13][28] ));
 sky130_fd_sc_hd__dfxtp_1 _15270_ (.CLK(clknet_leaf_214_clk),
    .D(_01885_),
    .Q(\core_pipeline.pipeline_registers.registers[13][29] ));
 sky130_fd_sc_hd__dfxtp_1 _15271_ (.CLK(clknet_leaf_236_clk),
    .D(_01886_),
    .Q(\core_pipeline.pipeline_registers.registers[13][30] ));
 sky130_fd_sc_hd__dfxtp_1 _15272_ (.CLK(clknet_leaf_173_clk),
    .D(_01887_),
    .Q(\core_pipeline.pipeline_registers.registers[13][31] ));
 sky130_fd_sc_hd__dfxtp_1 _15273_ (.CLK(clknet_leaf_254_clk),
    .D(_01888_),
    .Q(\core_pipeline.pipeline_registers.registers[12][0] ));
 sky130_fd_sc_hd__dfxtp_1 _15274_ (.CLK(clknet_leaf_166_clk),
    .D(_01889_),
    .Q(\core_pipeline.pipeline_registers.registers[12][1] ));
 sky130_fd_sc_hd__dfxtp_1 _15275_ (.CLK(clknet_leaf_192_clk),
    .D(_01890_),
    .Q(\core_pipeline.pipeline_registers.registers[12][2] ));
 sky130_fd_sc_hd__dfxtp_1 _15276_ (.CLK(clknet_leaf_234_clk),
    .D(_01891_),
    .Q(\core_pipeline.pipeline_registers.registers[12][3] ));
 sky130_fd_sc_hd__dfxtp_1 _15277_ (.CLK(clknet_leaf_0_clk),
    .D(_01892_),
    .Q(\core_pipeline.pipeline_registers.registers[12][4] ));
 sky130_fd_sc_hd__dfxtp_1 _15278_ (.CLK(clknet_leaf_201_clk),
    .D(_01893_),
    .Q(\core_pipeline.pipeline_registers.registers[12][5] ));
 sky130_fd_sc_hd__dfxtp_1 _15279_ (.CLK(clknet_leaf_240_clk),
    .D(_01894_),
    .Q(\core_pipeline.pipeline_registers.registers[12][6] ));
 sky130_fd_sc_hd__dfxtp_1 _15280_ (.CLK(clknet_leaf_1_clk),
    .D(_01895_),
    .Q(\core_pipeline.pipeline_registers.registers[12][7] ));
 sky130_fd_sc_hd__dfxtp_1 _15281_ (.CLK(clknet_leaf_241_clk),
    .D(_01896_),
    .Q(\core_pipeline.pipeline_registers.registers[12][8] ));
 sky130_fd_sc_hd__dfxtp_1 _15282_ (.CLK(clknet_leaf_10_clk),
    .D(_01897_),
    .Q(\core_pipeline.pipeline_registers.registers[12][9] ));
 sky130_fd_sc_hd__dfxtp_1 _15283_ (.CLK(clknet_leaf_13_clk),
    .D(_01898_),
    .Q(\core_pipeline.pipeline_registers.registers[12][10] ));
 sky130_fd_sc_hd__dfxtp_1 _15284_ (.CLK(clknet_leaf_1_clk),
    .D(_01899_),
    .Q(\core_pipeline.pipeline_registers.registers[12][11] ));
 sky130_fd_sc_hd__dfxtp_1 _15285_ (.CLK(clknet_leaf_247_clk),
    .D(_01900_),
    .Q(\core_pipeline.pipeline_registers.registers[12][12] ));
 sky130_fd_sc_hd__dfxtp_1 _15286_ (.CLK(clknet_leaf_12_clk),
    .D(_01901_),
    .Q(\core_pipeline.pipeline_registers.registers[12][13] ));
 sky130_fd_sc_hd__dfxtp_1 _15287_ (.CLK(clknet_leaf_15_clk),
    .D(_01902_),
    .Q(\core_pipeline.pipeline_registers.registers[12][14] ));
 sky130_fd_sc_hd__dfxtp_1 _15288_ (.CLK(clknet_leaf_19_clk),
    .D(_01903_),
    .Q(\core_pipeline.pipeline_registers.registers[12][15] ));
 sky130_fd_sc_hd__dfxtp_1 _15289_ (.CLK(clknet_leaf_252_clk),
    .D(_01904_),
    .Q(\core_pipeline.pipeline_registers.registers[12][16] ));
 sky130_fd_sc_hd__dfxtp_1 _15290_ (.CLK(clknet_leaf_213_clk),
    .D(_01905_),
    .Q(\core_pipeline.pipeline_registers.registers[12][17] ));
 sky130_fd_sc_hd__dfxtp_1 _15291_ (.CLK(clknet_leaf_186_clk),
    .D(_01906_),
    .Q(\core_pipeline.pipeline_registers.registers[12][18] ));
 sky130_fd_sc_hd__dfxtp_1 _15292_ (.CLK(clknet_leaf_191_clk),
    .D(_01907_),
    .Q(\core_pipeline.pipeline_registers.registers[12][19] ));
 sky130_fd_sc_hd__dfxtp_1 _15293_ (.CLK(clknet_leaf_189_clk),
    .D(_01908_),
    .Q(\core_pipeline.pipeline_registers.registers[12][20] ));
 sky130_fd_sc_hd__dfxtp_1 _15294_ (.CLK(clknet_leaf_171_clk),
    .D(_01909_),
    .Q(\core_pipeline.pipeline_registers.registers[12][21] ));
 sky130_fd_sc_hd__dfxtp_1 _15295_ (.CLK(clknet_leaf_203_clk),
    .D(_01910_),
    .Q(\core_pipeline.pipeline_registers.registers[12][22] ));
 sky130_fd_sc_hd__dfxtp_1 _15296_ (.CLK(clknet_leaf_217_clk),
    .D(_01911_),
    .Q(\core_pipeline.pipeline_registers.registers[12][23] ));
 sky130_fd_sc_hd__dfxtp_1 _15297_ (.CLK(clknet_leaf_235_clk),
    .D(_01912_),
    .Q(\core_pipeline.pipeline_registers.registers[12][24] ));
 sky130_fd_sc_hd__dfxtp_1 _15298_ (.CLK(clknet_leaf_14_clk),
    .D(_01913_),
    .Q(\core_pipeline.pipeline_registers.registers[12][25] ));
 sky130_fd_sc_hd__dfxtp_1 _15299_ (.CLK(clknet_leaf_19_clk),
    .D(_01914_),
    .Q(\core_pipeline.pipeline_registers.registers[12][26] ));
 sky130_fd_sc_hd__dfxtp_1 _15300_ (.CLK(clknet_leaf_171_clk),
    .D(_01915_),
    .Q(\core_pipeline.pipeline_registers.registers[12][27] ));
 sky130_fd_sc_hd__dfxtp_1 _15301_ (.CLK(clknet_leaf_175_clk),
    .D(_01916_),
    .Q(\core_pipeline.pipeline_registers.registers[12][28] ));
 sky130_fd_sc_hd__dfxtp_1 _15302_ (.CLK(clknet_leaf_213_clk),
    .D(_01917_),
    .Q(\core_pipeline.pipeline_registers.registers[12][29] ));
 sky130_fd_sc_hd__dfxtp_1 _15303_ (.CLK(clknet_leaf_236_clk),
    .D(_01918_),
    .Q(\core_pipeline.pipeline_registers.registers[12][30] ));
 sky130_fd_sc_hd__dfxtp_1 _15304_ (.CLK(clknet_leaf_173_clk),
    .D(_01919_),
    .Q(\core_pipeline.pipeline_registers.registers[12][31] ));
 sky130_fd_sc_hd__dfxtp_1 _15305_ (.CLK(clknet_leaf_158_clk),
    .D(_01920_),
    .Q(\core_pipeline.memory_to_writeback_ecause[3] ));
 sky130_fd_sc_hd__dfxtp_1 _15306_ (.CLK(clknet_leaf_46_clk),
    .D(_01921_),
    .Q(\core_pipeline.decode_to_execute_rs1_data[0] ));
 sky130_fd_sc_hd__dfxtp_1 _15307_ (.CLK(clknet_leaf_223_clk),
    .D(_01922_),
    .Q(\core_pipeline.decode_to_execute_rs1_data[1] ));
 sky130_fd_sc_hd__dfxtp_1 _15308_ (.CLK(clknet_leaf_216_clk),
    .D(_01923_),
    .Q(\core_pipeline.decode_to_execute_rs1_data[2] ));
 sky130_fd_sc_hd__dfxtp_1 _15309_ (.CLK(clknet_leaf_228_clk),
    .D(_01924_),
    .Q(\core_pipeline.decode_to_execute_rs1_data[3] ));
 sky130_fd_sc_hd__dfxtp_1 _15310_ (.CLK(clknet_leaf_28_clk),
    .D(_01925_),
    .Q(\core_pipeline.decode_to_execute_rs1_data[4] ));
 sky130_fd_sc_hd__dfxtp_1 _15311_ (.CLK(clknet_leaf_220_clk),
    .D(_01926_),
    .Q(\core_pipeline.decode_to_execute_rs1_data[5] ));
 sky130_fd_sc_hd__dfxtp_1 _15312_ (.CLK(clknet_leaf_219_clk),
    .D(_01927_),
    .Q(\core_pipeline.decode_to_execute_rs1_data[6] ));
 sky130_fd_sc_hd__dfxtp_1 _15313_ (.CLK(clknet_leaf_228_clk),
    .D(_01928_),
    .Q(\core_pipeline.decode_to_execute_rs1_data[7] ));
 sky130_fd_sc_hd__dfxtp_2 _15314_ (.CLK(clknet_leaf_232_clk),
    .D(_01929_),
    .Q(\core_pipeline.decode_to_execute_rs1_data[8] ));
 sky130_fd_sc_hd__dfxtp_2 _15315_ (.CLK(clknet_leaf_21_clk),
    .D(_01930_),
    .Q(\core_pipeline.decode_to_execute_rs1_data[9] ));
 sky130_fd_sc_hd__dfxtp_1 _15316_ (.CLK(clknet_leaf_20_clk),
    .D(_01931_),
    .Q(\core_pipeline.decode_to_execute_rs1_data[10] ));
 sky130_fd_sc_hd__dfxtp_1 _15317_ (.CLK(clknet_leaf_26_clk),
    .D(_01932_),
    .Q(\core_pipeline.decode_to_execute_rs1_data[11] ));
 sky130_fd_sc_hd__dfxtp_1 _15318_ (.CLK(clknet_leaf_230_clk),
    .D(_01933_),
    .Q(\core_pipeline.decode_to_execute_rs1_data[12] ));
 sky130_fd_sc_hd__dfxtp_1 _15319_ (.CLK(clknet_leaf_19_clk),
    .D(_01934_),
    .Q(\core_pipeline.decode_to_execute_rs1_data[13] ));
 sky130_fd_sc_hd__dfxtp_1 _15320_ (.CLK(clknet_leaf_19_clk),
    .D(_01935_),
    .Q(\core_pipeline.decode_to_execute_rs1_data[14] ));
 sky130_fd_sc_hd__dfxtp_1 _15321_ (.CLK(clknet_leaf_20_clk),
    .D(_01936_),
    .Q(\core_pipeline.decode_to_execute_rs1_data[15] ));
 sky130_fd_sc_hd__dfxtp_1 _15322_ (.CLK(clknet_leaf_228_clk),
    .D(_01937_),
    .Q(\core_pipeline.decode_to_execute_rs1_data[16] ));
 sky130_fd_sc_hd__dfxtp_2 _15323_ (.CLK(clknet_leaf_213_clk),
    .D(_01938_),
    .Q(\core_pipeline.decode_to_execute_rs1_data[17] ));
 sky130_fd_sc_hd__dfxtp_2 _15324_ (.CLK(clknet_leaf_178_clk),
    .D(_01939_),
    .Q(\core_pipeline.decode_to_execute_rs1_data[18] ));
 sky130_fd_sc_hd__dfxtp_1 _15325_ (.CLK(clknet_leaf_166_clk),
    .D(_01940_),
    .Q(\core_pipeline.decode_to_execute_rs1_data[19] ));
 sky130_fd_sc_hd__dfxtp_4 _15326_ (.CLK(clknet_leaf_176_clk),
    .D(_01941_),
    .Q(\core_pipeline.decode_to_execute_rs1_data[20] ));
 sky130_fd_sc_hd__dfxtp_2 _15327_ (.CLK(clknet_leaf_168_clk),
    .D(_01942_),
    .Q(\core_pipeline.decode_to_execute_rs1_data[21] ));
 sky130_fd_sc_hd__dfxtp_1 _15328_ (.CLK(clknet_leaf_217_clk),
    .D(_01943_),
    .Q(\core_pipeline.decode_to_execute_rs1_data[22] ));
 sky130_fd_sc_hd__dfxtp_1 _15329_ (.CLK(clknet_leaf_219_clk),
    .D(_01944_),
    .Q(\core_pipeline.decode_to_execute_rs1_data[23] ));
 sky130_fd_sc_hd__dfxtp_1 _15330_ (.CLK(clknet_leaf_224_clk),
    .D(_01945_),
    .Q(\core_pipeline.decode_to_execute_rs1_data[24] ));
 sky130_fd_sc_hd__dfxtp_2 _15331_ (.CLK(clknet_leaf_22_clk),
    .D(_01946_),
    .Q(\core_pipeline.decode_to_execute_rs1_data[25] ));
 sky130_fd_sc_hd__dfxtp_1 _15332_ (.CLK(clknet_leaf_19_clk),
    .D(_01947_),
    .Q(\core_pipeline.decode_to_execute_rs1_data[26] ));
 sky130_fd_sc_hd__dfxtp_2 _15333_ (.CLK(clknet_leaf_168_clk),
    .D(_01948_),
    .Q(\core_pipeline.decode_to_execute_rs1_data[27] ));
 sky130_fd_sc_hd__dfxtp_2 _15334_ (.CLK(clknet_leaf_165_clk),
    .D(_01949_),
    .Q(\core_pipeline.decode_to_execute_rs1_data[28] ));
 sky130_fd_sc_hd__dfxtp_2 _15335_ (.CLK(clknet_leaf_214_clk),
    .D(_01950_),
    .Q(\core_pipeline.decode_to_execute_rs1_data[29] ));
 sky130_fd_sc_hd__dfxtp_1 _15336_ (.CLK(clknet_leaf_218_clk),
    .D(_01951_),
    .Q(\core_pipeline.decode_to_execute_rs1_data[30] ));
 sky130_fd_sc_hd__dfxtp_2 _15337_ (.CLK(clknet_leaf_166_clk),
    .D(_01952_),
    .Q(\core_pipeline.decode_to_execute_rs1_data[31] ));
 sky130_fd_sc_hd__dfxtp_4 _15338_ (.CLK(clknet_leaf_147_clk),
    .D(_01953_),
    .Q(\core_pipeline.pipeline_fetch.pc[2] ));
 sky130_fd_sc_hd__dfxtp_2 _15339_ (.CLK(clknet_leaf_151_clk),
    .D(_01954_),
    .Q(\core_pipeline.pipeline_fetch.pc[3] ));
 sky130_fd_sc_hd__dfxtp_2 _15340_ (.CLK(clknet_leaf_93_clk),
    .D(_01955_),
    .Q(\core_pipeline.pipeline_fetch.pc[4] ));
 sky130_fd_sc_hd__dfxtp_4 _15341_ (.CLK(clknet_leaf_147_clk),
    .D(_01956_),
    .Q(\core_pipeline.pipeline_fetch.pc[5] ));
 sky130_fd_sc_hd__dfxtp_4 _15342_ (.CLK(clknet_leaf_95_clk),
    .D(_01957_),
    .Q(\core_pipeline.pipeline_fetch.pc[6] ));
 sky130_fd_sc_hd__dfxtp_2 _15343_ (.CLK(clknet_leaf_98_clk),
    .D(_01958_),
    .Q(\core_pipeline.pipeline_fetch.pc[7] ));
 sky130_fd_sc_hd__dfxtp_2 _15344_ (.CLK(clknet_leaf_103_clk),
    .D(_01959_),
    .Q(\core_pipeline.pipeline_fetch.pc[8] ));
 sky130_fd_sc_hd__dfxtp_4 _15345_ (.CLK(clknet_leaf_107_clk),
    .D(_01960_),
    .Q(\core_pipeline.pipeline_fetch.pc[9] ));
 sky130_fd_sc_hd__dfxtp_2 _15346_ (.CLK(clknet_leaf_107_clk),
    .D(_01961_),
    .Q(\core_pipeline.pipeline_fetch.pc[10] ));
 sky130_fd_sc_hd__dfxtp_4 _15347_ (.CLK(clknet_leaf_108_clk),
    .D(_01962_),
    .Q(\core_pipeline.pipeline_fetch.pc[11] ));
 sky130_fd_sc_hd__dfxtp_4 _15348_ (.CLK(clknet_leaf_108_clk),
    .D(_01963_),
    .Q(\core_pipeline.pipeline_fetch.pc[12] ));
 sky130_fd_sc_hd__dfxtp_2 _15349_ (.CLK(clknet_leaf_109_clk),
    .D(_01964_),
    .Q(\core_pipeline.pipeline_fetch.pc[13] ));
 sky130_fd_sc_hd__dfxtp_2 _15350_ (.CLK(clknet_leaf_108_clk),
    .D(_01965_),
    .Q(\core_pipeline.pipeline_fetch.pc[14] ));
 sky130_fd_sc_hd__dfxtp_4 _15351_ (.CLK(clknet_leaf_108_clk),
    .D(_01966_),
    .Q(\core_pipeline.pipeline_fetch.pc[15] ));
 sky130_fd_sc_hd__dfxtp_2 _15352_ (.CLK(clknet_leaf_108_clk),
    .D(_01967_),
    .Q(\core_pipeline.pipeline_fetch.pc[16] ));
 sky130_fd_sc_hd__dfxtp_2 _15353_ (.CLK(clknet_leaf_109_clk),
    .D(_01968_),
    .Q(\core_pipeline.pipeline_fetch.pc[17] ));
 sky130_fd_sc_hd__dfxtp_2 _15354_ (.CLK(clknet_leaf_111_clk),
    .D(_01969_),
    .Q(\core_pipeline.pipeline_fetch.pc[18] ));
 sky130_fd_sc_hd__dfxtp_2 _15355_ (.CLK(clknet_leaf_110_clk),
    .D(_01970_),
    .Q(\core_pipeline.pipeline_fetch.pc[19] ));
 sky130_fd_sc_hd__dfxtp_2 _15356_ (.CLK(clknet_leaf_115_clk),
    .D(_01971_),
    .Q(\core_pipeline.pipeline_fetch.pc[20] ));
 sky130_fd_sc_hd__dfxtp_2 _15357_ (.CLK(clknet_leaf_116_clk),
    .D(_01972_),
    .Q(\core_pipeline.pipeline_fetch.pc[21] ));
 sky130_fd_sc_hd__dfxtp_2 _15358_ (.CLK(clknet_leaf_101_clk),
    .D(_01973_),
    .Q(\core_pipeline.pipeline_fetch.pc[22] ));
 sky130_fd_sc_hd__dfxtp_1 _15359_ (.CLK(clknet_leaf_105_clk),
    .D(_01974_),
    .Q(\core_pipeline.pipeline_fetch.pc[23] ));
 sky130_fd_sc_hd__dfxtp_4 _15360_ (.CLK(clknet_leaf_117_clk),
    .D(_01975_),
    .Q(\core_pipeline.pipeline_fetch.pc[24] ));
 sky130_fd_sc_hd__dfxtp_2 _15361_ (.CLK(clknet_leaf_105_clk),
    .D(_01976_),
    .Q(\core_pipeline.pipeline_fetch.pc[25] ));
 sky130_fd_sc_hd__dfxtp_2 _15362_ (.CLK(clknet_leaf_102_clk),
    .D(_01977_),
    .Q(\core_pipeline.pipeline_fetch.pc[26] ));
 sky130_fd_sc_hd__dfxtp_2 _15363_ (.CLK(clknet_leaf_102_clk),
    .D(_01978_),
    .Q(\core_pipeline.pipeline_fetch.pc[27] ));
 sky130_fd_sc_hd__dfxtp_2 _15364_ (.CLK(clknet_leaf_99_clk),
    .D(_01979_),
    .Q(\core_pipeline.pipeline_fetch.pc[28] ));
 sky130_fd_sc_hd__dfxtp_2 _15365_ (.CLK(clknet_leaf_96_clk),
    .D(_01980_),
    .Q(\core_pipeline.pipeline_fetch.pc[29] ));
 sky130_fd_sc_hd__dfxtp_4 _15366_ (.CLK(clknet_leaf_94_clk),
    .D(_01981_),
    .Q(\core_pipeline.pipeline_fetch.pc[30] ));
 sky130_fd_sc_hd__dfxtp_2 _15367_ (.CLK(clknet_leaf_146_clk),
    .D(_01982_),
    .Q(\core_pipeline.pipeline_fetch.pc[31] ));
 sky130_fd_sc_hd__dfxtp_1 _15368_ (.CLK(clknet_leaf_140_clk),
    .D(_01983_),
    .Q(\core_pipeline.pipeline_csr.mtimecmp[0] ));
 sky130_fd_sc_hd__dfxtp_1 _15369_ (.CLK(clknet_leaf_142_clk),
    .D(_01984_),
    .Q(\core_pipeline.pipeline_csr.mtimecmp[1] ));
 sky130_fd_sc_hd__dfxtp_1 _15370_ (.CLK(clknet_leaf_140_clk),
    .D(_01985_),
    .Q(\core_pipeline.pipeline_csr.mtimecmp[2] ));
 sky130_fd_sc_hd__dfxtp_1 _15371_ (.CLK(clknet_leaf_142_clk),
    .D(_01986_),
    .Q(\core_pipeline.pipeline_csr.mtimecmp[3] ));
 sky130_fd_sc_hd__dfxtp_1 _15372_ (.CLK(clknet_leaf_142_clk),
    .D(_01987_),
    .Q(\core_pipeline.pipeline_csr.mtimecmp[4] ));
 sky130_fd_sc_hd__dfxtp_1 _15373_ (.CLK(clknet_leaf_144_clk),
    .D(_01988_),
    .Q(\core_pipeline.pipeline_csr.mtimecmp[5] ));
 sky130_fd_sc_hd__dfxtp_1 _15374_ (.CLK(clknet_leaf_144_clk),
    .D(_01989_),
    .Q(\core_pipeline.pipeline_csr.mtimecmp[6] ));
 sky130_fd_sc_hd__dfxtp_2 _15375_ (.CLK(clknet_leaf_100_clk),
    .D(_01990_),
    .Q(\core_pipeline.pipeline_csr.mtimecmp[7] ));
 sky130_fd_sc_hd__dfxtp_1 _15376_ (.CLK(clknet_leaf_118_clk),
    .D(_01991_),
    .Q(\core_pipeline.pipeline_csr.mtimecmp[8] ));
 sky130_fd_sc_hd__dfxtp_1 _15377_ (.CLK(clknet_leaf_118_clk),
    .D(_01992_),
    .Q(\core_pipeline.pipeline_csr.mtimecmp[9] ));
 sky130_fd_sc_hd__dfxtp_1 _15378_ (.CLK(clknet_leaf_117_clk),
    .D(_01993_),
    .Q(\core_pipeline.pipeline_csr.mtimecmp[10] ));
 sky130_fd_sc_hd__dfxtp_2 _15379_ (.CLK(clknet_leaf_114_clk),
    .D(_01994_),
    .Q(\core_pipeline.pipeline_csr.mtimecmp[11] ));
 sky130_fd_sc_hd__dfxtp_1 _15380_ (.CLK(clknet_leaf_113_clk),
    .D(_01995_),
    .Q(\core_pipeline.pipeline_csr.mtimecmp[12] ));
 sky130_fd_sc_hd__dfxtp_1 _15381_ (.CLK(clknet_leaf_113_clk),
    .D(_01996_),
    .Q(\core_pipeline.pipeline_csr.mtimecmp[13] ));
 sky130_fd_sc_hd__dfxtp_1 _15382_ (.CLK(clknet_leaf_121_clk),
    .D(_01997_),
    .Q(\core_pipeline.pipeline_csr.mtimecmp[14] ));
 sky130_fd_sc_hd__dfxtp_1 _15383_ (.CLK(clknet_leaf_121_clk),
    .D(_01998_),
    .Q(\core_pipeline.pipeline_csr.mtimecmp[15] ));
 sky130_fd_sc_hd__dfxtp_1 _15384_ (.CLK(clknet_leaf_123_clk),
    .D(_01999_),
    .Q(\core_pipeline.pipeline_csr.mtimecmp[16] ));
 sky130_fd_sc_hd__dfxtp_1 _15385_ (.CLK(clknet_leaf_123_clk),
    .D(_02000_),
    .Q(\core_pipeline.pipeline_csr.mtimecmp[17] ));
 sky130_fd_sc_hd__dfxtp_1 _15386_ (.CLK(clknet_leaf_124_clk),
    .D(_02001_),
    .Q(\core_pipeline.pipeline_csr.mtimecmp[18] ));
 sky130_fd_sc_hd__dfxtp_1 _15387_ (.CLK(clknet_leaf_120_clk),
    .D(_02002_),
    .Q(\core_pipeline.pipeline_csr.mtimecmp[19] ));
 sky130_fd_sc_hd__dfxtp_1 _15388_ (.CLK(clknet_leaf_120_clk),
    .D(_02003_),
    .Q(\core_pipeline.pipeline_csr.mtimecmp[20] ));
 sky130_fd_sc_hd__dfxtp_1 _15389_ (.CLK(clknet_leaf_120_clk),
    .D(_02004_),
    .Q(\core_pipeline.pipeline_csr.mtimecmp[21] ));
 sky130_fd_sc_hd__dfxtp_1 _15390_ (.CLK(clknet_leaf_130_clk),
    .D(_02005_),
    .Q(\core_pipeline.pipeline_csr.mtimecmp[22] ));
 sky130_fd_sc_hd__dfxtp_1 _15391_ (.CLK(clknet_leaf_130_clk),
    .D(_02006_),
    .Q(\core_pipeline.pipeline_csr.mtimecmp[23] ));
 sky130_fd_sc_hd__dfxtp_1 _15392_ (.CLK(clknet_leaf_130_clk),
    .D(_02007_),
    .Q(\core_pipeline.pipeline_csr.mtimecmp[24] ));
 sky130_fd_sc_hd__dfxtp_1 _15393_ (.CLK(clknet_leaf_130_clk),
    .D(_02008_),
    .Q(\core_pipeline.pipeline_csr.mtimecmp[25] ));
 sky130_fd_sc_hd__dfxtp_1 _15394_ (.CLK(clknet_leaf_132_clk),
    .D(_02009_),
    .Q(\core_pipeline.pipeline_csr.mtimecmp[26] ));
 sky130_fd_sc_hd__dfxtp_1 _15395_ (.CLK(clknet_leaf_132_clk),
    .D(_02010_),
    .Q(\core_pipeline.pipeline_csr.mtimecmp[27] ));
 sky130_fd_sc_hd__dfxtp_1 _15396_ (.CLK(clknet_leaf_132_clk),
    .D(_02011_),
    .Q(\core_pipeline.pipeline_csr.mtimecmp[28] ));
 sky130_fd_sc_hd__dfxtp_2 _15397_ (.CLK(clknet_leaf_132_clk),
    .D(_02012_),
    .Q(\core_pipeline.pipeline_csr.mtimecmp[29] ));
 sky130_fd_sc_hd__dfxtp_2 _15398_ (.CLK(clknet_leaf_133_clk),
    .D(_02013_),
    .Q(\core_pipeline.pipeline_csr.mtimecmp[30] ));
 sky130_fd_sc_hd__dfxtp_2 _15399_ (.CLK(clknet_leaf_143_clk),
    .D(_02014_),
    .Q(\core_pipeline.pipeline_csr.mtimecmp[31] ));
 sky130_fd_sc_hd__dfxtp_2 _15400_ (.CLK(clknet_leaf_152_clk),
    .D(_02015_),
    .Q(\core_pipeline.decode_to_execute_pc[2] ));
 sky130_fd_sc_hd__dfxtp_2 _15401_ (.CLK(clknet_leaf_93_clk),
    .D(_02016_),
    .Q(\core_pipeline.decode_to_execute_pc[3] ));
 sky130_fd_sc_hd__dfxtp_1 _15402_ (.CLK(clknet_leaf_39_clk),
    .D(_02017_),
    .Q(\core_pipeline.decode_to_execute_pc[4] ));
 sky130_fd_sc_hd__dfxtp_1 _15403_ (.CLK(clknet_leaf_36_clk),
    .D(_02018_),
    .Q(\core_pipeline.decode_to_execute_pc[5] ));
 sky130_fd_sc_hd__dfxtp_1 _15404_ (.CLK(clknet_leaf_40_clk),
    .D(_02019_),
    .Q(\core_pipeline.decode_to_execute_pc[6] ));
 sky130_fd_sc_hd__dfxtp_2 _15405_ (.CLK(clknet_leaf_94_clk),
    .D(_02020_),
    .Q(\core_pipeline.decode_to_execute_pc[7] ));
 sky130_fd_sc_hd__dfxtp_2 _15406_ (.CLK(clknet_leaf_83_clk),
    .D(_02021_),
    .Q(\core_pipeline.decode_to_execute_pc[8] ));
 sky130_fd_sc_hd__dfxtp_2 _15407_ (.CLK(clknet_leaf_73_clk),
    .D(_02022_),
    .Q(\core_pipeline.decode_to_execute_pc[9] ));
 sky130_fd_sc_hd__dfxtp_2 _15408_ (.CLK(clknet_leaf_77_clk),
    .D(_02023_),
    .Q(\core_pipeline.decode_to_execute_pc[10] ));
 sky130_fd_sc_hd__dfxtp_2 _15409_ (.CLK(clknet_leaf_71_clk),
    .D(_02024_),
    .Q(\core_pipeline.decode_to_execute_pc[11] ));
 sky130_fd_sc_hd__dfxtp_2 _15410_ (.CLK(clknet_leaf_71_clk),
    .D(_02025_),
    .Q(\core_pipeline.decode_to_execute_pc[12] ));
 sky130_fd_sc_hd__dfxtp_2 _15411_ (.CLK(clknet_leaf_72_clk),
    .D(_02026_),
    .Q(\core_pipeline.decode_to_execute_pc[13] ));
 sky130_fd_sc_hd__dfxtp_2 _15412_ (.CLK(clknet_leaf_76_clk),
    .D(_02027_),
    .Q(\core_pipeline.decode_to_execute_pc[14] ));
 sky130_fd_sc_hd__dfxtp_2 _15413_ (.CLK(clknet_leaf_71_clk),
    .D(_02028_),
    .Q(\core_pipeline.decode_to_execute_pc[15] ));
 sky130_fd_sc_hd__dfxtp_2 _15414_ (.CLK(clknet_leaf_72_clk),
    .D(_02029_),
    .Q(\core_pipeline.decode_to_execute_pc[16] ));
 sky130_fd_sc_hd__dfxtp_4 _15415_ (.CLK(clknet_leaf_109_clk),
    .D(_02030_),
    .Q(\core_pipeline.decode_to_execute_pc[17] ));
 sky130_fd_sc_hd__dfxtp_4 _15416_ (.CLK(clknet_leaf_110_clk),
    .D(_02031_),
    .Q(\core_pipeline.decode_to_execute_pc[18] ));
 sky130_fd_sc_hd__dfxtp_2 _15417_ (.CLK(clknet_leaf_107_clk),
    .D(_02032_),
    .Q(\core_pipeline.decode_to_execute_pc[19] ));
 sky130_fd_sc_hd__dfxtp_2 _15418_ (.CLK(clknet_leaf_116_clk),
    .D(_02033_),
    .Q(\core_pipeline.decode_to_execute_pc[20] ));
 sky130_fd_sc_hd__dfxtp_2 _15419_ (.CLK(clknet_leaf_101_clk),
    .D(_02034_),
    .Q(\core_pipeline.decode_to_execute_pc[21] ));
 sky130_fd_sc_hd__dfxtp_2 _15420_ (.CLK(clknet_leaf_101_clk),
    .D(_02035_),
    .Q(\core_pipeline.decode_to_execute_pc[22] ));
 sky130_fd_sc_hd__dfxtp_2 _15421_ (.CLK(clknet_leaf_79_clk),
    .D(_02036_),
    .Q(\core_pipeline.decode_to_execute_pc[23] ));
 sky130_fd_sc_hd__dfxtp_1 _15422_ (.CLK(clknet_leaf_82_clk),
    .D(_02037_),
    .Q(\core_pipeline.decode_to_execute_pc[24] ));
 sky130_fd_sc_hd__dfxtp_1 _15423_ (.CLK(clknet_leaf_78_clk),
    .D(_02038_),
    .Q(\core_pipeline.decode_to_execute_pc[25] ));
 sky130_fd_sc_hd__dfxtp_2 _15424_ (.CLK(clknet_leaf_103_clk),
    .D(_02039_),
    .Q(\core_pipeline.decode_to_execute_pc[26] ));
 sky130_fd_sc_hd__dfxtp_2 _15425_ (.CLK(clknet_leaf_97_clk),
    .D(_02040_),
    .Q(\core_pipeline.decode_to_execute_pc[27] ));
 sky130_fd_sc_hd__dfxtp_2 _15426_ (.CLK(clknet_leaf_97_clk),
    .D(_02041_),
    .Q(\core_pipeline.decode_to_execute_pc[28] ));
 sky130_fd_sc_hd__dfxtp_1 _15427_ (.CLK(clknet_leaf_87_clk),
    .D(_02042_),
    .Q(\core_pipeline.decode_to_execute_pc[29] ));
 sky130_fd_sc_hd__dfxtp_1 _15428_ (.CLK(clknet_leaf_40_clk),
    .D(_02043_),
    .Q(\core_pipeline.decode_to_execute_pc[30] ));
 sky130_fd_sc_hd__dfxtp_2 _15429_ (.CLK(clknet_leaf_147_clk),
    .D(_02044_),
    .Q(\core_pipeline.decode_to_execute_pc[31] ));
 sky130_fd_sc_hd__dfxtp_1 _15430_ (.CLK(clknet_leaf_91_clk),
    .D(_02045_),
    .Q(\core_pipeline.decode_to_execute_next_pc[0] ));
 sky130_fd_sc_hd__dfxtp_2 _15431_ (.CLK(clknet_leaf_152_clk),
    .D(_02046_),
    .Q(\core_pipeline.decode_to_execute_next_pc[1] ));
 sky130_fd_sc_hd__dfxtp_1 _15432_ (.CLK(clknet_leaf_150_clk),
    .D(_02047_),
    .Q(\core_pipeline.decode_to_execute_next_pc[2] ));
 sky130_fd_sc_hd__dfxtp_1 _15433_ (.CLK(clknet_leaf_151_clk),
    .D(_02048_),
    .Q(\core_pipeline.decode_to_execute_next_pc[3] ));
 sky130_fd_sc_hd__dfxtp_1 _15434_ (.CLK(clknet_leaf_91_clk),
    .D(_02049_),
    .Q(\core_pipeline.decode_to_execute_next_pc[4] ));
 sky130_fd_sc_hd__dfxtp_1 _15435_ (.CLK(clknet_leaf_94_clk),
    .D(_02050_),
    .Q(\core_pipeline.decode_to_execute_next_pc[5] ));
 sky130_fd_sc_hd__dfxtp_1 _15436_ (.CLK(clknet_leaf_95_clk),
    .D(_02051_),
    .Q(\core_pipeline.decode_to_execute_next_pc[6] ));
 sky130_fd_sc_hd__dfxtp_1 _15437_ (.CLK(clknet_leaf_97_clk),
    .D(_02052_),
    .Q(\core_pipeline.decode_to_execute_next_pc[7] ));
 sky130_fd_sc_hd__dfxtp_1 _15438_ (.CLK(clknet_leaf_104_clk),
    .D(_02053_),
    .Q(\core_pipeline.decode_to_execute_next_pc[8] ));
 sky130_fd_sc_hd__dfxtp_1 _15439_ (.CLK(clknet_leaf_76_clk),
    .D(_02054_),
    .Q(\core_pipeline.decode_to_execute_next_pc[9] ));
 sky130_fd_sc_hd__dfxtp_1 _15440_ (.CLK(clknet_leaf_77_clk),
    .D(_02055_),
    .Q(\core_pipeline.decode_to_execute_next_pc[10] ));
 sky130_fd_sc_hd__dfxtp_1 _15441_ (.CLK(clknet_leaf_76_clk),
    .D(_02056_),
    .Q(\core_pipeline.decode_to_execute_next_pc[11] ));
 sky130_fd_sc_hd__dfxtp_1 _15442_ (.CLK(clknet_leaf_74_clk),
    .D(_02057_),
    .Q(\core_pipeline.decode_to_execute_next_pc[12] ));
 sky130_fd_sc_hd__dfxtp_1 _15443_ (.CLK(clknet_leaf_76_clk),
    .D(_02058_),
    .Q(\core_pipeline.decode_to_execute_next_pc[13] ));
 sky130_fd_sc_hd__dfxtp_1 _15444_ (.CLK(clknet_leaf_108_clk),
    .D(_02059_),
    .Q(\core_pipeline.decode_to_execute_next_pc[14] ));
 sky130_fd_sc_hd__dfxtp_1 _15445_ (.CLK(clknet_leaf_74_clk),
    .D(_02060_),
    .Q(\core_pipeline.decode_to_execute_next_pc[15] ));
 sky130_fd_sc_hd__dfxtp_1 _15446_ (.CLK(clknet_leaf_75_clk),
    .D(_02061_),
    .Q(\core_pipeline.decode_to_execute_next_pc[16] ));
 sky130_fd_sc_hd__dfxtp_1 _15447_ (.CLK(clknet_5_27_0_clk),
    .D(_02062_),
    .Q(\core_pipeline.decode_to_execute_next_pc[17] ));
 sky130_fd_sc_hd__dfxtp_1 _15448_ (.CLK(clknet_leaf_109_clk),
    .D(_02063_),
    .Q(\core_pipeline.decode_to_execute_next_pc[18] ));
 sky130_fd_sc_hd__dfxtp_1 _15449_ (.CLK(clknet_leaf_110_clk),
    .D(_02064_),
    .Q(\core_pipeline.decode_to_execute_next_pc[19] ));
 sky130_fd_sc_hd__dfxtp_1 _15450_ (.CLK(clknet_leaf_110_clk),
    .D(_02065_),
    .Q(\core_pipeline.decode_to_execute_next_pc[20] ));
 sky130_fd_sc_hd__dfxtp_1 _15451_ (.CLK(clknet_leaf_116_clk),
    .D(_02066_),
    .Q(\core_pipeline.decode_to_execute_next_pc[21] ));
 sky130_fd_sc_hd__dfxtp_1 _15452_ (.CLK(clknet_leaf_102_clk),
    .D(_02067_),
    .Q(\core_pipeline.decode_to_execute_next_pc[22] ));
 sky130_fd_sc_hd__dfxtp_1 _15453_ (.CLK(clknet_leaf_107_clk),
    .D(_02068_),
    .Q(\core_pipeline.decode_to_execute_next_pc[23] ));
 sky130_fd_sc_hd__dfxtp_1 _15454_ (.CLK(clknet_leaf_79_clk),
    .D(_02069_),
    .Q(\core_pipeline.decode_to_execute_next_pc[24] ));
 sky130_fd_sc_hd__dfxtp_1 _15455_ (.CLK(clknet_leaf_105_clk),
    .D(_02070_),
    .Q(\core_pipeline.decode_to_execute_next_pc[25] ));
 sky130_fd_sc_hd__dfxtp_1 _15456_ (.CLK(clknet_leaf_106_clk),
    .D(_02071_),
    .Q(\core_pipeline.decode_to_execute_next_pc[26] ));
 sky130_fd_sc_hd__dfxtp_1 _15457_ (.CLK(clknet_leaf_106_clk),
    .D(_02072_),
    .Q(\core_pipeline.decode_to_execute_next_pc[27] ));
 sky130_fd_sc_hd__dfxtp_1 _15458_ (.CLK(clknet_leaf_99_clk),
    .D(_02073_),
    .Q(\core_pipeline.decode_to_execute_next_pc[28] ));
 sky130_fd_sc_hd__dfxtp_1 _15459_ (.CLK(clknet_leaf_96_clk),
    .D(_02074_),
    .Q(\core_pipeline.decode_to_execute_next_pc[29] ));
 sky130_fd_sc_hd__dfxtp_1 _15460_ (.CLK(clknet_leaf_95_clk),
    .D(_02075_),
    .Q(\core_pipeline.decode_to_execute_next_pc[30] ));
 sky130_fd_sc_hd__dfxtp_1 _15461_ (.CLK(clknet_leaf_146_clk),
    .D(_02076_),
    .Q(\core_pipeline.decode_to_execute_next_pc[31] ));
 sky130_fd_sc_hd__dfxtp_1 _15462_ (.CLK(clknet_leaf_38_clk),
    .D(_02077_),
    .Q(\core_pipeline.decode_to_execute_rs1_bypass[0] ));
 sky130_fd_sc_hd__dfxtp_1 _15463_ (.CLK(clknet_leaf_221_clk),
    .D(_02078_),
    .Q(\core_pipeline.decode_to_execute_rs1_bypass[1] ));
 sky130_fd_sc_hd__dfxtp_1 _15464_ (.CLK(clknet_leaf_216_clk),
    .D(_02079_),
    .Q(\core_pipeline.decode_to_execute_rs1_bypass[2] ));
 sky130_fd_sc_hd__dfxtp_1 _15465_ (.CLK(clknet_leaf_26_clk),
    .D(_02080_),
    .Q(\core_pipeline.decode_to_execute_rs1_bypass[3] ));
 sky130_fd_sc_hd__dfxtp_1 _15466_ (.CLK(clknet_leaf_28_clk),
    .D(_02081_),
    .Q(\core_pipeline.decode_to_execute_rs1_bypass[4] ));
 sky130_fd_sc_hd__dfxtp_1 _15467_ (.CLK(clknet_leaf_221_clk),
    .D(_02082_),
    .Q(\core_pipeline.decode_to_execute_rs1_bypass[5] ));
 sky130_fd_sc_hd__dfxtp_1 _15468_ (.CLK(clknet_leaf_224_clk),
    .D(_02083_),
    .Q(\core_pipeline.decode_to_execute_rs1_bypass[6] ));
 sky130_fd_sc_hd__dfxtp_1 _15469_ (.CLK(clknet_leaf_30_clk),
    .D(_02084_),
    .Q(\core_pipeline.decode_to_execute_rs1_bypass[7] ));
 sky130_fd_sc_hd__dfxtp_1 _15470_ (.CLK(clknet_leaf_31_clk),
    .D(_02085_),
    .Q(\core_pipeline.decode_to_execute_rs1_bypass[8] ));
 sky130_fd_sc_hd__dfxtp_1 _15471_ (.CLK(clknet_leaf_28_clk),
    .D(_02086_),
    .Q(\core_pipeline.decode_to_execute_rs1_bypass[9] ));
 sky130_fd_sc_hd__dfxtp_1 _15472_ (.CLK(clknet_leaf_29_clk),
    .D(_02087_),
    .Q(\core_pipeline.decode_to_execute_rs1_bypass[10] ));
 sky130_fd_sc_hd__dfxtp_1 _15473_ (.CLK(clknet_leaf_27_clk),
    .D(_02088_),
    .Q(\core_pipeline.decode_to_execute_rs1_bypass[11] ));
 sky130_fd_sc_hd__dfxtp_1 _15474_ (.CLK(clknet_leaf_30_clk),
    .D(_02089_),
    .Q(\core_pipeline.decode_to_execute_rs1_bypass[12] ));
 sky130_fd_sc_hd__dfxtp_1 _15475_ (.CLK(clknet_leaf_29_clk),
    .D(_02090_),
    .Q(\core_pipeline.decode_to_execute_rs1_bypass[13] ));
 sky130_fd_sc_hd__dfxtp_1 _15476_ (.CLK(clknet_leaf_30_clk),
    .D(_02091_),
    .Q(\core_pipeline.decode_to_execute_rs1_bypass[14] ));
 sky130_fd_sc_hd__dfxtp_1 _15477_ (.CLK(clknet_leaf_30_clk),
    .D(_02092_),
    .Q(\core_pipeline.decode_to_execute_rs1_bypass[15] ));
 sky130_fd_sc_hd__dfxtp_1 _15478_ (.CLK(clknet_leaf_227_clk),
    .D(_02093_),
    .Q(\core_pipeline.decode_to_execute_rs1_bypass[16] ));
 sky130_fd_sc_hd__dfxtp_1 _15479_ (.CLK(clknet_leaf_155_clk),
    .D(_02094_),
    .Q(\core_pipeline.decode_to_execute_rs1_bypass[17] ));
 sky130_fd_sc_hd__dfxtp_1 _15480_ (.CLK(clknet_leaf_156_clk),
    .D(_02095_),
    .Q(\core_pipeline.decode_to_execute_rs1_bypass[18] ));
 sky130_fd_sc_hd__dfxtp_1 _15481_ (.CLK(clknet_leaf_155_clk),
    .D(_02096_),
    .Q(\core_pipeline.decode_to_execute_rs1_bypass[19] ));
 sky130_fd_sc_hd__dfxtp_1 _15482_ (.CLK(clknet_leaf_220_clk),
    .D(_02097_),
    .Q(\core_pipeline.decode_to_execute_rs1_bypass[20] ));
 sky130_fd_sc_hd__dfxtp_1 _15483_ (.CLK(clknet_leaf_156_clk),
    .D(_02098_),
    .Q(\core_pipeline.decode_to_execute_rs1_bypass[21] ));
 sky130_fd_sc_hd__dfxtp_1 _15484_ (.CLK(clknet_leaf_221_clk),
    .D(_02099_),
    .Q(\core_pipeline.decode_to_execute_rs1_bypass[22] ));
 sky130_fd_sc_hd__dfxtp_1 _15485_ (.CLK(clknet_leaf_219_clk),
    .D(_02100_),
    .Q(\core_pipeline.decode_to_execute_rs1_bypass[23] ));
 sky130_fd_sc_hd__dfxtp_1 _15486_ (.CLK(clknet_leaf_223_clk),
    .D(_02101_),
    .Q(\core_pipeline.decode_to_execute_rs1_bypass[24] ));
 sky130_fd_sc_hd__dfxtp_1 _15487_ (.CLK(clknet_leaf_31_clk),
    .D(_02102_),
    .Q(\core_pipeline.decode_to_execute_rs1_bypass[25] ));
 sky130_fd_sc_hd__dfxtp_1 _15488_ (.CLK(clknet_leaf_30_clk),
    .D(_02103_),
    .Q(\core_pipeline.decode_to_execute_rs1_bypass[26] ));
 sky130_fd_sc_hd__dfxtp_1 _15489_ (.CLK(clknet_leaf_156_clk),
    .D(_02104_),
    .Q(\core_pipeline.decode_to_execute_rs1_bypass[27] ));
 sky130_fd_sc_hd__dfxtp_1 _15490_ (.CLK(clknet_leaf_215_clk),
    .D(_02105_),
    .Q(\core_pipeline.decode_to_execute_rs1_bypass[28] ));
 sky130_fd_sc_hd__dfxtp_1 _15491_ (.CLK(clknet_leaf_221_clk),
    .D(_02106_),
    .Q(\core_pipeline.decode_to_execute_rs1_bypass[29] ));
 sky130_fd_sc_hd__dfxtp_1 _15492_ (.CLK(clknet_leaf_221_clk),
    .D(_02107_),
    .Q(\core_pipeline.decode_to_execute_rs1_bypass[30] ));
 sky130_fd_sc_hd__dfxtp_1 _15493_ (.CLK(clknet_leaf_155_clk),
    .D(_02108_),
    .Q(\core_pipeline.decode_to_execute_rs1_bypass[31] ));
 sky130_fd_sc_hd__dfxtp_1 _15494_ (.CLK(clknet_leaf_28_clk),
    .D(_02109_),
    .Q(\core_pipeline.decode_to_execute_rs2_bypass[0] ));
 sky130_fd_sc_hd__dfxtp_1 _15495_ (.CLK(clknet_leaf_221_clk),
    .D(_02110_),
    .Q(\core_pipeline.decode_to_execute_rs2_bypass[1] ));
 sky130_fd_sc_hd__dfxtp_1 _15496_ (.CLK(clknet_leaf_220_clk),
    .D(_02111_),
    .Q(\core_pipeline.decode_to_execute_rs2_bypass[2] ));
 sky130_fd_sc_hd__dfxtp_1 _15497_ (.CLK(clknet_leaf_26_clk),
    .D(_02112_),
    .Q(\core_pipeline.decode_to_execute_rs2_bypass[3] ));
 sky130_fd_sc_hd__dfxtp_1 _15498_ (.CLK(clknet_leaf_28_clk),
    .D(_02113_),
    .Q(\core_pipeline.decode_to_execute_rs2_bypass[4] ));
 sky130_fd_sc_hd__dfxtp_1 _15499_ (.CLK(clknet_leaf_221_clk),
    .D(_02114_),
    .Q(\core_pipeline.decode_to_execute_rs2_bypass[5] ));
 sky130_fd_sc_hd__dfxtp_1 _15500_ (.CLK(clknet_leaf_224_clk),
    .D(_02115_),
    .Q(\core_pipeline.decode_to_execute_rs2_bypass[6] ));
 sky130_fd_sc_hd__dfxtp_1 _15501_ (.CLK(clknet_leaf_30_clk),
    .D(_02116_),
    .Q(\core_pipeline.decode_to_execute_rs2_bypass[7] ));
 sky130_fd_sc_hd__dfxtp_1 _15502_ (.CLK(clknet_leaf_27_clk),
    .D(_02117_),
    .Q(\core_pipeline.decode_to_execute_rs2_bypass[8] ));
 sky130_fd_sc_hd__dfxtp_1 _15503_ (.CLK(clknet_leaf_27_clk),
    .D(_02118_),
    .Q(\core_pipeline.decode_to_execute_rs2_bypass[9] ));
 sky130_fd_sc_hd__dfxtp_1 _15504_ (.CLK(clknet_leaf_28_clk),
    .D(_02119_),
    .Q(\core_pipeline.decode_to_execute_rs2_bypass[10] ));
 sky130_fd_sc_hd__dfxtp_1 _15505_ (.CLK(clknet_leaf_27_clk),
    .D(_02120_),
    .Q(\core_pipeline.decode_to_execute_rs2_bypass[11] ));
 sky130_fd_sc_hd__dfxtp_1 _15506_ (.CLK(clknet_leaf_31_clk),
    .D(_02121_),
    .Q(\core_pipeline.decode_to_execute_rs2_bypass[12] ));
 sky130_fd_sc_hd__dfxtp_1 _15507_ (.CLK(clknet_leaf_28_clk),
    .D(_02122_),
    .Q(\core_pipeline.decode_to_execute_rs2_bypass[13] ));
 sky130_fd_sc_hd__dfxtp_1 _15508_ (.CLK(clknet_leaf_27_clk),
    .D(_02123_),
    .Q(\core_pipeline.decode_to_execute_rs2_bypass[14] ));
 sky130_fd_sc_hd__dfxtp_1 _15509_ (.CLK(clknet_leaf_29_clk),
    .D(_02124_),
    .Q(\core_pipeline.decode_to_execute_rs2_bypass[15] ));
 sky130_fd_sc_hd__dfxtp_1 _15510_ (.CLK(clknet_leaf_228_clk),
    .D(_02125_),
    .Q(\core_pipeline.decode_to_execute_rs2_bypass[16] ));
 sky130_fd_sc_hd__dfxtp_1 _15511_ (.CLK(clknet_leaf_155_clk),
    .D(_02126_),
    .Q(\core_pipeline.decode_to_execute_rs2_bypass[17] ));
 sky130_fd_sc_hd__dfxtp_1 _15512_ (.CLK(clknet_leaf_155_clk),
    .D(_02127_),
    .Q(\core_pipeline.decode_to_execute_rs2_bypass[18] ));
 sky130_fd_sc_hd__dfxtp_1 _15513_ (.CLK(clknet_leaf_216_clk),
    .D(_02128_),
    .Q(\core_pipeline.decode_to_execute_rs2_bypass[19] ));
 sky130_fd_sc_hd__dfxtp_1 _15514_ (.CLK(clknet_leaf_220_clk),
    .D(_02129_),
    .Q(\core_pipeline.decode_to_execute_rs2_bypass[20] ));
 sky130_fd_sc_hd__dfxtp_1 _15515_ (.CLK(clknet_leaf_155_clk),
    .D(_02130_),
    .Q(\core_pipeline.decode_to_execute_rs2_bypass[21] ));
 sky130_fd_sc_hd__dfxtp_1 _15516_ (.CLK(clknet_leaf_219_clk),
    .D(_02131_),
    .Q(\core_pipeline.decode_to_execute_rs2_bypass[22] ));
 sky130_fd_sc_hd__dfxtp_1 _15517_ (.CLK(clknet_leaf_219_clk),
    .D(_02132_),
    .Q(\core_pipeline.decode_to_execute_rs2_bypass[23] ));
 sky130_fd_sc_hd__dfxtp_1 _15518_ (.CLK(clknet_leaf_227_clk),
    .D(_02133_),
    .Q(\core_pipeline.decode_to_execute_rs2_bypass[24] ));
 sky130_fd_sc_hd__dfxtp_1 _15519_ (.CLK(clknet_leaf_31_clk),
    .D(_02134_),
    .Q(\core_pipeline.decode_to_execute_rs2_bypass[25] ));
 sky130_fd_sc_hd__dfxtp_1 _15520_ (.CLK(clknet_leaf_29_clk),
    .D(_02135_),
    .Q(\core_pipeline.decode_to_execute_rs2_bypass[26] ));
 sky130_fd_sc_hd__dfxtp_1 _15521_ (.CLK(clknet_leaf_155_clk),
    .D(_02136_),
    .Q(\core_pipeline.decode_to_execute_rs2_bypass[27] ));
 sky130_fd_sc_hd__dfxtp_1 _15522_ (.CLK(clknet_leaf_216_clk),
    .D(_02137_),
    .Q(\core_pipeline.decode_to_execute_rs2_bypass[28] ));
 sky130_fd_sc_hd__dfxtp_1 _15523_ (.CLK(clknet_leaf_220_clk),
    .D(_02138_),
    .Q(\core_pipeline.decode_to_execute_rs2_bypass[29] ));
 sky130_fd_sc_hd__dfxtp_1 _15524_ (.CLK(clknet_leaf_225_clk),
    .D(_02139_),
    .Q(\core_pipeline.decode_to_execute_rs2_bypass[30] ));
 sky130_fd_sc_hd__dfxtp_1 _15525_ (.CLK(clknet_leaf_155_clk),
    .D(_02140_),
    .Q(\core_pipeline.decode_to_execute_rs2_bypass[31] ));
 sky130_fd_sc_hd__dfxtp_4 _15526_ (.CLK(clknet_leaf_215_clk),
    .D(_02141_),
    .Q(\core_pipeline.decode_to_execute_rs1_bypassed ));
 sky130_fd_sc_hd__dfxtp_4 _15527_ (.CLK(clknet_leaf_216_clk),
    .D(_02142_),
    .Q(\core_pipeline.decode_to_execute_rs2_bypassed ));
 sky130_fd_sc_hd__dfxtp_1 _15528_ (.CLK(clknet_leaf_223_clk),
    .D(_02143_),
    .Q(\core_pipeline.decode_to_execute_cmp_function[1] ));
 sky130_fd_sc_hd__dfxtp_1 _15529_ (.CLK(clknet_leaf_32_clk),
    .D(_02144_),
    .Q(\core_pipeline.decode_to_execute_cmp_function[2] ));
 sky130_fd_sc_hd__dfxtp_1 _15530_ (.CLK(clknet_leaf_222_clk),
    .D(_02145_),
    .Q(\core_pipeline.decode_to_execute_jump ));
 sky130_fd_sc_hd__dfxtp_1 _15531_ (.CLK(clknet_leaf_34_clk),
    .D(_02146_),
    .Q(\core_pipeline.decode_to_execute_branch ));
 sky130_fd_sc_hd__dfxtp_1 _15532_ (.CLK(clknet_leaf_158_clk),
    .D(_02147_),
    .Q(\core_pipeline.decode_to_execute_csr_readable ));
 sky130_fd_sc_hd__dfxtp_1 _15533_ (.CLK(clknet_leaf_158_clk),
    .D(_02148_),
    .Q(\core_pipeline.decode_to_execute_csr_writeable ));
 sky130_fd_sc_hd__dfxtp_1 _15534_ (.CLK(clknet_leaf_153_clk),
    .D(_02149_),
    .Q(\core_pipeline.decode_to_execute_load ));
 sky130_fd_sc_hd__dfxtp_1 _15535_ (.CLK(clknet_leaf_92_clk),
    .D(_02150_),
    .Q(\core_pipeline.decode_to_execute_store ));
 sky130_fd_sc_hd__dfxtp_1 _15536_ (.CLK(clknet_leaf_223_clk),
    .D(_02151_),
    .Q(\core_pipeline.decode_to_execute_cmp_function[0] ));
 sky130_fd_sc_hd__dfxtp_1 _15537_ (.CLK(clknet_leaf_34_clk),
    .D(_02152_),
    .Q(\core_pipeline.decode_to_execute_load_signed ));
 sky130_fd_sc_hd__dfxtp_1 _15538_ (.CLK(clknet_leaf_152_clk),
    .D(_02153_),
    .Q(\core_pipeline.decode_to_execute_mret ));
 sky130_fd_sc_hd__dfxtp_1 _15539_ (.CLK(clknet_leaf_152_clk),
    .D(_02154_),
    .Q(\core_pipeline.decode_to_execute_wfi ));
 sky130_fd_sc_hd__dfxtp_1 _15540_ (.CLK(clknet_leaf_154_clk),
    .D(_00037_),
    .Q(\core_pipeline.decode_to_execute_valid ));
 sky130_fd_sc_hd__dfxtp_1 _15541_ (.CLK(clknet_leaf_139_clk),
    .D(_02155_),
    .Q(\core_pipeline.decode_to_execute_csr_address[0] ));
 sky130_fd_sc_hd__dfxtp_1 _15542_ (.CLK(clknet_leaf_139_clk),
    .D(_02156_),
    .Q(\core_pipeline.decode_to_execute_csr_address[1] ));
 sky130_fd_sc_hd__dfxtp_1 _15543_ (.CLK(clknet_leaf_140_clk),
    .D(_02157_),
    .Q(\core_pipeline.decode_to_execute_csr_address[2] ));
 sky130_fd_sc_hd__dfxtp_1 _15544_ (.CLK(clknet_leaf_170_clk),
    .D(_02158_),
    .Q(\core_pipeline.decode_to_execute_csr_address[3] ));
 sky130_fd_sc_hd__dfxtp_1 _15545_ (.CLK(clknet_leaf_168_clk),
    .D(_02159_),
    .Q(\core_pipeline.decode_to_execute_csr_address[4] ));
 sky130_fd_sc_hd__dfxtp_1 _15546_ (.CLK(clknet_leaf_167_clk),
    .D(_02160_),
    .Q(\core_pipeline.decode_to_execute_csr_address[5] ));
 sky130_fd_sc_hd__dfxtp_1 _15547_ (.CLK(clknet_leaf_168_clk),
    .D(_02161_),
    .Q(\core_pipeline.decode_to_execute_csr_address[6] ));
 sky130_fd_sc_hd__dfxtp_1 _15548_ (.CLK(clknet_leaf_141_clk),
    .D(_02162_),
    .Q(\core_pipeline.decode_to_execute_csr_address[7] ));
 sky130_fd_sc_hd__dfxtp_1 _15549_ (.CLK(clknet_leaf_167_clk),
    .D(_02163_),
    .Q(\core_pipeline.decode_to_execute_csr_address[8] ));
 sky130_fd_sc_hd__dfxtp_1 _15550_ (.CLK(clknet_leaf_158_clk),
    .D(_02164_),
    .Q(\core_pipeline.decode_to_execute_csr_address[9] ));
 sky130_fd_sc_hd__dfxtp_1 _15551_ (.CLK(clknet_leaf_166_clk),
    .D(_02165_),
    .Q(\core_pipeline.decode_to_execute_csr_address[10] ));
 sky130_fd_sc_hd__dfxtp_1 _15552_ (.CLK(clknet_leaf_167_clk),
    .D(_02166_),
    .Q(\core_pipeline.decode_to_execute_csr_address[11] ));
 sky130_fd_sc_hd__dfxtp_1 _15553_ (.CLK(clknet_leaf_44_clk),
    .D(_02167_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_and_clr[0] ));
 sky130_fd_sc_hd__dfxtp_1 _15554_ (.CLK(clknet_leaf_48_clk),
    .D(_02168_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_and_clr[1] ));
 sky130_fd_sc_hd__dfxtp_1 _15555_ (.CLK(clknet_leaf_48_clk),
    .D(_02169_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_and_clr[2] ));
 sky130_fd_sc_hd__dfxtp_1 _15556_ (.CLK(clknet_leaf_48_clk),
    .D(_02170_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_and_clr[3] ));
 sky130_fd_sc_hd__dfxtp_1 _15557_ (.CLK(clknet_leaf_47_clk),
    .D(_02171_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_and_clr[4] ));
 sky130_fd_sc_hd__dfxtp_1 _15558_ (.CLK(clknet_leaf_47_clk),
    .D(_02172_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_and_clr[5] ));
 sky130_fd_sc_hd__dfxtp_1 _15559_ (.CLK(clknet_leaf_41_clk),
    .D(_02173_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_and_clr[6] ));
 sky130_fd_sc_hd__dfxtp_1 _15560_ (.CLK(clknet_leaf_39_clk),
    .D(_02174_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_and_clr[7] ));
 sky130_fd_sc_hd__dfxtp_1 _15561_ (.CLK(clknet_leaf_64_clk),
    .D(_02175_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_and_clr[8] ));
 sky130_fd_sc_hd__dfxtp_1 _15562_ (.CLK(clknet_leaf_62_clk),
    .D(_02176_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_and_clr[9] ));
 sky130_fd_sc_hd__dfxtp_1 _15563_ (.CLK(clknet_leaf_64_clk),
    .D(_02177_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_and_clr[10] ));
 sky130_fd_sc_hd__dfxtp_1 _15564_ (.CLK(clknet_leaf_62_clk),
    .D(_02178_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_and_clr[11] ));
 sky130_fd_sc_hd__dfxtp_1 _15565_ (.CLK(clknet_leaf_70_clk),
    .D(_02179_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_and_clr[12] ));
 sky130_fd_sc_hd__dfxtp_1 _15566_ (.CLK(clknet_leaf_62_clk),
    .D(_02180_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_and_clr[13] ));
 sky130_fd_sc_hd__dfxtp_1 _15567_ (.CLK(clknet_leaf_70_clk),
    .D(_02181_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_and_clr[14] ));
 sky130_fd_sc_hd__dfxtp_1 _15568_ (.CLK(clknet_leaf_68_clk),
    .D(_02182_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_and_clr[15] ));
 sky130_fd_sc_hd__dfxtp_1 _15569_ (.CLK(clknet_leaf_70_clk),
    .D(_02183_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_and_clr[16] ));
 sky130_fd_sc_hd__dfxtp_1 _15570_ (.CLK(clknet_leaf_64_clk),
    .D(_02184_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_and_clr[17] ));
 sky130_fd_sc_hd__dfxtp_1 _15571_ (.CLK(clknet_leaf_68_clk),
    .D(_02185_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_and_clr[18] ));
 sky130_fd_sc_hd__dfxtp_1 _15572_ (.CLK(clknet_leaf_68_clk),
    .D(_02186_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_and_clr[19] ));
 sky130_fd_sc_hd__dfxtp_1 _15573_ (.CLK(clknet_leaf_83_clk),
    .D(_02187_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_and_clr[20] ));
 sky130_fd_sc_hd__dfxtp_1 _15574_ (.CLK(clknet_leaf_42_clk),
    .D(_02188_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_and_clr[21] ));
 sky130_fd_sc_hd__dfxtp_1 _15575_ (.CLK(clknet_leaf_67_clk),
    .D(_02189_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_and_clr[22] ));
 sky130_fd_sc_hd__dfxtp_1 _15576_ (.CLK(clknet_leaf_41_clk),
    .D(_02190_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_and_clr[23] ));
 sky130_fd_sc_hd__dfxtp_1 _15577_ (.CLK(clknet_leaf_65_clk),
    .D(_02191_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_and_clr[24] ));
 sky130_fd_sc_hd__dfxtp_1 _15578_ (.CLK(clknet_leaf_67_clk),
    .D(_02192_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_and_clr[25] ));
 sky130_fd_sc_hd__dfxtp_1 _15579_ (.CLK(clknet_leaf_67_clk),
    .D(_02193_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_and_clr[26] ));
 sky130_fd_sc_hd__dfxtp_1 _15580_ (.CLK(clknet_leaf_62_clk),
    .D(_02194_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_and_clr[27] ));
 sky130_fd_sc_hd__dfxtp_1 _15581_ (.CLK(clknet_leaf_42_clk),
    .D(_02195_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_and_clr[28] ));
 sky130_fd_sc_hd__dfxtp_1 _15582_ (.CLK(clknet_leaf_55_clk),
    .D(_02196_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_and_clr[29] ));
 sky130_fd_sc_hd__dfxtp_1 _15583_ (.CLK(clknet_leaf_41_clk),
    .D(_02197_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_and_clr[30] ));
 sky130_fd_sc_hd__dfxtp_1 _15584_ (.CLK(clknet_leaf_43_clk),
    .D(_02198_),
    .Q(\core_pipeline.pipeline_execute.ex_alu.result_and_clr[31] ));
 sky130_fd_sc_hd__dfxtp_1 _15585_ (.CLK(clknet_leaf_152_clk),
    .D(_02199_),
    .Q(\core_pipeline.fetch_to_decode_pc[2] ));
 sky130_fd_sc_hd__dfxtp_1 _15586_ (.CLK(clknet_leaf_93_clk),
    .D(_02200_),
    .Q(\core_pipeline.fetch_to_decode_pc[3] ));
 sky130_fd_sc_hd__dfxtp_1 _15587_ (.CLK(clknet_leaf_39_clk),
    .D(_02201_),
    .Q(\core_pipeline.fetch_to_decode_pc[4] ));
 sky130_fd_sc_hd__dfxtp_1 _15588_ (.CLK(clknet_leaf_36_clk),
    .D(_02202_),
    .Q(\core_pipeline.fetch_to_decode_pc[5] ));
 sky130_fd_sc_hd__dfxtp_1 _15589_ (.CLK(clknet_leaf_40_clk),
    .D(_02203_),
    .Q(\core_pipeline.fetch_to_decode_pc[6] ));
 sky130_fd_sc_hd__dfxtp_1 _15590_ (.CLK(clknet_leaf_94_clk),
    .D(_02204_),
    .Q(\core_pipeline.fetch_to_decode_pc[7] ));
 sky130_fd_sc_hd__dfxtp_1 _15591_ (.CLK(clknet_leaf_83_clk),
    .D(_02205_),
    .Q(\core_pipeline.fetch_to_decode_pc[8] ));
 sky130_fd_sc_hd__dfxtp_1 _15592_ (.CLK(clknet_leaf_73_clk),
    .D(_02206_),
    .Q(\core_pipeline.fetch_to_decode_pc[9] ));
 sky130_fd_sc_hd__dfxtp_1 _15593_ (.CLK(clknet_leaf_77_clk),
    .D(_02207_),
    .Q(\core_pipeline.fetch_to_decode_pc[10] ));
 sky130_fd_sc_hd__dfxtp_1 _15594_ (.CLK(clknet_leaf_71_clk),
    .D(_02208_),
    .Q(\core_pipeline.fetch_to_decode_pc[11] ));
 sky130_fd_sc_hd__dfxtp_1 _15595_ (.CLK(clknet_leaf_71_clk),
    .D(_02209_),
    .Q(\core_pipeline.fetch_to_decode_pc[12] ));
 sky130_fd_sc_hd__dfxtp_1 _15596_ (.CLK(clknet_leaf_72_clk),
    .D(_02210_),
    .Q(\core_pipeline.fetch_to_decode_pc[13] ));
 sky130_fd_sc_hd__dfxtp_1 _15597_ (.CLK(clknet_leaf_76_clk),
    .D(_02211_),
    .Q(\core_pipeline.fetch_to_decode_pc[14] ));
 sky130_fd_sc_hd__dfxtp_1 _15598_ (.CLK(clknet_leaf_71_clk),
    .D(_02212_),
    .Q(\core_pipeline.fetch_to_decode_pc[15] ));
 sky130_fd_sc_hd__dfxtp_1 _15599_ (.CLK(clknet_leaf_71_clk),
    .D(_02213_),
    .Q(\core_pipeline.fetch_to_decode_pc[16] ));
 sky130_fd_sc_hd__dfxtp_1 _15600_ (.CLK(clknet_leaf_109_clk),
    .D(_02214_),
    .Q(\core_pipeline.fetch_to_decode_pc[17] ));
 sky130_fd_sc_hd__dfxtp_1 _15601_ (.CLK(clknet_leaf_110_clk),
    .D(_02215_),
    .Q(\core_pipeline.fetch_to_decode_pc[18] ));
 sky130_fd_sc_hd__dfxtp_1 _15602_ (.CLK(clknet_leaf_106_clk),
    .D(_02216_),
    .Q(\core_pipeline.fetch_to_decode_pc[19] ));
 sky130_fd_sc_hd__dfxtp_1 _15603_ (.CLK(clknet_leaf_116_clk),
    .D(_02217_),
    .Q(\core_pipeline.fetch_to_decode_pc[20] ));
 sky130_fd_sc_hd__dfxtp_1 _15604_ (.CLK(clknet_leaf_101_clk),
    .D(_02218_),
    .Q(\core_pipeline.fetch_to_decode_pc[21] ));
 sky130_fd_sc_hd__dfxtp_1 _15605_ (.CLK(clknet_leaf_101_clk),
    .D(_02219_),
    .Q(\core_pipeline.fetch_to_decode_pc[22] ));
 sky130_fd_sc_hd__dfxtp_1 _15606_ (.CLK(clknet_leaf_79_clk),
    .D(_02220_),
    .Q(\core_pipeline.fetch_to_decode_pc[23] ));
 sky130_fd_sc_hd__dfxtp_1 _15607_ (.CLK(clknet_leaf_81_clk),
    .D(_02221_),
    .Q(\core_pipeline.fetch_to_decode_pc[24] ));
 sky130_fd_sc_hd__dfxtp_1 _15608_ (.CLK(clknet_leaf_78_clk),
    .D(_02222_),
    .Q(\core_pipeline.fetch_to_decode_pc[25] ));
 sky130_fd_sc_hd__dfxtp_1 _15609_ (.CLK(clknet_leaf_105_clk),
    .D(_02223_),
    .Q(\core_pipeline.fetch_to_decode_pc[26] ));
 sky130_fd_sc_hd__dfxtp_1 _15610_ (.CLK(clknet_leaf_96_clk),
    .D(_02224_),
    .Q(\core_pipeline.fetch_to_decode_pc[27] ));
 sky130_fd_sc_hd__dfxtp_1 _15611_ (.CLK(clknet_leaf_97_clk),
    .D(_02225_),
    .Q(\core_pipeline.fetch_to_decode_pc[28] ));
 sky130_fd_sc_hd__dfxtp_1 _15612_ (.CLK(clknet_leaf_87_clk),
    .D(_02226_),
    .Q(\core_pipeline.fetch_to_decode_pc[29] ));
 sky130_fd_sc_hd__dfxtp_1 _15613_ (.CLK(clknet_leaf_41_clk),
    .D(_02227_),
    .Q(\core_pipeline.fetch_to_decode_pc[30] ));
 sky130_fd_sc_hd__dfxtp_1 _15614_ (.CLK(clknet_leaf_98_clk),
    .D(_02228_),
    .Q(\core_pipeline.fetch_to_decode_pc[31] ));
 sky130_fd_sc_hd__dfxtp_4 _15615_ (.CLK(clknet_leaf_149_clk),
    .D(_00004_),
    .Q(\core_pipeline.fetch_to_decode_valid ));
 sky130_fd_sc_hd__dfxtp_1 _15616_ (.CLK(clknet_leaf_92_clk),
    .D(_02229_),
    .Q(\core_pipeline.fetch_to_decode_next_pc[0] ));
 sky130_fd_sc_hd__dfxtp_1 _15617_ (.CLK(clknet_leaf_152_clk),
    .D(_02230_),
    .Q(\core_pipeline.fetch_to_decode_next_pc[1] ));
 sky130_fd_sc_hd__dfxtp_1 _15618_ (.CLK(clknet_leaf_150_clk),
    .D(_02231_),
    .Q(\core_pipeline.fetch_to_decode_next_pc[2] ));
 sky130_fd_sc_hd__dfxtp_1 _15619_ (.CLK(clknet_leaf_151_clk),
    .D(_02232_),
    .Q(\core_pipeline.fetch_to_decode_next_pc[3] ));
 sky130_fd_sc_hd__dfxtp_1 _15620_ (.CLK(clknet_leaf_93_clk),
    .D(_02233_),
    .Q(\core_pipeline.fetch_to_decode_next_pc[4] ));
 sky130_fd_sc_hd__dfxtp_1 _15621_ (.CLK(clknet_leaf_94_clk),
    .D(_02234_),
    .Q(\core_pipeline.fetch_to_decode_next_pc[5] ));
 sky130_fd_sc_hd__dfxtp_1 _15622_ (.CLK(clknet_leaf_95_clk),
    .D(_02235_),
    .Q(\core_pipeline.fetch_to_decode_next_pc[6] ));
 sky130_fd_sc_hd__dfxtp_1 _15623_ (.CLK(clknet_leaf_97_clk),
    .D(_02236_),
    .Q(\core_pipeline.fetch_to_decode_next_pc[7] ));
 sky130_fd_sc_hd__dfxtp_1 _15624_ (.CLK(clknet_leaf_103_clk),
    .D(_02237_),
    .Q(\core_pipeline.fetch_to_decode_next_pc[8] ));
 sky130_fd_sc_hd__dfxtp_1 _15625_ (.CLK(clknet_leaf_77_clk),
    .D(_02238_),
    .Q(\core_pipeline.fetch_to_decode_next_pc[9] ));
 sky130_fd_sc_hd__dfxtp_1 _15626_ (.CLK(clknet_leaf_77_clk),
    .D(_02239_),
    .Q(\core_pipeline.fetch_to_decode_next_pc[10] ));
 sky130_fd_sc_hd__dfxtp_1 _15627_ (.CLK(clknet_leaf_76_clk),
    .D(_02240_),
    .Q(\core_pipeline.fetch_to_decode_next_pc[11] ));
 sky130_fd_sc_hd__dfxtp_1 _15628_ (.CLK(clknet_leaf_74_clk),
    .D(_02241_),
    .Q(\core_pipeline.fetch_to_decode_next_pc[12] ));
 sky130_fd_sc_hd__dfxtp_1 _15629_ (.CLK(clknet_leaf_76_clk),
    .D(_02242_),
    .Q(\core_pipeline.fetch_to_decode_next_pc[13] ));
 sky130_fd_sc_hd__dfxtp_1 _15630_ (.CLK(clknet_leaf_108_clk),
    .D(_02243_),
    .Q(\core_pipeline.fetch_to_decode_next_pc[14] ));
 sky130_fd_sc_hd__dfxtp_1 _15631_ (.CLK(clknet_leaf_76_clk),
    .D(_02244_),
    .Q(\core_pipeline.fetch_to_decode_next_pc[15] ));
 sky130_fd_sc_hd__dfxtp_1 _15632_ (.CLK(clknet_leaf_76_clk),
    .D(_02245_),
    .Q(\core_pipeline.fetch_to_decode_next_pc[16] ));
 sky130_fd_sc_hd__dfxtp_1 _15633_ (.CLK(clknet_leaf_109_clk),
    .D(_02246_),
    .Q(\core_pipeline.fetch_to_decode_next_pc[17] ));
 sky130_fd_sc_hd__dfxtp_1 _15634_ (.CLK(clknet_leaf_109_clk),
    .D(_02247_),
    .Q(\core_pipeline.fetch_to_decode_next_pc[18] ));
 sky130_fd_sc_hd__dfxtp_1 _15635_ (.CLK(clknet_leaf_110_clk),
    .D(_02248_),
    .Q(\core_pipeline.fetch_to_decode_next_pc[19] ));
 sky130_fd_sc_hd__dfxtp_1 _15636_ (.CLK(clknet_leaf_115_clk),
    .D(_02249_),
    .Q(\core_pipeline.fetch_to_decode_next_pc[20] ));
 sky130_fd_sc_hd__dfxtp_1 _15637_ (.CLK(clknet_leaf_116_clk),
    .D(_02250_),
    .Q(\core_pipeline.fetch_to_decode_next_pc[21] ));
 sky130_fd_sc_hd__dfxtp_1 _15638_ (.CLK(clknet_leaf_101_clk),
    .D(_02251_),
    .Q(\core_pipeline.fetch_to_decode_next_pc[22] ));
 sky130_fd_sc_hd__dfxtp_1 _15639_ (.CLK(clknet_leaf_105_clk),
    .D(_02252_),
    .Q(\core_pipeline.fetch_to_decode_next_pc[23] ));
 sky130_fd_sc_hd__dfxtp_1 _15640_ (.CLK(clknet_leaf_106_clk),
    .D(_02253_),
    .Q(\core_pipeline.fetch_to_decode_next_pc[24] ));
 sky130_fd_sc_hd__dfxtp_1 _15641_ (.CLK(clknet_leaf_105_clk),
    .D(_02254_),
    .Q(\core_pipeline.fetch_to_decode_next_pc[25] ));
 sky130_fd_sc_hd__dfxtp_1 _15642_ (.CLK(clknet_leaf_106_clk),
    .D(_02255_),
    .Q(\core_pipeline.fetch_to_decode_next_pc[26] ));
 sky130_fd_sc_hd__dfxtp_1 _15643_ (.CLK(clknet_leaf_106_clk),
    .D(_02256_),
    .Q(\core_pipeline.fetch_to_decode_next_pc[27] ));
 sky130_fd_sc_hd__dfxtp_1 _15644_ (.CLK(clknet_leaf_99_clk),
    .D(_02257_),
    .Q(\core_pipeline.fetch_to_decode_next_pc[28] ));
 sky130_fd_sc_hd__dfxtp_1 _15645_ (.CLK(clknet_leaf_96_clk),
    .D(_02258_),
    .Q(\core_pipeline.fetch_to_decode_next_pc[29] ));
 sky130_fd_sc_hd__dfxtp_1 _15646_ (.CLK(clknet_leaf_94_clk),
    .D(_02259_),
    .Q(\core_pipeline.fetch_to_decode_next_pc[30] ));
 sky130_fd_sc_hd__dfxtp_1 _15647_ (.CLK(clknet_leaf_98_clk),
    .D(_02260_),
    .Q(\core_pipeline.fetch_to_decode_next_pc[31] ));
 sky130_fd_sc_hd__dfxtp_1 _15648_ (.CLK(clknet_leaf_158_clk),
    .D(_02261_),
    .Q(\core_pipeline.memory_to_writeback_ecause[0] ));
 sky130_fd_sc_hd__dfxtp_1 _15649_ (.CLK(clknet_leaf_250_clk),
    .D(_02262_),
    .Q(\core_pipeline.pipeline_registers.registers[18][0] ));
 sky130_fd_sc_hd__dfxtp_1 _15650_ (.CLK(clknet_leaf_161_clk),
    .D(_02263_),
    .Q(\core_pipeline.pipeline_registers.registers[18][1] ));
 sky130_fd_sc_hd__dfxtp_1 _15651_ (.CLK(clknet_leaf_197_clk),
    .D(_02264_),
    .Q(\core_pipeline.pipeline_registers.registers[18][2] ));
 sky130_fd_sc_hd__dfxtp_1 _15652_ (.CLK(clknet_leaf_235_clk),
    .D(_02265_),
    .Q(\core_pipeline.pipeline_registers.registers[18][3] ));
 sky130_fd_sc_hd__dfxtp_1 _15653_ (.CLK(clknet_leaf_5_clk),
    .D(_02266_),
    .Q(\core_pipeline.pipeline_registers.registers[18][4] ));
 sky130_fd_sc_hd__dfxtp_1 _15654_ (.CLK(clknet_leaf_198_clk),
    .D(_02267_),
    .Q(\core_pipeline.pipeline_registers.registers[18][5] ));
 sky130_fd_sc_hd__dfxtp_1 _15655_ (.CLK(clknet_leaf_206_clk),
    .D(_02268_),
    .Q(\core_pipeline.pipeline_registers.registers[18][6] ));
 sky130_fd_sc_hd__dfxtp_1 _15656_ (.CLK(clknet_leaf_232_clk),
    .D(_02269_),
    .Q(\core_pipeline.pipeline_registers.registers[18][7] ));
 sky130_fd_sc_hd__dfxtp_1 _15657_ (.CLK(clknet_leaf_242_clk),
    .D(_02270_),
    .Q(\core_pipeline.pipeline_registers.registers[18][8] ));
 sky130_fd_sc_hd__dfxtp_1 _15658_ (.CLK(clknet_leaf_6_clk),
    .D(_02271_),
    .Q(\core_pipeline.pipeline_registers.registers[18][9] ));
 sky130_fd_sc_hd__dfxtp_1 _15659_ (.CLK(clknet_leaf_9_clk),
    .D(_02272_),
    .Q(\core_pipeline.pipeline_registers.registers[18][10] ));
 sky130_fd_sc_hd__dfxtp_1 _15660_ (.CLK(clknet_leaf_5_clk),
    .D(_02273_),
    .Q(\core_pipeline.pipeline_registers.registers[18][11] ));
 sky130_fd_sc_hd__dfxtp_1 _15661_ (.CLK(clknet_leaf_230_clk),
    .D(_02274_),
    .Q(\core_pipeline.pipeline_registers.registers[18][12] ));
 sky130_fd_sc_hd__dfxtp_1 _15662_ (.CLK(clknet_leaf_13_clk),
    .D(_02275_),
    .Q(\core_pipeline.pipeline_registers.registers[18][13] ));
 sky130_fd_sc_hd__dfxtp_1 _15663_ (.CLK(clknet_leaf_4_clk),
    .D(_02276_),
    .Q(\core_pipeline.pipeline_registers.registers[18][14] ));
 sky130_fd_sc_hd__dfxtp_1 _15664_ (.CLK(clknet_leaf_20_clk),
    .D(_02277_),
    .Q(\core_pipeline.pipeline_registers.registers[18][15] ));
 sky130_fd_sc_hd__dfxtp_1 _15665_ (.CLK(clknet_leaf_245_clk),
    .D(_02278_),
    .Q(\core_pipeline.pipeline_registers.registers[18][16] ));
 sky130_fd_sc_hd__dfxtp_1 _15666_ (.CLK(clknet_leaf_213_clk),
    .D(_02279_),
    .Q(\core_pipeline.pipeline_registers.registers[18][17] ));
 sky130_fd_sc_hd__dfxtp_1 _15667_ (.CLK(clknet_leaf_179_clk),
    .D(_02280_),
    .Q(\core_pipeline.pipeline_registers.registers[18][18] ));
 sky130_fd_sc_hd__dfxtp_1 _15668_ (.CLK(clknet_leaf_195_clk),
    .D(_02281_),
    .Q(\core_pipeline.pipeline_registers.registers[18][19] ));
 sky130_fd_sc_hd__dfxtp_1 _15669_ (.CLK(clknet_leaf_187_clk),
    .D(_02282_),
    .Q(\core_pipeline.pipeline_registers.registers[18][20] ));
 sky130_fd_sc_hd__dfxtp_1 _15670_ (.CLK(clknet_leaf_168_clk),
    .D(_02283_),
    .Q(\core_pipeline.pipeline_registers.registers[18][21] ));
 sky130_fd_sc_hd__dfxtp_1 _15671_ (.CLK(clknet_leaf_207_clk),
    .D(_02284_),
    .Q(\core_pipeline.pipeline_registers.registers[18][22] ));
 sky130_fd_sc_hd__dfxtp_1 _15672_ (.CLK(clknet_leaf_209_clk),
    .D(_02285_),
    .Q(\core_pipeline.pipeline_registers.registers[18][23] ));
 sky130_fd_sc_hd__dfxtp_1 _15673_ (.CLK(clknet_leaf_225_clk),
    .D(_02286_),
    .Q(\core_pipeline.pipeline_registers.registers[18][24] ));
 sky130_fd_sc_hd__dfxtp_1 _15674_ (.CLK(clknet_leaf_10_clk),
    .D(_02287_),
    .Q(\core_pipeline.pipeline_registers.registers[18][25] ));
 sky130_fd_sc_hd__dfxtp_1 _15675_ (.CLK(clknet_leaf_18_clk),
    .D(_02288_),
    .Q(\core_pipeline.pipeline_registers.registers[18][26] ));
 sky130_fd_sc_hd__dfxtp_1 _15676_ (.CLK(clknet_leaf_166_clk),
    .D(_02289_),
    .Q(\core_pipeline.pipeline_registers.registers[18][27] ));
 sky130_fd_sc_hd__dfxtp_1 _15677_ (.CLK(clknet_leaf_182_clk),
    .D(_02290_),
    .Q(\core_pipeline.pipeline_registers.registers[18][28] ));
 sky130_fd_sc_hd__dfxtp_1 _15678_ (.CLK(clknet_leaf_210_clk),
    .D(_02291_),
    .Q(\core_pipeline.pipeline_registers.registers[18][29] ));
 sky130_fd_sc_hd__dfxtp_1 _15679_ (.CLK(clknet_leaf_207_clk),
    .D(_02292_),
    .Q(\core_pipeline.pipeline_registers.registers[18][30] ));
 sky130_fd_sc_hd__dfxtp_1 _15680_ (.CLK(clknet_leaf_177_clk),
    .D(_02293_),
    .Q(\core_pipeline.pipeline_registers.registers[18][31] ));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_1_0_0_clk (.A(clknet_0_clk),
    .X(clknet_1_0_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_1_0_1_clk (.A(clknet_1_0_0_clk),
    .X(clknet_1_0_1_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_1_1_0_clk (.A(clknet_0_clk),
    .X(clknet_1_1_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_1_1_1_clk (.A(clknet_1_1_0_clk),
    .X(clknet_1_1_1_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_0_0_clk (.A(clknet_1_0_1_clk),
    .X(clknet_2_0_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_0_1_clk (.A(clknet_2_0_0_clk),
    .X(clknet_2_0_1_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_1_0_clk (.A(clknet_1_0_1_clk),
    .X(clknet_2_1_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_1_1_clk (.A(clknet_2_1_0_clk),
    .X(clknet_2_1_1_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_2_0_clk (.A(clknet_1_1_1_clk),
    .X(clknet_2_2_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_2_1_clk (.A(clknet_2_2_0_clk),
    .X(clknet_2_2_1_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_3_0_clk (.A(clknet_1_1_1_clk),
    .X(clknet_2_3_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_3_1_clk (.A(clknet_2_3_0_clk),
    .X(clknet_2_3_1_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_0_0_clk (.A(clknet_2_0_1_clk),
    .X(clknet_3_0_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_1_0_clk (.A(clknet_2_0_1_clk),
    .X(clknet_3_1_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_2_0_clk (.A(clknet_2_1_1_clk),
    .X(clknet_3_2_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_3_0_clk (.A(clknet_2_1_1_clk),
    .X(clknet_3_3_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_4_0_clk (.A(clknet_2_2_1_clk),
    .X(clknet_3_4_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_5_0_clk (.A(clknet_2_2_1_clk),
    .X(clknet_3_5_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_6_0_clk (.A(clknet_2_3_1_clk),
    .X(clknet_3_6_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_7_0_clk (.A(clknet_2_3_1_clk),
    .X(clknet_3_7_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_0_0_clk (.A(clknet_3_0_0_clk),
    .X(clknet_4_0_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_10_0_clk (.A(clknet_3_5_0_clk),
    .X(clknet_4_10_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_11_0_clk (.A(clknet_3_5_0_clk),
    .X(clknet_4_11_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_12_0_clk (.A(clknet_3_6_0_clk),
    .X(clknet_4_12_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_13_0_clk (.A(clknet_3_6_0_clk),
    .X(clknet_4_13_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_14_0_clk (.A(clknet_3_7_0_clk),
    .X(clknet_4_14_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_15_0_clk (.A(clknet_3_7_0_clk),
    .X(clknet_4_15_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_1_0_clk (.A(clknet_3_0_0_clk),
    .X(clknet_4_1_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_2_0_clk (.A(clknet_3_1_0_clk),
    .X(clknet_4_2_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_3_0_clk (.A(clknet_3_1_0_clk),
    .X(clknet_4_3_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_4_0_clk (.A(clknet_3_2_0_clk),
    .X(clknet_4_4_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_5_0_clk (.A(clknet_3_2_0_clk),
    .X(clknet_4_5_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_6_0_clk (.A(clknet_3_3_0_clk),
    .X(clknet_4_6_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_7_0_clk (.A(clknet_3_3_0_clk),
    .X(clknet_4_7_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_8_0_clk (.A(clknet_3_4_0_clk),
    .X(clknet_4_8_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_9_0_clk (.A(clknet_3_4_0_clk),
    .X(clknet_4_9_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_5_0_0_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_0_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_5_10_0_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_10_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_5_11_0_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_11_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_5_12_0_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_12_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_5_13_0_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_13_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_5_14_0_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_14_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_5_15_0_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_15_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_5_16_0_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_16_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_5_17_0_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_17_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_5_18_0_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_18_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_5_19_0_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_19_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_5_1_0_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_1_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_5_20_0_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_20_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_5_21_0_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_21_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_5_22_0_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_22_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_5_23_0_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_23_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_5_24_0_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_24_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_5_25_0_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_25_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_5_26_0_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_26_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_5_27_0_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_27_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_5_28_0_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_28_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_5_29_0_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_29_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_5_2_0_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_2_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_5_30_0_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_30_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_5_31_0_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_31_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_5_3_0_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_3_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_5_4_0_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_4_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_5_5_0_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_5_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_5_6_0_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_6_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_5_7_0_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_7_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_5_8_0_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_8_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_5_9_0_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_9_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_0_clk (.A(clknet_5_0_0_clk),
    .X(clknet_leaf_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_100_clk (.A(clknet_5_27_0_clk),
    .X(clknet_leaf_100_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_101_clk (.A(clknet_5_27_0_clk),
    .X(clknet_leaf_101_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_102_clk (.A(clknet_5_26_0_clk),
    .X(clknet_leaf_102_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_103_clk (.A(clknet_5_26_0_clk),
    .X(clknet_leaf_103_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_104_clk (.A(clknet_5_26_0_clk),
    .X(clknet_leaf_104_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_105_clk (.A(clknet_5_26_0_clk),
    .X(clknet_leaf_105_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_106_clk (.A(clknet_5_26_0_clk),
    .X(clknet_leaf_106_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_107_clk (.A(clknet_5_26_0_clk),
    .X(clknet_leaf_107_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_108_clk (.A(clknet_5_26_0_clk),
    .X(clknet_leaf_108_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_109_clk (.A(clknet_5_26_0_clk),
    .X(clknet_leaf_109_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_10_clk (.A(clknet_5_2_0_clk),
    .X(clknet_leaf_10_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_110_clk (.A(clknet_5_26_0_clk),
    .X(clknet_leaf_110_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_111_clk (.A(clknet_5_27_0_clk),
    .X(clknet_leaf_111_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_113_clk (.A(clknet_5_27_0_clk),
    .X(clknet_leaf_113_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_114_clk (.A(clknet_5_27_0_clk),
    .X(clknet_leaf_114_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_115_clk (.A(clknet_5_27_0_clk),
    .X(clknet_leaf_115_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_116_clk (.A(clknet_5_27_0_clk),
    .X(clknet_leaf_116_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_117_clk (.A(clknet_5_27_0_clk),
    .X(clknet_leaf_117_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_118_clk (.A(clknet_5_30_0_clk),
    .X(clknet_leaf_118_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_119_clk (.A(clknet_5_30_0_clk),
    .X(clknet_leaf_119_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_11_clk (.A(clknet_5_2_0_clk),
    .X(clknet_leaf_11_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_120_clk (.A(clknet_5_30_0_clk),
    .X(clknet_leaf_120_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_121_clk (.A(clknet_5_30_0_clk),
    .X(clknet_leaf_121_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_122_clk (.A(clknet_5_30_0_clk),
    .X(clknet_leaf_122_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_123_clk (.A(clknet_5_31_0_clk),
    .X(clknet_leaf_123_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_124_clk (.A(clknet_5_31_0_clk),
    .X(clknet_leaf_124_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_125_clk (.A(clknet_5_31_0_clk),
    .X(clknet_leaf_125_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_126_clk (.A(clknet_5_31_0_clk),
    .X(clknet_leaf_126_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_127_clk (.A(clknet_5_31_0_clk),
    .X(clknet_leaf_127_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_128_clk (.A(clknet_5_31_0_clk),
    .X(clknet_leaf_128_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_129_clk (.A(clknet_5_31_0_clk),
    .X(clknet_leaf_129_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_12_clk (.A(clknet_5_2_0_clk),
    .X(clknet_leaf_12_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_130_clk (.A(clknet_5_30_0_clk),
    .X(clknet_leaf_130_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_131_clk (.A(clknet_5_28_0_clk),
    .X(clknet_leaf_131_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_132_clk (.A(clknet_5_28_0_clk),
    .X(clknet_leaf_132_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_133_clk (.A(clknet_5_29_0_clk),
    .X(clknet_leaf_133_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_134_clk (.A(clknet_5_29_0_clk),
    .X(clknet_leaf_134_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_135_clk (.A(clknet_5_29_0_clk),
    .X(clknet_leaf_135_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_136_clk (.A(clknet_5_29_0_clk),
    .X(clknet_leaf_136_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_137_clk (.A(clknet_5_29_0_clk),
    .X(clknet_leaf_137_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_138_clk (.A(clknet_5_29_0_clk),
    .X(clknet_leaf_138_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_139_clk (.A(clknet_5_29_0_clk),
    .X(clknet_leaf_139_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_13_clk (.A(clknet_5_2_0_clk),
    .X(clknet_leaf_13_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_140_clk (.A(clknet_5_29_0_clk),
    .X(clknet_leaf_140_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_141_clk (.A(clknet_5_28_0_clk),
    .X(clknet_leaf_141_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_142_clk (.A(clknet_5_28_0_clk),
    .X(clknet_leaf_142_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_143_clk (.A(clknet_5_28_0_clk),
    .X(clknet_leaf_143_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_144_clk (.A(clknet_5_28_0_clk),
    .X(clknet_leaf_144_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_145_clk (.A(clknet_5_28_0_clk),
    .X(clknet_leaf_145_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_146_clk (.A(clknet_5_25_0_clk),
    .X(clknet_leaf_146_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_147_clk (.A(clknet_5_25_0_clk),
    .X(clknet_leaf_147_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_148_clk (.A(clknet_5_25_0_clk),
    .X(clknet_leaf_148_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_149_clk (.A(clknet_5_25_0_clk),
    .X(clknet_leaf_149_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_14_clk (.A(clknet_5_2_0_clk),
    .X(clknet_leaf_14_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_150_clk (.A(clknet_5_25_0_clk),
    .X(clknet_leaf_150_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_151_clk (.A(clknet_5_24_0_clk),
    .X(clknet_leaf_151_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_152_clk (.A(clknet_5_24_0_clk),
    .X(clknet_leaf_152_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_153_clk (.A(clknet_5_24_0_clk),
    .X(clknet_leaf_153_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_154_clk (.A(clknet_5_24_0_clk),
    .X(clknet_leaf_154_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_155_clk (.A(clknet_5_18_0_clk),
    .X(clknet_leaf_155_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_156_clk (.A(clknet_5_19_0_clk),
    .X(clknet_leaf_156_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_157_clk (.A(clknet_5_25_0_clk),
    .X(clknet_leaf_157_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_158_clk (.A(clknet_5_19_0_clk),
    .X(clknet_leaf_158_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_159_clk (.A(clknet_5_19_0_clk),
    .X(clknet_leaf_159_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_15_clk (.A(clknet_5_2_0_clk),
    .X(clknet_leaf_15_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_160_clk (.A(clknet_5_19_0_clk),
    .X(clknet_leaf_160_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_161_clk (.A(clknet_5_19_0_clk),
    .X(clknet_leaf_161_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_162_clk (.A(clknet_5_19_0_clk),
    .X(clknet_leaf_162_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_163_clk (.A(clknet_5_22_0_clk),
    .X(clknet_leaf_163_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_164_clk (.A(clknet_5_22_0_clk),
    .X(clknet_leaf_164_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_165_clk (.A(clknet_5_22_0_clk),
    .X(clknet_leaf_165_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_166_clk (.A(clknet_5_22_0_clk),
    .X(clknet_leaf_166_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_167_clk (.A(clknet_5_22_0_clk),
    .X(clknet_leaf_167_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_168_clk (.A(clknet_5_22_0_clk),
    .X(clknet_leaf_168_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_169_clk (.A(clknet_5_23_0_clk),
    .X(clknet_leaf_169_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_16_clk (.A(clknet_5_2_0_clk),
    .X(clknet_leaf_16_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_170_clk (.A(clknet_5_23_0_clk),
    .X(clknet_leaf_170_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_171_clk (.A(clknet_5_23_0_clk),
    .X(clknet_leaf_171_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_172_clk (.A(clknet_5_23_0_clk),
    .X(clknet_leaf_172_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_173_clk (.A(clknet_5_23_0_clk),
    .X(clknet_leaf_173_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_174_clk (.A(clknet_5_23_0_clk),
    .X(clknet_leaf_174_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_175_clk (.A(clknet_5_23_0_clk),
    .X(clknet_leaf_175_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_176_clk (.A(clknet_5_23_0_clk),
    .X(clknet_leaf_176_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_177_clk (.A(clknet_5_23_0_clk),
    .X(clknet_leaf_177_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_178_clk (.A(clknet_5_22_0_clk),
    .X(clknet_leaf_178_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_179_clk (.A(clknet_5_22_0_clk),
    .X(clknet_leaf_179_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_17_clk (.A(clknet_5_2_0_clk),
    .X(clknet_leaf_17_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_180_clk (.A(clknet_5_22_0_clk),
    .X(clknet_leaf_180_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_181_clk (.A(clknet_5_20_0_clk),
    .X(clknet_leaf_181_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_182_clk (.A(clknet_5_20_0_clk),
    .X(clknet_leaf_182_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_183_clk (.A(clknet_5_21_0_clk),
    .X(clknet_leaf_183_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_184_clk (.A(clknet_5_21_0_clk),
    .X(clknet_leaf_184_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_185_clk (.A(clknet_5_21_0_clk),
    .X(clknet_leaf_185_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_186_clk (.A(clknet_5_21_0_clk),
    .X(clknet_leaf_186_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_187_clk (.A(clknet_5_21_0_clk),
    .X(clknet_leaf_187_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_188_clk (.A(clknet_5_21_0_clk),
    .X(clknet_leaf_188_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_189_clk (.A(clknet_5_21_0_clk),
    .X(clknet_leaf_189_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_18_clk (.A(clknet_5_2_0_clk),
    .X(clknet_leaf_18_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_190_clk (.A(clknet_5_20_0_clk),
    .X(clknet_leaf_190_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_191_clk (.A(clknet_5_20_0_clk),
    .X(clknet_leaf_191_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_192_clk (.A(clknet_5_20_0_clk),
    .X(clknet_leaf_192_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_193_clk (.A(clknet_5_20_0_clk),
    .X(clknet_leaf_193_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_194_clk (.A(clknet_5_20_0_clk),
    .X(clknet_leaf_194_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_195_clk (.A(clknet_5_20_0_clk),
    .X(clknet_leaf_195_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_196_clk (.A(clknet_5_17_0_clk),
    .X(clknet_leaf_196_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_197_clk (.A(clknet_5_17_0_clk),
    .X(clknet_leaf_197_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_198_clk (.A(clknet_5_17_0_clk),
    .X(clknet_leaf_198_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_199_clk (.A(clknet_5_17_0_clk),
    .X(clknet_leaf_199_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_19_clk (.A(clknet_5_3_0_clk),
    .X(clknet_leaf_19_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_1_clk (.A(clknet_5_0_0_clk),
    .X(clknet_leaf_1_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_200_clk (.A(clknet_5_17_0_clk),
    .X(clknet_leaf_200_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_201_clk (.A(clknet_5_17_0_clk),
    .X(clknet_leaf_201_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_202_clk (.A(clknet_5_16_0_clk),
    .X(clknet_leaf_202_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_203_clk (.A(clknet_5_16_0_clk),
    .X(clknet_leaf_203_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_204_clk (.A(clknet_5_16_0_clk),
    .X(clknet_leaf_204_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_205_clk (.A(clknet_5_16_0_clk),
    .X(clknet_leaf_205_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_206_clk (.A(clknet_5_16_0_clk),
    .X(clknet_leaf_206_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_207_clk (.A(clknet_5_16_0_clk),
    .X(clknet_leaf_207_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_208_clk (.A(clknet_5_16_0_clk),
    .X(clknet_leaf_208_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_209_clk (.A(clknet_5_16_0_clk),
    .X(clknet_leaf_209_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_20_clk (.A(clknet_5_3_0_clk),
    .X(clknet_leaf_20_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_210_clk (.A(clknet_5_16_0_clk),
    .X(clknet_leaf_210_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_211_clk (.A(clknet_5_16_0_clk),
    .X(clknet_leaf_211_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_212_clk (.A(clknet_5_17_0_clk),
    .X(clknet_leaf_212_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_213_clk (.A(clknet_5_19_0_clk),
    .X(clknet_leaf_213_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_214_clk (.A(clknet_5_18_0_clk),
    .X(clknet_leaf_214_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_215_clk (.A(clknet_5_19_0_clk),
    .X(clknet_leaf_215_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_216_clk (.A(clknet_5_18_0_clk),
    .X(clknet_leaf_216_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_217_clk (.A(clknet_5_18_0_clk),
    .X(clknet_leaf_217_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_218_clk (.A(clknet_5_18_0_clk),
    .X(clknet_leaf_218_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_219_clk (.A(clknet_5_18_0_clk),
    .X(clknet_leaf_219_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_21_clk (.A(clknet_5_3_0_clk),
    .X(clknet_leaf_21_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_220_clk (.A(clknet_5_18_0_clk),
    .X(clknet_leaf_220_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_221_clk (.A(clknet_5_18_0_clk),
    .X(clknet_leaf_221_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_222_clk (.A(clknet_opt_1_0_clk),
    .X(clknet_leaf_222_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_223_clk (.A(clknet_5_7_0_clk),
    .X(clknet_leaf_223_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_224_clk (.A(clknet_5_7_0_clk),
    .X(clknet_leaf_224_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_225_clk (.A(clknet_5_7_0_clk),
    .X(clknet_leaf_225_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_226_clk (.A(clknet_5_7_0_clk),
    .X(clknet_leaf_226_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_227_clk (.A(clknet_5_7_0_clk),
    .X(clknet_leaf_227_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_228_clk (.A(clknet_5_6_0_clk),
    .X(clknet_leaf_228_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_229_clk (.A(clknet_5_6_0_clk),
    .X(clknet_leaf_229_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_22_clk (.A(clknet_5_3_0_clk),
    .X(clknet_leaf_22_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_230_clk (.A(clknet_5_6_0_clk),
    .X(clknet_leaf_230_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_231_clk (.A(clknet_5_4_0_clk),
    .X(clknet_leaf_231_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_232_clk (.A(clknet_5_4_0_clk),
    .X(clknet_leaf_232_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_233_clk (.A(clknet_5_4_0_clk),
    .X(clknet_leaf_233_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_234_clk (.A(clknet_5_5_0_clk),
    .X(clknet_leaf_234_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_235_clk (.A(clknet_5_5_0_clk),
    .X(clknet_leaf_235_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_236_clk (.A(clknet_5_5_0_clk),
    .X(clknet_leaf_236_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_237_clk (.A(clknet_5_5_0_clk),
    .X(clknet_leaf_237_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_238_clk (.A(clknet_5_5_0_clk),
    .X(clknet_leaf_238_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_239_clk (.A(clknet_5_5_0_clk),
    .X(clknet_leaf_239_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_23_clk (.A(clknet_5_3_0_clk),
    .X(clknet_leaf_23_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_240_clk (.A(clknet_5_5_0_clk),
    .X(clknet_leaf_240_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_241_clk (.A(clknet_5_5_0_clk),
    .X(clknet_leaf_241_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_242_clk (.A(clknet_5_5_0_clk),
    .X(clknet_leaf_242_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_243_clk (.A(clknet_5_4_0_clk),
    .X(clknet_leaf_243_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_244_clk (.A(clknet_5_4_0_clk),
    .X(clknet_leaf_244_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_245_clk (.A(clknet_5_4_0_clk),
    .X(clknet_leaf_245_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_246_clk (.A(clknet_5_4_0_clk),
    .X(clknet_leaf_246_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_247_clk (.A(clknet_5_4_0_clk),
    .X(clknet_leaf_247_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_248_clk (.A(clknet_5_4_0_clk),
    .X(clknet_leaf_248_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_249_clk (.A(clknet_5_1_0_clk),
    .X(clknet_leaf_249_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_24_clk (.A(clknet_5_3_0_clk),
    .X(clknet_leaf_24_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_250_clk (.A(clknet_5_1_0_clk),
    .X(clknet_leaf_250_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_251_clk (.A(clknet_5_1_0_clk),
    .X(clknet_leaf_251_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_252_clk (.A(clknet_5_1_0_clk),
    .X(clknet_leaf_252_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_253_clk (.A(clknet_5_1_0_clk),
    .X(clknet_leaf_253_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_254_clk (.A(clknet_5_0_0_clk),
    .X(clknet_leaf_254_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_255_clk (.A(clknet_5_0_0_clk),
    .X(clknet_leaf_255_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_256_clk (.A(clknet_5_0_0_clk),
    .X(clknet_leaf_256_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_25_clk (.A(clknet_5_6_0_clk),
    .X(clknet_leaf_25_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_26_clk (.A(clknet_5_6_0_clk),
    .X(clknet_leaf_26_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_27_clk (.A(clknet_5_6_0_clk),
    .X(clknet_leaf_27_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_28_clk (.A(clknet_5_6_0_clk),
    .X(clknet_leaf_28_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_29_clk (.A(clknet_opt_2_0_clk),
    .X(clknet_leaf_29_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_2_clk (.A(clknet_5_0_0_clk),
    .X(clknet_leaf_2_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_30_clk (.A(clknet_5_6_0_clk),
    .X(clknet_leaf_30_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_31_clk (.A(clknet_5_7_0_clk),
    .X(clknet_leaf_31_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_32_clk (.A(clknet_5_7_0_clk),
    .X(clknet_leaf_32_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_33_clk (.A(clknet_5_13_0_clk),
    .X(clknet_leaf_33_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_34_clk (.A(clknet_5_13_0_clk),
    .X(clknet_leaf_34_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_35_clk (.A(clknet_5_13_0_clk),
    .X(clknet_leaf_35_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_36_clk (.A(clknet_5_12_0_clk),
    .X(clknet_leaf_36_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_37_clk (.A(clknet_5_12_0_clk),
    .X(clknet_leaf_37_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_38_clk (.A(clknet_5_9_0_clk),
    .X(clknet_leaf_38_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_39_clk (.A(clknet_5_12_0_clk),
    .X(clknet_leaf_39_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_3_clk (.A(clknet_5_0_0_clk),
    .X(clknet_leaf_3_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_40_clk (.A(clknet_5_12_0_clk),
    .X(clknet_leaf_40_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_41_clk (.A(clknet_5_9_0_clk),
    .X(clknet_leaf_41_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_42_clk (.A(clknet_5_9_0_clk),
    .X(clknet_leaf_42_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_43_clk (.A(clknet_5_9_0_clk),
    .X(clknet_leaf_43_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_44_clk (.A(clknet_5_9_0_clk),
    .X(clknet_leaf_44_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_45_clk (.A(clknet_5_9_0_clk),
    .X(clknet_leaf_45_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_46_clk (.A(clknet_5_9_0_clk),
    .X(clknet_leaf_46_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_47_clk (.A(clknet_5_8_0_clk),
    .X(clknet_leaf_47_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_48_clk (.A(clknet_5_8_0_clk),
    .X(clknet_leaf_48_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_49_clk (.A(clknet_5_8_0_clk),
    .X(clknet_leaf_49_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_4_clk (.A(clknet_5_0_0_clk),
    .X(clknet_leaf_4_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_50_clk (.A(clknet_5_8_0_clk),
    .X(clknet_leaf_50_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_51_clk (.A(clknet_5_8_0_clk),
    .X(clknet_leaf_51_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_52_clk (.A(clknet_5_8_0_clk),
    .X(clknet_leaf_52_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_54_clk (.A(clknet_5_8_0_clk),
    .X(clknet_leaf_54_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_55_clk (.A(clknet_5_11_0_clk),
    .X(clknet_leaf_55_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_56_clk (.A(clknet_5_11_0_clk),
    .X(clknet_leaf_56_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_57_clk (.A(clknet_5_11_0_clk),
    .X(clknet_leaf_57_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_58_clk (.A(clknet_5_10_0_clk),
    .X(clknet_leaf_58_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_59_clk (.A(clknet_5_10_0_clk),
    .X(clknet_leaf_59_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_5_clk (.A(clknet_5_1_0_clk),
    .X(clknet_leaf_5_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_60_clk (.A(clknet_5_10_0_clk),
    .X(clknet_leaf_60_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_61_clk (.A(clknet_5_10_0_clk),
    .X(clknet_leaf_61_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_62_clk (.A(clknet_5_10_0_clk),
    .X(clknet_leaf_62_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_63_clk (.A(clknet_5_11_0_clk),
    .X(clknet_leaf_63_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_64_clk (.A(clknet_5_11_0_clk),
    .X(clknet_leaf_64_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_65_clk (.A(clknet_5_11_0_clk),
    .X(clknet_leaf_65_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_66_clk (.A(clknet_5_11_0_clk),
    .X(clknet_leaf_66_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_67_clk (.A(clknet_5_11_0_clk),
    .X(clknet_leaf_67_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_68_clk (.A(clknet_5_14_0_clk),
    .X(clknet_leaf_68_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_69_clk (.A(clknet_5_14_0_clk),
    .X(clknet_leaf_69_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_6_clk (.A(clknet_5_1_0_clk),
    .X(clknet_leaf_6_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_70_clk (.A(clknet_5_14_0_clk),
    .X(clknet_leaf_70_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_71_clk (.A(clknet_5_14_0_clk),
    .X(clknet_leaf_71_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_72_clk (.A(clknet_5_14_0_clk),
    .X(clknet_leaf_72_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_73_clk (.A(clknet_5_14_0_clk),
    .X(clknet_leaf_73_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_74_clk (.A(clknet_5_15_0_clk),
    .X(clknet_leaf_74_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_75_clk (.A(clknet_5_15_0_clk),
    .X(clknet_leaf_75_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_76_clk (.A(clknet_5_15_0_clk),
    .X(clknet_leaf_76_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_77_clk (.A(clknet_5_15_0_clk),
    .X(clknet_leaf_77_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_78_clk (.A(clknet_5_15_0_clk),
    .X(clknet_leaf_78_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_79_clk (.A(clknet_5_15_0_clk),
    .X(clknet_leaf_79_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_7_clk (.A(clknet_5_1_0_clk),
    .X(clknet_leaf_7_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_80_clk (.A(clknet_5_15_0_clk),
    .X(clknet_leaf_80_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_81_clk (.A(clknet_5_15_0_clk),
    .X(clknet_leaf_81_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_82_clk (.A(clknet_5_15_0_clk),
    .X(clknet_leaf_82_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_83_clk (.A(clknet_5_14_0_clk),
    .X(clknet_leaf_83_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_84_clk (.A(clknet_5_12_0_clk),
    .X(clknet_leaf_84_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_85_clk (.A(clknet_5_12_0_clk),
    .X(clknet_leaf_85_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_86_clk (.A(clknet_5_13_0_clk),
    .X(clknet_leaf_86_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_87_clk (.A(clknet_5_13_0_clk),
    .X(clknet_leaf_87_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_88_clk (.A(clknet_5_13_0_clk),
    .X(clknet_leaf_88_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_89_clk (.A(clknet_5_13_0_clk),
    .X(clknet_leaf_89_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_8_clk (.A(clknet_5_3_0_clk),
    .X(clknet_leaf_8_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_90_clk (.A(clknet_5_13_0_clk),
    .X(clknet_leaf_90_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_91_clk (.A(clknet_5_13_0_clk),
    .X(clknet_leaf_91_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_92_clk (.A(clknet_5_24_0_clk),
    .X(clknet_leaf_92_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_93_clk (.A(clknet_5_24_0_clk),
    .X(clknet_leaf_93_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_94_clk (.A(clknet_5_24_0_clk),
    .X(clknet_leaf_94_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_95_clk (.A(clknet_5_24_0_clk),
    .X(clknet_leaf_95_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_96_clk (.A(clknet_5_24_0_clk),
    .X(clknet_leaf_96_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_97_clk (.A(clknet_5_24_0_clk),
    .X(clknet_leaf_97_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_98_clk (.A(clknet_5_25_0_clk),
    .X(clknet_leaf_98_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_99_clk (.A(clknet_5_25_0_clk),
    .X(clknet_leaf_99_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_9_clk (.A(clknet_5_2_0_clk),
    .X(clknet_leaf_9_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_1_0_clk (.A(clknet_5_7_0_clk),
    .X(clknet_opt_1_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_2_0_clk (.A(clknet_5_12_0_clk),
    .X(clknet_opt_2_0_clk));
 sky130_fd_sc_hd__conb_1 core_648 (.LO(net648));
 sky130_fd_sc_hd__conb_1 core_649 (.LO(net649));
 sky130_fd_sc_hd__conb_1 core_650 (.HI(net650));
 sky130_fd_sc_hd__clkbuf_16 fanout103 (.A(net104),
    .X(net103));
 sky130_fd_sc_hd__buf_12 fanout104 (.A(_02924_),
    .X(net104));
 sky130_fd_sc_hd__buf_12 fanout105 (.A(_02923_),
    .X(net105));
 sky130_fd_sc_hd__clkbuf_8 fanout106 (.A(_02923_),
    .X(net106));
 sky130_fd_sc_hd__buf_12 fanout107 (.A(net112),
    .X(net107));
 sky130_fd_sc_hd__buf_8 fanout108 (.A(net112),
    .X(net108));
 sky130_fd_sc_hd__buf_12 fanout109 (.A(net112),
    .X(net109));
 sky130_fd_sc_hd__buf_12 fanout110 (.A(net112),
    .X(net110));
 sky130_fd_sc_hd__buf_12 fanout111 (.A(net112),
    .X(net111));
 sky130_fd_sc_hd__buf_12 fanout112 (.A(_03505_),
    .X(net112));
 sky130_fd_sc_hd__buf_12 fanout113 (.A(_03187_),
    .X(net113));
 sky130_fd_sc_hd__buf_8 fanout114 (.A(_03187_),
    .X(net114));
 sky130_fd_sc_hd__clkbuf_16 fanout115 (.A(_03124_),
    .X(net115));
 sky130_fd_sc_hd__buf_8 fanout116 (.A(_03124_),
    .X(net116));
 sky130_fd_sc_hd__clkbuf_16 fanout117 (.A(_03122_),
    .X(net117));
 sky130_fd_sc_hd__buf_8 fanout118 (.A(_03122_),
    .X(net118));
 sky130_fd_sc_hd__clkbuf_16 fanout119 (.A(_03197_),
    .X(net119));
 sky130_fd_sc_hd__buf_8 fanout120 (.A(_03197_),
    .X(net120));
 sky130_fd_sc_hd__buf_8 fanout121 (.A(net123),
    .X(net121));
 sky130_fd_sc_hd__buf_8 fanout122 (.A(net123),
    .X(net122));
 sky130_fd_sc_hd__buf_6 fanout123 (.A(net138),
    .X(net123));
 sky130_fd_sc_hd__clkbuf_16 fanout124 (.A(net138),
    .X(net124));
 sky130_fd_sc_hd__buf_6 fanout125 (.A(net138),
    .X(net125));
 sky130_fd_sc_hd__clkbuf_16 fanout126 (.A(net127),
    .X(net126));
 sky130_fd_sc_hd__buf_6 fanout127 (.A(net138),
    .X(net127));
 sky130_fd_sc_hd__buf_12 fanout128 (.A(net129),
    .X(net128));
 sky130_fd_sc_hd__buf_12 fanout129 (.A(net138),
    .X(net129));
 sky130_fd_sc_hd__clkbuf_16 fanout130 (.A(net131),
    .X(net130));
 sky130_fd_sc_hd__buf_8 fanout131 (.A(net138),
    .X(net131));
 sky130_fd_sc_hd__buf_12 fanout132 (.A(net138),
    .X(net132));
 sky130_fd_sc_hd__buf_6 fanout133 (.A(net138),
    .X(net133));
 sky130_fd_sc_hd__buf_12 fanout134 (.A(net135),
    .X(net134));
 sky130_fd_sc_hd__buf_8 fanout135 (.A(net138),
    .X(net135));
 sky130_fd_sc_hd__buf_12 fanout136 (.A(net137),
    .X(net136));
 sky130_fd_sc_hd__buf_12 fanout137 (.A(net138),
    .X(net137));
 sky130_fd_sc_hd__buf_12 fanout138 (.A(_03435_),
    .X(net138));
 sky130_fd_sc_hd__buf_12 fanout139 (.A(net148),
    .X(net139));
 sky130_fd_sc_hd__clkbuf_8 fanout140 (.A(net148),
    .X(net140));
 sky130_fd_sc_hd__buf_12 fanout141 (.A(net143),
    .X(net141));
 sky130_fd_sc_hd__clkbuf_16 fanout142 (.A(net143),
    .X(net142));
 sky130_fd_sc_hd__buf_8 fanout143 (.A(net148),
    .X(net143));
 sky130_fd_sc_hd__buf_12 fanout144 (.A(net148),
    .X(net144));
 sky130_fd_sc_hd__buf_12 fanout145 (.A(net148),
    .X(net145));
 sky130_fd_sc_hd__clkbuf_16 fanout146 (.A(net147),
    .X(net146));
 sky130_fd_sc_hd__buf_12 fanout147 (.A(net148),
    .X(net147));
 sky130_fd_sc_hd__buf_12 fanout148 (.A(_03434_),
    .X(net148));
 sky130_fd_sc_hd__buf_12 fanout149 (.A(net156),
    .X(net149));
 sky130_fd_sc_hd__buf_8 fanout150 (.A(net151),
    .X(net150));
 sky130_fd_sc_hd__buf_6 fanout151 (.A(net156),
    .X(net151));
 sky130_fd_sc_hd__buf_12 fanout152 (.A(net156),
    .X(net152));
 sky130_fd_sc_hd__buf_12 fanout153 (.A(net156),
    .X(net153));
 sky130_fd_sc_hd__buf_6 fanout154 (.A(net155),
    .X(net154));
 sky130_fd_sc_hd__buf_12 fanout155 (.A(net156),
    .X(net155));
 sky130_fd_sc_hd__buf_12 fanout156 (.A(_03434_),
    .X(net156));
 sky130_fd_sc_hd__buf_12 fanout157 (.A(net159),
    .X(net157));
 sky130_fd_sc_hd__clkbuf_16 fanout158 (.A(net159),
    .X(net158));
 sky130_fd_sc_hd__buf_12 fanout159 (.A(_03434_),
    .X(net159));
 sky130_fd_sc_hd__buf_12 fanout160 (.A(net162),
    .X(net160));
 sky130_fd_sc_hd__buf_8 fanout161 (.A(net162),
    .X(net161));
 sky130_fd_sc_hd__clkbuf_16 fanout162 (.A(_03434_),
    .X(net162));
 sky130_fd_sc_hd__buf_12 fanout163 (.A(_03311_),
    .X(net163));
 sky130_fd_sc_hd__buf_12 fanout164 (.A(_03311_),
    .X(net164));
 sky130_fd_sc_hd__buf_12 fanout165 (.A(net166),
    .X(net165));
 sky130_fd_sc_hd__buf_12 fanout166 (.A(_03111_),
    .X(net166));
 sky130_fd_sc_hd__buf_12 fanout167 (.A(_06582_),
    .X(net167));
 sky130_fd_sc_hd__buf_12 fanout168 (.A(_06582_),
    .X(net168));
 sky130_fd_sc_hd__buf_12 fanout169 (.A(_06581_),
    .X(net169));
 sky130_fd_sc_hd__buf_12 fanout170 (.A(_06581_),
    .X(net170));
 sky130_fd_sc_hd__buf_12 fanout171 (.A(_06580_),
    .X(net171));
 sky130_fd_sc_hd__buf_12 fanout172 (.A(_06580_),
    .X(net172));
 sky130_fd_sc_hd__buf_12 fanout173 (.A(_06575_),
    .X(net173));
 sky130_fd_sc_hd__buf_12 fanout174 (.A(_06575_),
    .X(net174));
 sky130_fd_sc_hd__buf_12 fanout175 (.A(_06574_),
    .X(net175));
 sky130_fd_sc_hd__buf_12 fanout176 (.A(_06574_),
    .X(net176));
 sky130_fd_sc_hd__buf_12 fanout177 (.A(_06572_),
    .X(net177));
 sky130_fd_sc_hd__buf_12 fanout178 (.A(_06572_),
    .X(net178));
 sky130_fd_sc_hd__buf_12 fanout179 (.A(_06571_),
    .X(net179));
 sky130_fd_sc_hd__buf_12 fanout180 (.A(_06571_),
    .X(net180));
 sky130_fd_sc_hd__buf_12 fanout181 (.A(_05608_),
    .X(net181));
 sky130_fd_sc_hd__buf_12 fanout182 (.A(_05608_),
    .X(net182));
 sky130_fd_sc_hd__buf_12 fanout183 (.A(_05607_),
    .X(net183));
 sky130_fd_sc_hd__buf_12 fanout184 (.A(_05607_),
    .X(net184));
 sky130_fd_sc_hd__buf_12 fanout185 (.A(_05605_),
    .X(net185));
 sky130_fd_sc_hd__buf_12 fanout186 (.A(_05605_),
    .X(net186));
 sky130_fd_sc_hd__buf_12 fanout187 (.A(_05604_),
    .X(net187));
 sky130_fd_sc_hd__buf_12 fanout188 (.A(_05604_),
    .X(net188));
 sky130_fd_sc_hd__buf_12 fanout189 (.A(_05603_),
    .X(net189));
 sky130_fd_sc_hd__buf_12 fanout190 (.A(_05603_),
    .X(net190));
 sky130_fd_sc_hd__buf_12 fanout191 (.A(_05602_),
    .X(net191));
 sky130_fd_sc_hd__buf_12 fanout192 (.A(_05602_),
    .X(net192));
 sky130_fd_sc_hd__buf_12 fanout193 (.A(_05601_),
    .X(net193));
 sky130_fd_sc_hd__buf_12 fanout194 (.A(_05601_),
    .X(net194));
 sky130_fd_sc_hd__buf_12 fanout195 (.A(_05600_),
    .X(net195));
 sky130_fd_sc_hd__buf_12 fanout196 (.A(_05600_),
    .X(net196));
 sky130_fd_sc_hd__buf_12 fanout197 (.A(_05599_),
    .X(net197));
 sky130_fd_sc_hd__buf_12 fanout198 (.A(_05599_),
    .X(net198));
 sky130_fd_sc_hd__buf_12 fanout199 (.A(_05595_),
    .X(net199));
 sky130_fd_sc_hd__buf_12 fanout200 (.A(_05595_),
    .X(net200));
 sky130_fd_sc_hd__buf_12 fanout201 (.A(_05594_),
    .X(net201));
 sky130_fd_sc_hd__buf_12 fanout202 (.A(_05594_),
    .X(net202));
 sky130_fd_sc_hd__buf_12 fanout203 (.A(_05593_),
    .X(net203));
 sky130_fd_sc_hd__buf_12 fanout204 (.A(_05593_),
    .X(net204));
 sky130_fd_sc_hd__buf_12 fanout205 (.A(_05591_),
    .X(net205));
 sky130_fd_sc_hd__buf_12 fanout206 (.A(_05591_),
    .X(net206));
 sky130_fd_sc_hd__buf_12 fanout207 (.A(_05590_),
    .X(net207));
 sky130_fd_sc_hd__buf_12 fanout208 (.A(_05590_),
    .X(net208));
 sky130_fd_sc_hd__buf_12 fanout209 (.A(_05588_),
    .X(net209));
 sky130_fd_sc_hd__buf_12 fanout210 (.A(_05588_),
    .X(net210));
 sky130_fd_sc_hd__buf_12 fanout211 (.A(_05587_),
    .X(net211));
 sky130_fd_sc_hd__buf_12 fanout212 (.A(_05587_),
    .X(net212));
 sky130_fd_sc_hd__buf_12 fanout213 (.A(_05585_),
    .X(net213));
 sky130_fd_sc_hd__buf_12 fanout214 (.A(_05585_),
    .X(net214));
 sky130_fd_sc_hd__buf_12 fanout215 (.A(_04940_),
    .X(net215));
 sky130_fd_sc_hd__buf_12 fanout216 (.A(_04940_),
    .X(net216));
 sky130_fd_sc_hd__buf_12 fanout217 (.A(_04938_),
    .X(net217));
 sky130_fd_sc_hd__buf_12 fanout218 (.A(_04938_),
    .X(net218));
 sky130_fd_sc_hd__buf_12 fanout219 (.A(_04935_),
    .X(net219));
 sky130_fd_sc_hd__buf_12 fanout220 (.A(_04935_),
    .X(net220));
 sky130_fd_sc_hd__buf_12 fanout221 (.A(_04390_),
    .X(net221));
 sky130_fd_sc_hd__buf_12 fanout222 (.A(_04390_),
    .X(net222));
 sky130_fd_sc_hd__buf_6 fanout223 (.A(net224),
    .X(net223));
 sky130_fd_sc_hd__clkbuf_16 fanout224 (.A(_04295_),
    .X(net224));
 sky130_fd_sc_hd__buf_6 fanout225 (.A(net226),
    .X(net225));
 sky130_fd_sc_hd__buf_8 fanout226 (.A(_04295_),
    .X(net226));
 sky130_fd_sc_hd__buf_6 fanout227 (.A(net228),
    .X(net227));
 sky130_fd_sc_hd__buf_6 fanout228 (.A(_04112_),
    .X(net228));
 sky130_fd_sc_hd__buf_6 fanout229 (.A(net230),
    .X(net229));
 sky130_fd_sc_hd__buf_8 fanout230 (.A(_04112_),
    .X(net230));
 sky130_fd_sc_hd__buf_8 fanout231 (.A(_04022_),
    .X(net231));
 sky130_fd_sc_hd__buf_4 fanout232 (.A(_04022_),
    .X(net232));
 sky130_fd_sc_hd__buf_6 fanout233 (.A(net234),
    .X(net233));
 sky130_fd_sc_hd__buf_8 fanout234 (.A(_04022_),
    .X(net234));
 sky130_fd_sc_hd__buf_12 fanout235 (.A(net236),
    .X(net235));
 sky130_fd_sc_hd__buf_12 fanout236 (.A(_04019_),
    .X(net236));
 sky130_fd_sc_hd__buf_12 fanout237 (.A(_03649_),
    .X(net237));
 sky130_fd_sc_hd__buf_12 fanout238 (.A(_03649_),
    .X(net238));
 sky130_fd_sc_hd__clkbuf_16 fanout239 (.A(net240),
    .X(net239));
 sky130_fd_sc_hd__buf_12 fanout240 (.A(_03114_),
    .X(net240));
 sky130_fd_sc_hd__buf_12 fanout241 (.A(_05609_),
    .X(net241));
 sky130_fd_sc_hd__buf_12 fanout242 (.A(_05609_),
    .X(net242));
 sky130_fd_sc_hd__buf_12 fanout243 (.A(_05597_),
    .X(net243));
 sky130_fd_sc_hd__buf_12 fanout244 (.A(_05597_),
    .X(net244));
 sky130_fd_sc_hd__buf_12 fanout245 (.A(net246),
    .X(net245));
 sky130_fd_sc_hd__buf_12 fanout246 (.A(_04718_),
    .X(net246));
 sky130_fd_sc_hd__buf_12 fanout247 (.A(_04717_),
    .X(net247));
 sky130_fd_sc_hd__clkbuf_16 fanout248 (.A(_04717_),
    .X(net248));
 sky130_fd_sc_hd__buf_12 fanout249 (.A(_04708_),
    .X(net249));
 sky130_fd_sc_hd__clkbuf_16 fanout250 (.A(_04708_),
    .X(net250));
 sky130_fd_sc_hd__buf_12 fanout251 (.A(_04705_),
    .X(net251));
 sky130_fd_sc_hd__clkbuf_16 fanout252 (.A(_04705_),
    .X(net252));
 sky130_fd_sc_hd__buf_12 fanout253 (.A(_04470_),
    .X(net253));
 sky130_fd_sc_hd__buf_12 fanout254 (.A(_04470_),
    .X(net254));
 sky130_fd_sc_hd__buf_6 fanout255 (.A(net256),
    .X(net255));
 sky130_fd_sc_hd__buf_8 fanout256 (.A(_04203_),
    .X(net256));
 sky130_fd_sc_hd__buf_8 fanout257 (.A(net258),
    .X(net257));
 sky130_fd_sc_hd__clkbuf_16 fanout258 (.A(_04203_),
    .X(net258));
 sky130_fd_sc_hd__buf_12 fanout259 (.A(_03916_),
    .X(net259));
 sky130_fd_sc_hd__buf_12 fanout260 (.A(_03916_),
    .X(net260));
 sky130_fd_sc_hd__buf_12 fanout261 (.A(net262),
    .X(net261));
 sky130_fd_sc_hd__buf_12 fanout262 (.A(_03429_),
    .X(net262));
 sky130_fd_sc_hd__buf_8 fanout263 (.A(net264),
    .X(net263));
 sky130_fd_sc_hd__buf_12 fanout264 (.A(_03190_),
    .X(net264));
 sky130_fd_sc_hd__buf_12 fanout265 (.A(_04719_),
    .X(net265));
 sky130_fd_sc_hd__buf_12 fanout266 (.A(_04719_),
    .X(net266));
 sky130_fd_sc_hd__buf_12 fanout267 (.A(_04711_),
    .X(net267));
 sky130_fd_sc_hd__clkbuf_16 fanout268 (.A(_04711_),
    .X(net268));
 sky130_fd_sc_hd__buf_12 fanout269 (.A(_04700_),
    .X(net269));
 sky130_fd_sc_hd__buf_8 fanout270 (.A(_04700_),
    .X(net270));
 sky130_fd_sc_hd__buf_12 fanout271 (.A(_04697_),
    .X(net271));
 sky130_fd_sc_hd__buf_6 fanout272 (.A(_04697_),
    .X(net272));
 sky130_fd_sc_hd__buf_12 fanout273 (.A(_04690_),
    .X(net273));
 sky130_fd_sc_hd__buf_6 fanout274 (.A(_04690_),
    .X(net274));
 sky130_fd_sc_hd__buf_12 fanout275 (.A(_03712_),
    .X(net275));
 sky130_fd_sc_hd__buf_12 fanout276 (.A(net277),
    .X(net276));
 sky130_fd_sc_hd__buf_12 fanout277 (.A(_04698_),
    .X(net277));
 sky130_fd_sc_hd__buf_12 fanout278 (.A(net279),
    .X(net278));
 sky130_fd_sc_hd__buf_12 fanout279 (.A(_04683_),
    .X(net279));
 sky130_fd_sc_hd__clkbuf_16 fanout280 (.A(_04481_),
    .X(net280));
 sky130_fd_sc_hd__buf_6 fanout282 (.A(net283),
    .X(net282));
 sky130_fd_sc_hd__buf_6 fanout283 (.A(_04015_),
    .X(net283));
 sky130_fd_sc_hd__buf_6 fanout284 (.A(net285),
    .X(net284));
 sky130_fd_sc_hd__buf_6 fanout285 (.A(_04012_),
    .X(net285));
 sky130_fd_sc_hd__buf_6 fanout286 (.A(net287),
    .X(net286));
 sky130_fd_sc_hd__clkbuf_4 fanout287 (.A(net288),
    .X(net287));
 sky130_fd_sc_hd__buf_4 fanout288 (.A(_04009_),
    .X(net288));
 sky130_fd_sc_hd__buf_6 fanout289 (.A(net290),
    .X(net289));
 sky130_fd_sc_hd__buf_6 fanout290 (.A(_04006_),
    .X(net290));
 sky130_fd_sc_hd__buf_6 fanout291 (.A(_04003_),
    .X(net291));
 sky130_fd_sc_hd__buf_4 fanout292 (.A(_04003_),
    .X(net292));
 sky130_fd_sc_hd__buf_6 fanout293 (.A(net294),
    .X(net293));
 sky130_fd_sc_hd__buf_8 fanout294 (.A(_04000_),
    .X(net294));
 sky130_fd_sc_hd__buf_6 fanout295 (.A(net296),
    .X(net295));
 sky130_fd_sc_hd__buf_8 fanout296 (.A(_03997_),
    .X(net296));
 sky130_fd_sc_hd__buf_6 fanout297 (.A(net298),
    .X(net297));
 sky130_fd_sc_hd__buf_6 fanout298 (.A(_03994_),
    .X(net298));
 sky130_fd_sc_hd__buf_6 fanout299 (.A(net300),
    .X(net299));
 sky130_fd_sc_hd__buf_6 fanout300 (.A(_03991_),
    .X(net300));
 sky130_fd_sc_hd__buf_6 fanout301 (.A(_03988_),
    .X(net301));
 sky130_fd_sc_hd__buf_4 fanout302 (.A(_03988_),
    .X(net302));
 sky130_fd_sc_hd__buf_6 fanout303 (.A(net304),
    .X(net303));
 sky130_fd_sc_hd__buf_6 fanout304 (.A(_03985_),
    .X(net304));
 sky130_fd_sc_hd__buf_6 fanout305 (.A(net306),
    .X(net305));
 sky130_fd_sc_hd__clkbuf_4 fanout306 (.A(net307),
    .X(net306));
 sky130_fd_sc_hd__buf_6 fanout307 (.A(_03982_),
    .X(net307));
 sky130_fd_sc_hd__buf_6 fanout308 (.A(net309),
    .X(net308));
 sky130_fd_sc_hd__buf_6 fanout309 (.A(_03979_),
    .X(net309));
 sky130_fd_sc_hd__buf_6 fanout310 (.A(_03976_),
    .X(net310));
 sky130_fd_sc_hd__buf_4 fanout311 (.A(_03976_),
    .X(net311));
 sky130_fd_sc_hd__buf_6 fanout312 (.A(net314),
    .X(net312));
 sky130_fd_sc_hd__buf_2 fanout313 (.A(net314),
    .X(net313));
 sky130_fd_sc_hd__clkbuf_8 fanout314 (.A(_03973_),
    .X(net314));
 sky130_fd_sc_hd__buf_6 fanout315 (.A(_03970_),
    .X(net315));
 sky130_fd_sc_hd__buf_4 fanout316 (.A(_03970_),
    .X(net316));
 sky130_fd_sc_hd__buf_6 fanout317 (.A(net318),
    .X(net317));
 sky130_fd_sc_hd__buf_8 fanout318 (.A(_03967_),
    .X(net318));
 sky130_fd_sc_hd__buf_6 fanout319 (.A(_03964_),
    .X(net319));
 sky130_fd_sc_hd__buf_8 fanout320 (.A(_03964_),
    .X(net320));
 sky130_fd_sc_hd__buf_6 fanout321 (.A(net322),
    .X(net321));
 sky130_fd_sc_hd__buf_8 fanout322 (.A(_03961_),
    .X(net322));
 sky130_fd_sc_hd__buf_6 fanout323 (.A(_03958_),
    .X(net323));
 sky130_fd_sc_hd__buf_4 fanout324 (.A(_03958_),
    .X(net324));
 sky130_fd_sc_hd__buf_6 fanout325 (.A(_03955_),
    .X(net325));
 sky130_fd_sc_hd__buf_6 fanout326 (.A(_03955_),
    .X(net326));
 sky130_fd_sc_hd__buf_6 fanout327 (.A(net328),
    .X(net327));
 sky130_fd_sc_hd__clkbuf_16 fanout328 (.A(_03952_),
    .X(net328));
 sky130_fd_sc_hd__buf_6 fanout329 (.A(net330),
    .X(net329));
 sky130_fd_sc_hd__buf_8 fanout330 (.A(_03949_),
    .X(net330));
 sky130_fd_sc_hd__buf_6 fanout331 (.A(_03946_),
    .X(net331));
 sky130_fd_sc_hd__buf_4 fanout332 (.A(_03946_),
    .X(net332));
 sky130_fd_sc_hd__buf_6 fanout333 (.A(net334),
    .X(net333));
 sky130_fd_sc_hd__clkbuf_16 fanout334 (.A(_03943_),
    .X(net334));
 sky130_fd_sc_hd__buf_6 fanout335 (.A(net336),
    .X(net335));
 sky130_fd_sc_hd__buf_6 fanout336 (.A(_03940_),
    .X(net336));
 sky130_fd_sc_hd__buf_6 fanout337 (.A(net339),
    .X(net337));
 sky130_fd_sc_hd__clkbuf_4 fanout338 (.A(net339),
    .X(net338));
 sky130_fd_sc_hd__buf_6 fanout339 (.A(_03937_),
    .X(net339));
 sky130_fd_sc_hd__buf_6 fanout340 (.A(net341),
    .X(net340));
 sky130_fd_sc_hd__buf_6 fanout341 (.A(_03934_),
    .X(net341));
 sky130_fd_sc_hd__buf_6 fanout342 (.A(net343),
    .X(net342));
 sky130_fd_sc_hd__buf_6 fanout343 (.A(_03931_),
    .X(net343));
 sky130_fd_sc_hd__buf_6 fanout344 (.A(_03928_),
    .X(net344));
 sky130_fd_sc_hd__buf_4 fanout345 (.A(_03928_),
    .X(net345));
 sky130_fd_sc_hd__buf_6 fanout346 (.A(net347),
    .X(net346));
 sky130_fd_sc_hd__buf_6 fanout347 (.A(_03925_),
    .X(net347));
 sky130_fd_sc_hd__buf_6 fanout348 (.A(net349),
    .X(net348));
 sky130_fd_sc_hd__buf_6 fanout349 (.A(_03922_),
    .X(net349));
 sky130_fd_sc_hd__buf_12 fanout350 (.A(net351),
    .X(net350));
 sky130_fd_sc_hd__buf_12 fanout351 (.A(_03510_),
    .X(net351));
 sky130_fd_sc_hd__buf_8 fanout352 (.A(net353),
    .X(net352));
 sky130_fd_sc_hd__buf_12 fanout353 (.A(_05842_),
    .X(net353));
 sky130_fd_sc_hd__buf_12 fanout354 (.A(net355),
    .X(net354));
 sky130_fd_sc_hd__buf_12 fanout355 (.A(_05837_),
    .X(net355));
 sky130_fd_sc_hd__buf_12 fanout356 (.A(net357),
    .X(net356));
 sky130_fd_sc_hd__buf_12 fanout357 (.A(_05831_),
    .X(net357));
 sky130_fd_sc_hd__clkbuf_16 fanout358 (.A(net359),
    .X(net358));
 sky130_fd_sc_hd__buf_12 fanout359 (.A(_05830_),
    .X(net359));
 sky130_fd_sc_hd__buf_12 fanout361 (.A(_04706_),
    .X(net361));
 sky130_fd_sc_hd__buf_12 fanout362 (.A(_04706_),
    .X(net362));
 sky130_fd_sc_hd__buf_12 fanout363 (.A(net364),
    .X(net363));
 sky130_fd_sc_hd__buf_12 fanout364 (.A(_04695_),
    .X(net364));
 sky130_fd_sc_hd__buf_12 fanout365 (.A(net366),
    .X(net365));
 sky130_fd_sc_hd__buf_12 fanout366 (.A(_04695_),
    .X(net366));
 sky130_fd_sc_hd__buf_12 fanout367 (.A(net368),
    .X(net367));
 sky130_fd_sc_hd__buf_12 fanout368 (.A(_04694_),
    .X(net368));
 sky130_fd_sc_hd__buf_12 fanout369 (.A(net370),
    .X(net369));
 sky130_fd_sc_hd__buf_12 fanout370 (.A(_04694_),
    .X(net370));
 sky130_fd_sc_hd__buf_6 fanout372 (.A(net373),
    .X(net372));
 sky130_fd_sc_hd__buf_6 fanout373 (.A(net374),
    .X(net373));
 sky130_fd_sc_hd__buf_8 fanout374 (.A(_04491_),
    .X(net374));
 sky130_fd_sc_hd__buf_6 fanout375 (.A(net376),
    .X(net375));
 sky130_fd_sc_hd__buf_6 fanout376 (.A(net377),
    .X(net376));
 sky130_fd_sc_hd__clkbuf_16 fanout377 (.A(_04490_),
    .X(net377));
 sky130_fd_sc_hd__buf_8 fanout378 (.A(net379),
    .X(net378));
 sky130_fd_sc_hd__buf_12 fanout379 (.A(_04488_),
    .X(net379));
 sky130_fd_sc_hd__buf_12 fanout380 (.A(net383),
    .X(net380));
 sky130_fd_sc_hd__clkbuf_16 fanout381 (.A(net382),
    .X(net381));
 sky130_fd_sc_hd__buf_12 fanout382 (.A(net383),
    .X(net382));
 sky130_fd_sc_hd__buf_6 fanout383 (.A(_04487_),
    .X(net383));
 sky130_fd_sc_hd__buf_12 fanout384 (.A(_04485_),
    .X(net384));
 sky130_fd_sc_hd__buf_8 fanout385 (.A(_04485_),
    .X(net385));
 sky130_fd_sc_hd__buf_12 fanout386 (.A(net388),
    .X(net386));
 sky130_fd_sc_hd__clkbuf_8 fanout387 (.A(net388),
    .X(net387));
 sky130_fd_sc_hd__buf_12 fanout388 (.A(_04484_),
    .X(net388));
 sky130_fd_sc_hd__clkbuf_16 fanout389 (.A(_04480_),
    .X(net389));
 sky130_fd_sc_hd__buf_6 fanout390 (.A(net391),
    .X(net390));
 sky130_fd_sc_hd__buf_12 fanout391 (.A(_04480_),
    .X(net391));
 sky130_fd_sc_hd__buf_8 fanout392 (.A(net393),
    .X(net392));
 sky130_fd_sc_hd__buf_12 fanout393 (.A(_04479_),
    .X(net393));
 sky130_fd_sc_hd__buf_8 fanout394 (.A(net395),
    .X(net394));
 sky130_fd_sc_hd__buf_12 fanout395 (.A(_04477_),
    .X(net395));
 sky130_fd_sc_hd__buf_8 fanout396 (.A(net398),
    .X(net396));
 sky130_fd_sc_hd__clkbuf_4 fanout397 (.A(net398),
    .X(net397));
 sky130_fd_sc_hd__buf_12 fanout398 (.A(net399),
    .X(net398));
 sky130_fd_sc_hd__buf_12 fanout399 (.A(_04476_),
    .X(net399));
 sky130_fd_sc_hd__buf_12 fanout400 (.A(net401),
    .X(net400));
 sky130_fd_sc_hd__clkbuf_16 fanout401 (.A(_03478_),
    .X(net401));
 sky130_fd_sc_hd__buf_12 fanout402 (.A(net403),
    .X(net402));
 sky130_fd_sc_hd__buf_12 fanout403 (.A(_03478_),
    .X(net403));
 sky130_fd_sc_hd__buf_6 fanout404 (.A(net405),
    .X(net404));
 sky130_fd_sc_hd__buf_8 fanout405 (.A(_03244_),
    .X(net405));
 sky130_fd_sc_hd__buf_8 fanout406 (.A(_03244_),
    .X(net406));
 sky130_fd_sc_hd__clkbuf_16 fanout407 (.A(net409),
    .X(net407));
 sky130_fd_sc_hd__buf_4 fanout408 (.A(net409),
    .X(net408));
 sky130_fd_sc_hd__buf_12 fanout409 (.A(_06315_),
    .X(net409));
 sky130_fd_sc_hd__buf_12 fanout410 (.A(net411),
    .X(net410));
 sky130_fd_sc_hd__buf_12 fanout411 (.A(_06214_),
    .X(net411));
 sky130_fd_sc_hd__buf_12 fanout412 (.A(_06025_),
    .X(net412));
 sky130_fd_sc_hd__buf_6 fanout413 (.A(_06025_),
    .X(net413));
 sky130_fd_sc_hd__clkbuf_16 fanout414 (.A(_05968_),
    .X(net414));
 sky130_fd_sc_hd__buf_8 fanout415 (.A(net417),
    .X(net415));
 sky130_fd_sc_hd__clkbuf_4 fanout416 (.A(net417),
    .X(net416));
 sky130_fd_sc_hd__buf_6 fanout417 (.A(_05968_),
    .X(net417));
 sky130_fd_sc_hd__buf_12 fanout418 (.A(net419),
    .X(net418));
 sky130_fd_sc_hd__buf_12 fanout419 (.A(_05838_),
    .X(net419));
 sky130_fd_sc_hd__buf_8 fanout420 (.A(net421),
    .X(net420));
 sky130_fd_sc_hd__buf_12 fanout421 (.A(_05835_),
    .X(net421));
 sky130_fd_sc_hd__clkbuf_16 fanout422 (.A(net423),
    .X(net422));
 sky130_fd_sc_hd__buf_12 fanout423 (.A(_05829_),
    .X(net423));
 sky130_fd_sc_hd__buf_12 fanout424 (.A(net425),
    .X(net424));
 sky130_fd_sc_hd__buf_12 fanout425 (.A(_04681_),
    .X(net425));
 sky130_fd_sc_hd__buf_12 fanout426 (.A(net427),
    .X(net426));
 sky130_fd_sc_hd__buf_12 fanout427 (.A(_04681_),
    .X(net427));
 sky130_fd_sc_hd__buf_12 fanout428 (.A(net429),
    .X(net428));
 sky130_fd_sc_hd__buf_12 fanout429 (.A(_04680_),
    .X(net429));
 sky130_fd_sc_hd__buf_12 fanout430 (.A(_04680_),
    .X(net430));
 sky130_fd_sc_hd__buf_12 fanout431 (.A(net432),
    .X(net431));
 sky130_fd_sc_hd__buf_12 fanout432 (.A(_04493_),
    .X(net432));
 sky130_fd_sc_hd__buf_12 fanout433 (.A(net434),
    .X(net433));
 sky130_fd_sc_hd__buf_12 fanout434 (.A(_04474_),
    .X(net434));
 sky130_fd_sc_hd__clkbuf_16 fanout435 (.A(_04472_),
    .X(net435));
 sky130_fd_sc_hd__buf_6 fanout436 (.A(_04472_),
    .X(net436));
 sky130_fd_sc_hd__clkbuf_16 fanout439 (.A(net440),
    .X(net439));
 sky130_fd_sc_hd__buf_12 fanout440 (.A(_03920_),
    .X(net440));
 sky130_fd_sc_hd__buf_12 fanout441 (.A(net442),
    .X(net441));
 sky130_fd_sc_hd__buf_12 fanout442 (.A(_03919_),
    .X(net442));
 sky130_fd_sc_hd__clkbuf_16 fanout443 (.A(net444),
    .X(net443));
 sky130_fd_sc_hd__buf_12 fanout444 (.A(_03918_),
    .X(net444));
 sky130_fd_sc_hd__buf_12 fanout445 (.A(_03513_),
    .X(net445));
 sky130_fd_sc_hd__buf_12 fanout446 (.A(net448),
    .X(net446));
 sky130_fd_sc_hd__clkbuf_8 fanout447 (.A(net448),
    .X(net447));
 sky130_fd_sc_hd__buf_12 fanout448 (.A(_03432_),
    .X(net448));
 sky130_fd_sc_hd__buf_12 fanout449 (.A(net450),
    .X(net449));
 sky130_fd_sc_hd__buf_12 fanout450 (.A(_03432_),
    .X(net450));
 sky130_fd_sc_hd__clkbuf_16 fanout451 (.A(net452),
    .X(net451));
 sky130_fd_sc_hd__buf_8 fanout452 (.A(net453),
    .X(net452));
 sky130_fd_sc_hd__buf_8 fanout453 (.A(_03432_),
    .X(net453));
 sky130_fd_sc_hd__buf_12 fanout454 (.A(net455),
    .X(net454));
 sky130_fd_sc_hd__buf_12 fanout455 (.A(_03432_),
    .X(net455));
 sky130_fd_sc_hd__buf_12 fanout456 (.A(_03432_),
    .X(net456));
 sky130_fd_sc_hd__buf_6 fanout457 (.A(_03432_),
    .X(net457));
 sky130_fd_sc_hd__buf_12 fanout458 (.A(_03431_),
    .X(net458));
 sky130_fd_sc_hd__buf_12 fanout459 (.A(_03423_),
    .X(net459));
 sky130_fd_sc_hd__buf_12 fanout460 (.A(net461),
    .X(net460));
 sky130_fd_sc_hd__buf_12 fanout461 (.A(_03330_),
    .X(net461));
 sky130_fd_sc_hd__buf_12 fanout462 (.A(_03329_),
    .X(net462));
 sky130_fd_sc_hd__buf_12 fanout463 (.A(_03329_),
    .X(net463));
 sky130_fd_sc_hd__buf_12 fanout464 (.A(net465),
    .X(net464));
 sky130_fd_sc_hd__buf_12 fanout465 (.A(_03329_),
    .X(net465));
 sky130_fd_sc_hd__buf_12 fanout466 (.A(net467),
    .X(net466));
 sky130_fd_sc_hd__buf_12 fanout467 (.A(_03326_),
    .X(net467));
 sky130_fd_sc_hd__buf_12 fanout468 (.A(net469),
    .X(net468));
 sky130_fd_sc_hd__buf_12 fanout469 (.A(_03325_),
    .X(net469));
 sky130_fd_sc_hd__buf_12 fanout470 (.A(net471),
    .X(net470));
 sky130_fd_sc_hd__buf_12 fanout471 (.A(_03325_),
    .X(net471));
 sky130_fd_sc_hd__buf_12 fanout472 (.A(net474),
    .X(net472));
 sky130_fd_sc_hd__buf_12 fanout473 (.A(net474),
    .X(net473));
 sky130_fd_sc_hd__clkbuf_16 fanout474 (.A(net481),
    .X(net474));
 sky130_fd_sc_hd__buf_12 fanout475 (.A(net476),
    .X(net475));
 sky130_fd_sc_hd__buf_12 fanout476 (.A(net481),
    .X(net476));
 sky130_fd_sc_hd__buf_12 fanout477 (.A(net481),
    .X(net477));
 sky130_fd_sc_hd__buf_12 fanout478 (.A(net481),
    .X(net478));
 sky130_fd_sc_hd__buf_12 fanout479 (.A(net480),
    .X(net479));
 sky130_fd_sc_hd__buf_8 fanout480 (.A(net481),
    .X(net480));
 sky130_fd_sc_hd__buf_12 fanout481 (.A(_03324_),
    .X(net481));
 sky130_fd_sc_hd__buf_12 fanout482 (.A(_03323_),
    .X(net482));
 sky130_fd_sc_hd__clkbuf_16 fanout483 (.A(_03323_),
    .X(net483));
 sky130_fd_sc_hd__buf_12 fanout484 (.A(net485),
    .X(net484));
 sky130_fd_sc_hd__buf_12 fanout485 (.A(_03323_),
    .X(net485));
 sky130_fd_sc_hd__buf_12 fanout486 (.A(net487),
    .X(net486));
 sky130_fd_sc_hd__buf_12 fanout487 (.A(\core_pipeline.decode_to_execute_rs2_bypassed ),
    .X(net487));
 sky130_fd_sc_hd__buf_12 fanout488 (.A(\core_pipeline.decode_to_execute_rs1_bypassed ),
    .X(net488));
 sky130_fd_sc_hd__buf_12 fanout489 (.A(\core_pipeline.decode_to_execute_rs1_bypassed ),
    .X(net489));
 sky130_fd_sc_hd__clkbuf_16 fanout490 (.A(net492),
    .X(net490));
 sky130_fd_sc_hd__buf_4 fanout491 (.A(net492),
    .X(net491));
 sky130_fd_sc_hd__buf_12 fanout492 (.A(\core_busio.mem_address[1] ),
    .X(net492));
 sky130_fd_sc_hd__buf_12 fanout493 (.A(\core_busio.mem_address[0] ),
    .X(net493));
 sky130_fd_sc_hd__clkbuf_16 fanout494 (.A(\core_busio.mem_address[0] ),
    .X(net494));
 sky130_fd_sc_hd__buf_12 fanout495 (.A(\core_busio.mem_address[0] ),
    .X(net495));
 sky130_fd_sc_hd__buf_8 fanout496 (.A(net497),
    .X(net496));
 sky130_fd_sc_hd__buf_6 fanout497 (.A(\core_busio.mem_address[0] ),
    .X(net497));
 sky130_fd_sc_hd__buf_12 fanout498 (.A(net499),
    .X(net498));
 sky130_fd_sc_hd__buf_12 fanout499 (.A(\core_pipeline.execute_to_memory_write_select[0] ),
    .X(net499));
 sky130_fd_sc_hd__buf_6 fanout500 (.A(net501),
    .X(net500));
 sky130_fd_sc_hd__buf_12 fanout501 (.A(\core_pipeline.pipeline_decode.alu_select_b_out[2] ),
    .X(net501));
 sky130_fd_sc_hd__buf_6 fanout502 (.A(net503),
    .X(net502));
 sky130_fd_sc_hd__buf_12 fanout503 (.A(\core_pipeline.pipeline_decode.alu_select_b_out[1] ),
    .X(net503));
 sky130_fd_sc_hd__buf_12 fanout504 (.A(net505),
    .X(net504));
 sky130_fd_sc_hd__buf_12 fanout505 (.A(\core_pipeline.memory_to_writeback_wfi ),
    .X(net505));
 sky130_fd_sc_hd__buf_6 fanout506 (.A(net507),
    .X(net506));
 sky130_fd_sc_hd__buf_4 fanout507 (.A(net508),
    .X(net507));
 sky130_fd_sc_hd__buf_8 fanout508 (.A(\core_pipeline.memory_to_writeback_write_select[1] ),
    .X(net508));
 sky130_fd_sc_hd__buf_8 fanout509 (.A(net510),
    .X(net509));
 sky130_fd_sc_hd__buf_12 fanout510 (.A(\core_pipeline.memory_to_writeback_write_select[0] ),
    .X(net510));
 sky130_fd_sc_hd__buf_12 fanout511 (.A(\core_pipeline.decode_to_csr_read_address[4] ),
    .X(net511));
 sky130_fd_sc_hd__buf_12 fanout512 (.A(\core_pipeline.decode_to_csr_read_address[4] ),
    .X(net512));
 sky130_fd_sc_hd__buf_8 fanout513 (.A(\core_pipeline.decode_to_csr_read_address[4] ),
    .X(net513));
 sky130_fd_sc_hd__buf_12 fanout514 (.A(net515),
    .X(net514));
 sky130_fd_sc_hd__buf_12 fanout515 (.A(\core_pipeline.decode_to_csr_read_address[3] ),
    .X(net515));
 sky130_fd_sc_hd__buf_12 fanout516 (.A(net518),
    .X(net516));
 sky130_fd_sc_hd__buf_12 fanout517 (.A(net518),
    .X(net517));
 sky130_fd_sc_hd__buf_12 fanout518 (.A(\core_pipeline.decode_to_csr_read_address[3] ),
    .X(net518));
 sky130_fd_sc_hd__buf_12 fanout519 (.A(net521),
    .X(net519));
 sky130_fd_sc_hd__clkbuf_8 fanout520 (.A(net521),
    .X(net520));
 sky130_fd_sc_hd__buf_12 fanout521 (.A(\core_pipeline.decode_to_csr_read_address[2] ),
    .X(net521));
 sky130_fd_sc_hd__buf_12 fanout522 (.A(net524),
    .X(net522));
 sky130_fd_sc_hd__buf_12 fanout523 (.A(net524),
    .X(net523));
 sky130_fd_sc_hd__buf_12 fanout524 (.A(\core_pipeline.decode_to_csr_read_address[2] ),
    .X(net524));
 sky130_fd_sc_hd__buf_12 fanout525 (.A(net528),
    .X(net525));
 sky130_fd_sc_hd__buf_12 fanout526 (.A(net528),
    .X(net526));
 sky130_fd_sc_hd__buf_6 fanout527 (.A(net528),
    .X(net527));
 sky130_fd_sc_hd__clkbuf_16 fanout528 (.A(net543),
    .X(net528));
 sky130_fd_sc_hd__buf_12 fanout529 (.A(net531),
    .X(net529));
 sky130_fd_sc_hd__buf_12 fanout530 (.A(net531),
    .X(net530));
 sky130_fd_sc_hd__clkbuf_16 fanout531 (.A(net543),
    .X(net531));
 sky130_fd_sc_hd__buf_12 fanout532 (.A(net533),
    .X(net532));
 sky130_fd_sc_hd__buf_12 fanout533 (.A(net543),
    .X(net533));
 sky130_fd_sc_hd__buf_12 fanout534 (.A(net536),
    .X(net534));
 sky130_fd_sc_hd__buf_12 fanout535 (.A(net536),
    .X(net535));
 sky130_fd_sc_hd__buf_12 fanout536 (.A(net543),
    .X(net536));
 sky130_fd_sc_hd__buf_12 fanout537 (.A(net539),
    .X(net537));
 sky130_fd_sc_hd__buf_12 fanout538 (.A(net539),
    .X(net538));
 sky130_fd_sc_hd__clkbuf_16 fanout539 (.A(net543),
    .X(net539));
 sky130_fd_sc_hd__buf_12 fanout540 (.A(net541),
    .X(net540));
 sky130_fd_sc_hd__buf_8 fanout541 (.A(net542),
    .X(net541));
 sky130_fd_sc_hd__buf_12 fanout542 (.A(net543),
    .X(net542));
 sky130_fd_sc_hd__buf_12 fanout543 (.A(\core_pipeline.decode_to_csr_read_address[1] ),
    .X(net543));
 sky130_fd_sc_hd__buf_12 fanout544 (.A(net547),
    .X(net544));
 sky130_fd_sc_hd__buf_8 fanout545 (.A(net547),
    .X(net545));
 sky130_fd_sc_hd__buf_12 fanout546 (.A(net547),
    .X(net546));
 sky130_fd_sc_hd__buf_12 fanout547 (.A(net566),
    .X(net547));
 sky130_fd_sc_hd__buf_12 fanout548 (.A(net551),
    .X(net548));
 sky130_fd_sc_hd__buf_6 fanout549 (.A(net551),
    .X(net549));
 sky130_fd_sc_hd__buf_12 fanout550 (.A(net551),
    .X(net550));
 sky130_fd_sc_hd__clkbuf_16 fanout551 (.A(net566),
    .X(net551));
 sky130_fd_sc_hd__buf_12 fanout552 (.A(net554),
    .X(net552));
 sky130_fd_sc_hd__buf_6 fanout553 (.A(net554),
    .X(net553));
 sky130_fd_sc_hd__buf_8 fanout554 (.A(net566),
    .X(net554));
 sky130_fd_sc_hd__buf_12 fanout555 (.A(net566),
    .X(net555));
 sky130_fd_sc_hd__buf_6 fanout556 (.A(net566),
    .X(net556));
 sky130_fd_sc_hd__buf_12 fanout557 (.A(net566),
    .X(net557));
 sky130_fd_sc_hd__buf_8 fanout558 (.A(net566),
    .X(net558));
 sky130_fd_sc_hd__buf_12 fanout559 (.A(net562),
    .X(net559));
 sky130_fd_sc_hd__buf_8 fanout560 (.A(net562),
    .X(net560));
 sky130_fd_sc_hd__buf_12 fanout561 (.A(net562),
    .X(net561));
 sky130_fd_sc_hd__buf_12 fanout562 (.A(net566),
    .X(net562));
 sky130_fd_sc_hd__buf_12 fanout563 (.A(net564),
    .X(net563));
 sky130_fd_sc_hd__buf_8 fanout564 (.A(net565),
    .X(net564));
 sky130_fd_sc_hd__buf_12 fanout565 (.A(net566),
    .X(net565));
 sky130_fd_sc_hd__buf_12 fanout566 (.A(\core_pipeline.decode_to_csr_read_address[0] ),
    .X(net566));
 sky130_fd_sc_hd__buf_12 fanout567 (.A(net569),
    .X(net567));
 sky130_fd_sc_hd__buf_12 fanout568 (.A(net569),
    .X(net568));
 sky130_fd_sc_hd__buf_12 fanout569 (.A(\core_pipeline.decode_to_regfile_rs1_address[4] ),
    .X(net569));
 sky130_fd_sc_hd__buf_12 fanout570 (.A(net572),
    .X(net570));
 sky130_fd_sc_hd__clkbuf_16 fanout571 (.A(net572),
    .X(net571));
 sky130_fd_sc_hd__buf_12 fanout572 (.A(\core_pipeline.decode_to_regfile_rs1_address[3] ),
    .X(net572));
 sky130_fd_sc_hd__buf_12 fanout573 (.A(net575),
    .X(net573));
 sky130_fd_sc_hd__buf_12 fanout574 (.A(net575),
    .X(net574));
 sky130_fd_sc_hd__buf_12 fanout575 (.A(\core_pipeline.decode_to_regfile_rs1_address[3] ),
    .X(net575));
 sky130_fd_sc_hd__buf_12 fanout576 (.A(net577),
    .X(net576));
 sky130_fd_sc_hd__buf_12 fanout577 (.A(net578),
    .X(net577));
 sky130_fd_sc_hd__buf_12 fanout578 (.A(\core_pipeline.decode_to_regfile_rs1_address[2] ),
    .X(net578));
 sky130_fd_sc_hd__buf_12 fanout579 (.A(net581),
    .X(net579));
 sky130_fd_sc_hd__buf_12 fanout580 (.A(net581),
    .X(net580));
 sky130_fd_sc_hd__buf_12 fanout581 (.A(\core_pipeline.decode_to_regfile_rs1_address[2] ),
    .X(net581));
 sky130_fd_sc_hd__buf_12 fanout582 (.A(net589),
    .X(net582));
 sky130_fd_sc_hd__buf_6 fanout583 (.A(net589),
    .X(net583));
 sky130_fd_sc_hd__buf_12 fanout584 (.A(net585),
    .X(net584));
 sky130_fd_sc_hd__clkbuf_16 fanout585 (.A(net589),
    .X(net585));
 sky130_fd_sc_hd__clkbuf_16 fanout586 (.A(net589),
    .X(net586));
 sky130_fd_sc_hd__buf_6 fanout587 (.A(net589),
    .X(net587));
 sky130_fd_sc_hd__clkbuf_16 fanout588 (.A(net589),
    .X(net588));
 sky130_fd_sc_hd__buf_12 fanout589 (.A(\core_pipeline.decode_to_regfile_rs1_address[1] ),
    .X(net589));
 sky130_fd_sc_hd__buf_12 fanout590 (.A(net591),
    .X(net590));
 sky130_fd_sc_hd__buf_6 fanout591 (.A(\core_pipeline.decode_to_regfile_rs1_address[1] ),
    .X(net591));
 sky130_fd_sc_hd__buf_12 fanout592 (.A(net600),
    .X(net592));
 sky130_fd_sc_hd__clkbuf_8 fanout593 (.A(net600),
    .X(net593));
 sky130_fd_sc_hd__buf_12 fanout594 (.A(net600),
    .X(net594));
 sky130_fd_sc_hd__buf_6 fanout595 (.A(net600),
    .X(net595));
 sky130_fd_sc_hd__buf_12 fanout596 (.A(net600),
    .X(net596));
 sky130_fd_sc_hd__buf_4 fanout597 (.A(net600),
    .X(net597));
 sky130_fd_sc_hd__buf_12 fanout598 (.A(net600),
    .X(net598));
 sky130_fd_sc_hd__buf_6 fanout599 (.A(net600),
    .X(net599));
 sky130_fd_sc_hd__buf_12 fanout600 (.A(\core_pipeline.decode_to_regfile_rs1_address[1] ),
    .X(net600));
 sky130_fd_sc_hd__buf_12 fanout601 (.A(net602),
    .X(net601));
 sky130_fd_sc_hd__clkbuf_16 fanout602 (.A(\core_pipeline.decode_to_regfile_rs1_address[1] ),
    .X(net602));
 sky130_fd_sc_hd__buf_12 fanout603 (.A(net611),
    .X(net603));
 sky130_fd_sc_hd__clkbuf_16 fanout604 (.A(net611),
    .X(net604));
 sky130_fd_sc_hd__buf_12 fanout605 (.A(net606),
    .X(net605));
 sky130_fd_sc_hd__buf_12 fanout606 (.A(net611),
    .X(net606));
 sky130_fd_sc_hd__buf_12 fanout607 (.A(net608),
    .X(net607));
 sky130_fd_sc_hd__buf_12 fanout608 (.A(net611),
    .X(net608));
 sky130_fd_sc_hd__buf_12 fanout609 (.A(net611),
    .X(net609));
 sky130_fd_sc_hd__buf_12 fanout610 (.A(net611),
    .X(net610));
 sky130_fd_sc_hd__buf_12 fanout611 (.A(net614),
    .X(net611));
 sky130_fd_sc_hd__buf_12 fanout612 (.A(net614),
    .X(net612));
 sky130_fd_sc_hd__buf_12 fanout613 (.A(net614),
    .X(net613));
 sky130_fd_sc_hd__buf_12 fanout614 (.A(\core_pipeline.decode_to_regfile_rs1_address[0] ),
    .X(net614));
 sky130_fd_sc_hd__buf_12 fanout615 (.A(net623),
    .X(net615));
 sky130_fd_sc_hd__buf_12 fanout616 (.A(net623),
    .X(net616));
 sky130_fd_sc_hd__buf_12 fanout617 (.A(net623),
    .X(net617));
 sky130_fd_sc_hd__buf_6 fanout618 (.A(net623),
    .X(net618));
 sky130_fd_sc_hd__buf_12 fanout619 (.A(net623),
    .X(net619));
 sky130_fd_sc_hd__buf_12 fanout620 (.A(net623),
    .X(net620));
 sky130_fd_sc_hd__buf_12 fanout621 (.A(net622),
    .X(net621));
 sky130_fd_sc_hd__buf_12 fanout622 (.A(net623),
    .X(net622));
 sky130_fd_sc_hd__buf_12 fanout623 (.A(\core_pipeline.decode_to_regfile_rs1_address[0] ),
    .X(net623));
 sky130_fd_sc_hd__buf_12 fanout624 (.A(net626),
    .X(net624));
 sky130_fd_sc_hd__buf_6 fanout625 (.A(net626),
    .X(net625));
 sky130_fd_sc_hd__buf_12 fanout626 (.A(\core_pipeline.decode_to_regfile_rs1_address[0] ),
    .X(net626));
 sky130_fd_sc_hd__buf_8 fanout627 (.A(net628),
    .X(net627));
 sky130_fd_sc_hd__buf_12 fanout628 (.A(\core_pipeline.pipeline_decode.alu_select_a_out[2] ),
    .X(net628));
 sky130_fd_sc_hd__buf_8 fanout629 (.A(net630),
    .X(net629));
 sky130_fd_sc_hd__buf_12 fanout630 (.A(\core_pipeline.pipeline_decode.alu_select_a_out[1] ),
    .X(net630));
 sky130_fd_sc_hd__buf_12 fanout631 (.A(net632),
    .X(net631));
 sky130_fd_sc_hd__clkbuf_16 fanout632 (.A(\core_pipeline.decode_to_execute_alu_function_modifier ),
    .X(net632));
 sky130_fd_sc_hd__buf_8 fanout633 (.A(\core_pipeline.decode_to_execute_alu_function_modifier ),
    .X(net633));
 sky130_fd_sc_hd__buf_6 fanout634 (.A(net635),
    .X(net634));
 sky130_fd_sc_hd__clkbuf_16 fanout635 (.A(\core_pipeline.decode_to_execute_alu_function_modifier ),
    .X(net635));
 sky130_fd_sc_hd__clkbuf_16 fanout636 (.A(net647),
    .X(net636));
 sky130_fd_sc_hd__buf_6 fanout637 (.A(net647),
    .X(net637));
 sky130_fd_sc_hd__buf_12 fanout638 (.A(net647),
    .X(net638));
 sky130_fd_sc_hd__buf_8 fanout639 (.A(net647),
    .X(net639));
 sky130_fd_sc_hd__buf_4 fanout640 (.A(net647),
    .X(net640));
 sky130_fd_sc_hd__buf_8 fanout641 (.A(net647),
    .X(net641));
 sky130_fd_sc_hd__clkbuf_8 fanout642 (.A(net647),
    .X(net642));
 sky130_fd_sc_hd__buf_8 fanout643 (.A(net646),
    .X(net643));
 sky130_fd_sc_hd__buf_8 fanout644 (.A(net646),
    .X(net644));
 sky130_fd_sc_hd__buf_6 fanout645 (.A(net646),
    .X(net645));
 sky130_fd_sc_hd__buf_8 fanout646 (.A(net647),
    .X(net646));
 sky130_fd_sc_hd__buf_12 fanout647 (.A(_03338_),
    .X(net647));
 sky130_fd_sc_hd__bufbuf_16 hold1 (.A(\core_pipeline.decode_to_execute_branch ),
    .X(net651));
 sky130_fd_sc_hd__bufbuf_16 hold2 (.A(\core_pipeline.decode_to_execute_next_pc[17] ),
    .X(net652));
 sky130_fd_sc_hd__bufbuf_16 hold3 (.A(\core_pipeline.decode_to_execute_load_signed ),
    .X(net653));
 sky130_fd_sc_hd__bufbuf_16 hold4 (.A(\core_pipeline.fetch_to_decode_instruction[10] ),
    .X(net654));
 sky130_fd_sc_hd__bufbuf_16 hold5 (.A(\core_pipeline.fetch_to_decode_instruction[7] ),
    .X(net655));
 sky130_fd_sc_hd__bufbuf_16 hold6 (.A(\core_pipeline.execute_to_memory_pc[29] ),
    .X(net656));
 sky130_fd_sc_hd__bufbuf_16 hold7 (.A(\core_pipeline.execute_to_memory_next_pc[8] ),
    .X(net657));
 sky130_fd_sc_hd__bufbuf_16 hold8 (.A(\core_pipeline.fetch_to_decode_instruction[11] ),
    .X(net658));
 sky130_fd_sc_hd__bufbuf_16 hold9 (.A(\core_pipeline.decode_to_execute_next_pc[25] ),
    .X(net659));
 sky130_fd_sc_hd__buf_4 input1 (.A(ext_read_data[0]),
    .X(net1));
 sky130_fd_sc_hd__buf_6 input10 (.A(ext_read_data[18]),
    .X(net10));
 sky130_fd_sc_hd__buf_4 input11 (.A(ext_read_data[19]),
    .X(net11));
 sky130_fd_sc_hd__buf_6 input12 (.A(ext_read_data[1]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_4 input13 (.A(ext_read_data[20]),
    .X(net13));
 sky130_fd_sc_hd__buf_4 input14 (.A(ext_read_data[21]),
    .X(net14));
 sky130_fd_sc_hd__buf_4 input15 (.A(ext_read_data[22]),
    .X(net15));
 sky130_fd_sc_hd__buf_8 input16 (.A(ext_read_data[23]),
    .X(net16));
 sky130_fd_sc_hd__buf_6 input17 (.A(ext_read_data[24]),
    .X(net17));
 sky130_fd_sc_hd__buf_6 input18 (.A(ext_read_data[25]),
    .X(net18));
 sky130_fd_sc_hd__buf_8 input19 (.A(ext_read_data[26]),
    .X(net19));
 sky130_fd_sc_hd__buf_6 input2 (.A(ext_read_data[10]),
    .X(net2));
 sky130_fd_sc_hd__buf_8 input20 (.A(ext_read_data[27]),
    .X(net20));
 sky130_fd_sc_hd__buf_8 input21 (.A(ext_read_data[28]),
    .X(net21));
 sky130_fd_sc_hd__buf_6 input22 (.A(ext_read_data[29]),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_4 input23 (.A(ext_read_data[2]),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_16 input24 (.A(ext_read_data[30]),
    .X(net24));
 sky130_fd_sc_hd__buf_6 input25 (.A(ext_read_data[31]),
    .X(net25));
 sky130_fd_sc_hd__buf_6 input26 (.A(ext_read_data[3]),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_8 input27 (.A(ext_read_data[4]),
    .X(net27));
 sky130_fd_sc_hd__buf_6 input28 (.A(ext_read_data[5]),
    .X(net28));
 sky130_fd_sc_hd__buf_6 input29 (.A(ext_read_data[6]),
    .X(net29));
 sky130_fd_sc_hd__buf_6 input3 (.A(ext_read_data[11]),
    .X(net3));
 sky130_fd_sc_hd__buf_4 input30 (.A(ext_read_data[7]),
    .X(net30));
 sky130_fd_sc_hd__buf_8 input31 (.A(ext_read_data[8]),
    .X(net31));
 sky130_fd_sc_hd__buf_4 input32 (.A(ext_read_data[9]),
    .X(net32));
 sky130_fd_sc_hd__buf_4 input33 (.A(ext_ready),
    .X(net33));
 sky130_fd_sc_hd__buf_6 input34 (.A(meip),
    .X(net34));
 sky130_fd_sc_hd__buf_12 input35 (.A(reset),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_8 input4 (.A(ext_read_data[12]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_8 input5 (.A(ext_read_data[13]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_4 input6 (.A(ext_read_data[14]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_4 input7 (.A(ext_read_data[15]),
    .X(net7));
 sky130_fd_sc_hd__buf_4 input8 (.A(ext_read_data[16]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_4 input9 (.A(ext_read_data[17]),
    .X(net9));
 sky130_fd_sc_hd__buf_2 max_cap281 (.A(_04111_),
    .X(net281));
 sky130_fd_sc_hd__buf_6 max_cap371 (.A(_04590_),
    .X(net371));
 sky130_fd_sc_hd__buf_4 max_cap437 (.A(net438),
    .X(net437));
 sky130_fd_sc_hd__clkbuf_2 output100 (.A(net100),
    .X(ext_write_strobe[1]));
 sky130_fd_sc_hd__clkbuf_2 output101 (.A(net101),
    .X(ext_write_strobe[2]));
 sky130_fd_sc_hd__clkbuf_2 output102 (.A(net102),
    .X(ext_write_strobe[3]));
 sky130_fd_sc_hd__clkbuf_2 output36 (.A(net36),
    .X(ext_address[10]));
 sky130_fd_sc_hd__clkbuf_2 output37 (.A(net37),
    .X(ext_address[11]));
 sky130_fd_sc_hd__clkbuf_2 output38 (.A(net38),
    .X(ext_address[12]));
 sky130_fd_sc_hd__clkbuf_2 output39 (.A(net39),
    .X(ext_address[13]));
 sky130_fd_sc_hd__clkbuf_2 output40 (.A(net40),
    .X(ext_address[14]));
 sky130_fd_sc_hd__clkbuf_2 output41 (.A(net41),
    .X(ext_address[15]));
 sky130_fd_sc_hd__clkbuf_2 output42 (.A(net42),
    .X(ext_address[16]));
 sky130_fd_sc_hd__clkbuf_2 output43 (.A(net43),
    .X(ext_address[17]));
 sky130_fd_sc_hd__clkbuf_2 output44 (.A(net44),
    .X(ext_address[18]));
 sky130_fd_sc_hd__clkbuf_2 output45 (.A(net45),
    .X(ext_address[19]));
 sky130_fd_sc_hd__clkbuf_2 output46 (.A(net46),
    .X(ext_address[20]));
 sky130_fd_sc_hd__clkbuf_2 output47 (.A(net47),
    .X(ext_address[21]));
 sky130_fd_sc_hd__clkbuf_2 output48 (.A(net48),
    .X(ext_address[22]));
 sky130_fd_sc_hd__clkbuf_2 output49 (.A(net49),
    .X(ext_address[23]));
 sky130_fd_sc_hd__clkbuf_2 output50 (.A(net50),
    .X(ext_address[24]));
 sky130_fd_sc_hd__clkbuf_2 output51 (.A(net51),
    .X(ext_address[25]));
 sky130_fd_sc_hd__clkbuf_2 output52 (.A(net52),
    .X(ext_address[26]));
 sky130_fd_sc_hd__clkbuf_2 output53 (.A(net53),
    .X(ext_address[27]));
 sky130_fd_sc_hd__clkbuf_2 output54 (.A(net54),
    .X(ext_address[28]));
 sky130_fd_sc_hd__clkbuf_2 output55 (.A(net55),
    .X(ext_address[29]));
 sky130_fd_sc_hd__clkbuf_2 output56 (.A(net56),
    .X(ext_address[2]));
 sky130_fd_sc_hd__clkbuf_2 output57 (.A(net57),
    .X(ext_address[30]));
 sky130_fd_sc_hd__clkbuf_2 output58 (.A(net58),
    .X(ext_address[31]));
 sky130_fd_sc_hd__clkbuf_2 output59 (.A(net59),
    .X(ext_address[3]));
 sky130_fd_sc_hd__clkbuf_2 output60 (.A(net60),
    .X(ext_address[4]));
 sky130_fd_sc_hd__clkbuf_2 output61 (.A(net61),
    .X(ext_address[5]));
 sky130_fd_sc_hd__clkbuf_2 output62 (.A(net62),
    .X(ext_address[6]));
 sky130_fd_sc_hd__clkbuf_2 output63 (.A(net63),
    .X(ext_address[7]));
 sky130_fd_sc_hd__clkbuf_2 output64 (.A(net64),
    .X(ext_address[8]));
 sky130_fd_sc_hd__clkbuf_2 output65 (.A(net65),
    .X(ext_address[9]));
 sky130_fd_sc_hd__clkbuf_2 output66 (.A(net66),
    .X(ext_instruction));
 sky130_fd_sc_hd__clkbuf_2 output67 (.A(net67),
    .X(ext_write_data[0]));
 sky130_fd_sc_hd__clkbuf_2 output68 (.A(net68),
    .X(ext_write_data[10]));
 sky130_fd_sc_hd__clkbuf_2 output69 (.A(net69),
    .X(ext_write_data[11]));
 sky130_fd_sc_hd__clkbuf_2 output70 (.A(net70),
    .X(ext_write_data[12]));
 sky130_fd_sc_hd__clkbuf_2 output71 (.A(net71),
    .X(ext_write_data[13]));
 sky130_fd_sc_hd__clkbuf_2 output72 (.A(net72),
    .X(ext_write_data[14]));
 sky130_fd_sc_hd__clkbuf_2 output73 (.A(net73),
    .X(ext_write_data[15]));
 sky130_fd_sc_hd__clkbuf_2 output74 (.A(net74),
    .X(ext_write_data[16]));
 sky130_fd_sc_hd__clkbuf_2 output75 (.A(net75),
    .X(ext_write_data[17]));
 sky130_fd_sc_hd__clkbuf_2 output76 (.A(net76),
    .X(ext_write_data[18]));
 sky130_fd_sc_hd__clkbuf_2 output77 (.A(net77),
    .X(ext_write_data[19]));
 sky130_fd_sc_hd__clkbuf_2 output78 (.A(net78),
    .X(ext_write_data[1]));
 sky130_fd_sc_hd__clkbuf_2 output79 (.A(net79),
    .X(ext_write_data[20]));
 sky130_fd_sc_hd__clkbuf_2 output80 (.A(net80),
    .X(ext_write_data[21]));
 sky130_fd_sc_hd__clkbuf_2 output81 (.A(net81),
    .X(ext_write_data[22]));
 sky130_fd_sc_hd__clkbuf_2 output82 (.A(net82),
    .X(ext_write_data[23]));
 sky130_fd_sc_hd__clkbuf_2 output83 (.A(net83),
    .X(ext_write_data[24]));
 sky130_fd_sc_hd__clkbuf_2 output84 (.A(net84),
    .X(ext_write_data[25]));
 sky130_fd_sc_hd__clkbuf_2 output85 (.A(net85),
    .X(ext_write_data[26]));
 sky130_fd_sc_hd__clkbuf_2 output86 (.A(net86),
    .X(ext_write_data[27]));
 sky130_fd_sc_hd__clkbuf_2 output87 (.A(net87),
    .X(ext_write_data[28]));
 sky130_fd_sc_hd__clkbuf_2 output88 (.A(net88),
    .X(ext_write_data[29]));
 sky130_fd_sc_hd__clkbuf_2 output89 (.A(net89),
    .X(ext_write_data[2]));
 sky130_fd_sc_hd__clkbuf_2 output90 (.A(net90),
    .X(ext_write_data[30]));
 sky130_fd_sc_hd__clkbuf_2 output91 (.A(net91),
    .X(ext_write_data[31]));
 sky130_fd_sc_hd__clkbuf_2 output92 (.A(net92),
    .X(ext_write_data[3]));
 sky130_fd_sc_hd__clkbuf_2 output93 (.A(net93),
    .X(ext_write_data[4]));
 sky130_fd_sc_hd__clkbuf_2 output94 (.A(net94),
    .X(ext_write_data[5]));
 sky130_fd_sc_hd__clkbuf_2 output95 (.A(net95),
    .X(ext_write_data[6]));
 sky130_fd_sc_hd__clkbuf_2 output96 (.A(net96),
    .X(ext_write_data[7]));
 sky130_fd_sc_hd__clkbuf_2 output97 (.A(net97),
    .X(ext_write_data[8]));
 sky130_fd_sc_hd__clkbuf_2 output98 (.A(net98),
    .X(ext_write_data[9]));
 sky130_fd_sc_hd__clkbuf_2 output99 (.A(net99),
    .X(ext_write_strobe[0]));
 sky130_fd_sc_hd__buf_6 wire360 (.A(_05724_),
    .X(net360));
 sky130_fd_sc_hd__buf_4 wire438 (.A(_04471_),
    .X(net438));
 assign ext_address[0] = net648;
 assign ext_address[1] = net649;
 assign ext_valid = net650;
endmodule

